module ray_dispatch(
  input         clock,
  input         reset,
  input         io_dispatch,
  input         io_dispatch_2,
  output [31:0] io_rayid_id,
  output [31:0] io_rayid_id_2,
  output        io_ray_out,
  output        io_ray_out_2,
  output        io_ray_finish
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] count; // @[ray_dispatch.scala 21:37]
  reg [31:0] ray_id; // @[ray_dispatch.scala 22:37]
  reg [31:0] ray_id_2; // @[ray_dispatch.scala 23:33]
  reg  ray_out; // @[ray_dispatch.scala 25:35]
  reg  ray_out_2; // @[ray_dispatch.scala 26:32]
  reg [31:0] base; // @[ray_dispatch.scala 28:38]
  wire [31:0] _T_2 = count - 32'h2; // @[ray_dispatch.scala 33:39]
  wire [31:0] _T_5 = base + 32'h1; // @[ray_dispatch.scala 39:38]
  wire [31:0] _T_7 = base + 32'h2; // @[ray_dispatch.scala 40:35]
  wire  _GEN_5 = count >= 32'h1 | ray_out; // @[ray_dispatch.scala 38:27 ray_dispatch.scala 44:29 ray_dispatch.scala 25:35]
  wire  _GEN_6 = count >= 32'h1 | ray_out_2; // @[ray_dispatch.scala 38:27 ray_dispatch.scala 45:26 ray_dispatch.scala 26:32]
  wire  _GEN_11 = count == 32'h46 | _GEN_5; // @[ray_dispatch.scala 30:23 ray_dispatch.scala 35:29]
  wire  _GEN_12 = count == 32'h46 | _GEN_6; // @[ray_dispatch.scala 30:23 ray_dispatch.scala 36:26]
  wire [20:0] _T_17 = 21'h1e8480 - 21'h1; // @[ray_dispatch.scala 67:80]
  wire [31:0] _GEN_47 = {{11'd0}, _T_17}; // @[ray_dispatch.scala 67:67]
  wire  _T_18 = ray_id < _GEN_47; // @[ray_dispatch.scala 67:67]
  wire  _T_41 = io_dispatch & io_dispatch_2 & _T_18; // @[ray_dispatch.scala 83:63]
  wire [31:0] _GEN_19 = io_dispatch & io_dispatch_2 & _T_18 ? _T_5 : ray_id; // @[ray_dispatch.scala 83:91 ray_dispatch.scala 84:30]
  wire [31:0] _GEN_20 = io_dispatch & io_dispatch_2 & _T_18 ? _T_7 : ray_id_2; // @[ray_dispatch.scala 83:91 ray_dispatch.scala 85:27]
  wire [31:0] _GEN_21 = io_dispatch & io_dispatch_2 & _T_18 ? _T_7 : base; // @[ray_dispatch.scala 83:91 ray_dispatch.scala 86:31]
  wire  _GEN_29 = ~io_dispatch & io_dispatch_2 & _T_18 ? 1'h0 : _T_41; // @[ray_dispatch.scala 75:91 ray_dispatch.scala 80:28]
  wire  _GEN_30 = ~io_dispatch & io_dispatch_2 & _T_18 | _T_41; // @[ray_dispatch.scala 75:91 ray_dispatch.scala 81:26]
  wire  _GEN_36 = io_dispatch & ~io_dispatch_2 & ray_id < _GEN_47 | _GEN_29; // @[ray_dispatch.scala 67:85 ray_dispatch.scala 72:28]
  assign io_rayid_id = ray_id; // @[ray_dispatch.scala 122:25]
  assign io_rayid_id_2 = ray_id_2; // @[ray_dispatch.scala 123:22]
  assign io_ray_out = ray_out; // @[ray_dispatch.scala 125:25]
  assign io_ray_out_2 = ray_out_2; // @[ray_dispatch.scala 126:22]
  assign io_ray_finish = ray_id == 32'h1e8480; // @[ray_dispatch.scala 116:17]
  always @(posedge clock) begin
    if (reset) begin // @[ray_dispatch.scala 21:37]
      count <= 32'h46; // @[ray_dispatch.scala 21:37]
    end else if (count == 32'h46) begin // @[ray_dispatch.scala 30:23]
      count <= _T_2; // @[ray_dispatch.scala 33:30]
    end else if (count >= 32'h1) begin // @[ray_dispatch.scala 38:27]
      count <= _T_2; // @[ray_dispatch.scala 42:30]
    end
    if (reset) begin // @[ray_dispatch.scala 22:37]
      ray_id <= 32'h0; // @[ray_dispatch.scala 22:37]
    end else if (count == 32'h0) begin // @[ray_dispatch.scala 66:23]
      if (io_dispatch & ~io_dispatch_2 & ray_id < _GEN_47) begin // @[ray_dispatch.scala 67:85]
        ray_id <= _T_5; // @[ray_dispatch.scala 68:30]
      end else if (!(~io_dispatch & io_dispatch_2 & _T_18)) begin // @[ray_dispatch.scala 75:91]
        ray_id <= _GEN_19;
      end
    end else if (count == 32'h46) begin // @[ray_dispatch.scala 30:23]
      ray_id <= 32'h0; // @[ray_dispatch.scala 31:30]
    end else if (count >= 32'h1) begin // @[ray_dispatch.scala 38:27]
      ray_id <= _T_5; // @[ray_dispatch.scala 39:30]
    end
    if (reset) begin // @[ray_dispatch.scala 23:33]
      ray_id_2 <= 32'h0; // @[ray_dispatch.scala 23:33]
    end else if (count == 32'h0) begin // @[ray_dispatch.scala 66:23]
      if (!(io_dispatch & ~io_dispatch_2 & ray_id < _GEN_47)) begin // @[ray_dispatch.scala 67:85]
        if (~io_dispatch & io_dispatch_2 & _T_18) begin // @[ray_dispatch.scala 75:91]
          ray_id_2 <= _T_5; // @[ray_dispatch.scala 77:27]
        end else begin
          ray_id_2 <= _GEN_20;
        end
      end
    end else if (count == 32'h46) begin // @[ray_dispatch.scala 30:23]
      ray_id_2 <= 32'h1; // @[ray_dispatch.scala 32:27]
    end else if (count >= 32'h1) begin // @[ray_dispatch.scala 38:27]
      ray_id_2 <= _T_7; // @[ray_dispatch.scala 40:27]
    end
    if (reset) begin // @[ray_dispatch.scala 25:35]
      ray_out <= 1'h0; // @[ray_dispatch.scala 25:35]
    end else if (count == 32'h0) begin // @[ray_dispatch.scala 66:23]
      ray_out <= _GEN_36;
    end else begin
      ray_out <= _GEN_11;
    end
    if (reset) begin // @[ray_dispatch.scala 26:32]
      ray_out_2 <= 1'h0; // @[ray_dispatch.scala 26:32]
    end else if (count == 32'h0) begin // @[ray_dispatch.scala 66:23]
      if (io_dispatch & ~io_dispatch_2 & ray_id < _GEN_47) begin // @[ray_dispatch.scala 67:85]
        ray_out_2 <= 1'h0; // @[ray_dispatch.scala 73:25]
      end else begin
        ray_out_2 <= _GEN_30;
      end
    end else begin
      ray_out_2 <= _GEN_12;
    end
    if (reset) begin // @[ray_dispatch.scala 28:38]
      base <= 32'h0; // @[ray_dispatch.scala 28:38]
    end else if (count == 32'h0) begin // @[ray_dispatch.scala 66:23]
      if (io_dispatch & ~io_dispatch_2 & ray_id < _GEN_47) begin // @[ray_dispatch.scala 67:85]
        base <= _T_5; // @[ray_dispatch.scala 70:31]
      end else if (~io_dispatch & io_dispatch_2 & _T_18) begin // @[ray_dispatch.scala 75:91]
        base <= _T_5; // @[ray_dispatch.scala 78:31]
      end else begin
        base <= _GEN_21;
      end
    end else if (count == 32'h46) begin // @[ray_dispatch.scala 30:23]
      base <= 32'h1; // @[ray_dispatch.scala 37:33]
    end else if (count >= 32'h1) begin // @[ray_dispatch.scala 38:27]
      base <= _T_7; // @[ray_dispatch.scala 41:31]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  ray_id = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  ray_id_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  ray_out = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  ray_out_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  base = _RAND_5[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ray_memory(
  input         clock,
  input  [31:0] io_Ray_id,
  input  [31:0] io_Ray_id_2,
  output [31:0] io_Ray_out,
  output [31:0] io_Ray_out_2
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] mem [0:2073599]; // @[ray_memory.scala 16:26]
  wire [31:0] mem_MPORT_data; // @[ray_memory.scala 16:26]
  wire [20:0] mem_MPORT_addr; // @[ray_memory.scala 16:26]
  wire [31:0] mem_MPORT_1_data; // @[ray_memory.scala 16:26]
  wire [20:0] mem_MPORT_1_addr; // @[ray_memory.scala 16:26]
  wire [31:0] mem_MPORT_2_data; // @[ray_memory.scala 16:26]
  wire [20:0] mem_MPORT_2_addr; // @[ray_memory.scala 16:26]
  wire  mem_MPORT_2_mask; // @[ray_memory.scala 16:26]
  wire  mem_MPORT_2_en; // @[ray_memory.scala 16:26]
  reg [20:0] mem_MPORT_addr_pipe_0;
  reg [20:0] mem_MPORT_1_addr_pipe_0;
  assign mem_MPORT_addr = mem_MPORT_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_data = mem[mem_MPORT_addr]; // @[ray_memory.scala 16:26]
  `else
  assign mem_MPORT_data = mem_MPORT_addr >= 21'h1fa400 ? _RAND_1[31:0] : mem[mem_MPORT_addr]; // @[ray_memory.scala 16:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_1_addr = mem_MPORT_1_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_1_data = mem[mem_MPORT_1_addr]; // @[ray_memory.scala 16:26]
  `else
  assign mem_MPORT_1_data = mem_MPORT_1_addr >= 21'h1fa400 ? _RAND_2[31:0] : mem[mem_MPORT_1_addr]; // @[ray_memory.scala 16:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_2_data = 32'h0;
  assign mem_MPORT_2_addr = 21'h0;
  assign mem_MPORT_2_mask = 1'h1;
  assign mem_MPORT_2_en = 1'h0;
  assign io_Ray_out = mem_MPORT_data; // @[ray_memory.scala 18:16]
  assign io_Ray_out_2 = mem_MPORT_1_data; // @[ray_memory.scala 19:18]
  always @(posedge clock) begin
    if(mem_MPORT_2_en & mem_MPORT_2_mask) begin
      mem[mem_MPORT_2_addr] <= mem_MPORT_2_data; // @[ray_memory.scala 16:26]
    end
    mem_MPORT_addr_pipe_0 <= io_Ray_id[20:0];
    mem_MPORT_1_addr_pipe_0 <= io_Ray_id_2[20:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {1{`RANDOM}};
  _RAND_2 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2073600; initvar = initvar+1)
    mem[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  mem_MPORT_addr_pipe_0 = _RAND_3[20:0];
  _RAND_4 = {1{`RANDOM}};
  mem_MPORT_1_addr_pipe_0 = _RAND_4[20:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BVH_memory(
  input         clock,
  input  [31:0] io_BVH_id,
  input  [31:0] io_BVH_id_2,
  output [31:0] io_BVH_out,
  output [31:0] io_BVH_out_2
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg /* sparse */ [31:0] mem [0:21005099]; // @[BVH_memory.scala 16:26]
  wire [31:0] mem_MPORT_data; // @[BVH_memory.scala 16:26]
  wire [24:0] mem_MPORT_addr; // @[BVH_memory.scala 16:26]
  wire [31:0] mem_MPORT_1_data; // @[BVH_memory.scala 16:26]
  wire [24:0] mem_MPORT_1_addr; // @[BVH_memory.scala 16:26]
  wire [31:0] mem_MPORT_2_data; // @[BVH_memory.scala 16:26]
  wire [24:0] mem_MPORT_2_addr; // @[BVH_memory.scala 16:26]
  wire  mem_MPORT_2_mask; // @[BVH_memory.scala 16:26]
  wire  mem_MPORT_2_en; // @[BVH_memory.scala 16:26]
  reg [24:0] mem_MPORT_addr_pipe_0;
  reg [24:0] mem_MPORT_1_addr_pipe_0;
  wire [31:0] _T = io_BVH_id; // @[BVH_memory.scala 18:38]
  wire [31:0] _T_2 = io_BVH_id_2; // @[BVH_memory.scala 19:42]
  assign mem_MPORT_addr = mem_MPORT_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_data = mem[mem_MPORT_addr]; // @[BVH_memory.scala 16:26]
  `else
  assign mem_MPORT_data = mem_MPORT_addr >= 25'h140832c ? _RAND_1[31:0] : mem[mem_MPORT_addr]; // @[BVH_memory.scala 16:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_1_addr = mem_MPORT_1_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_1_data = mem[mem_MPORT_1_addr]; // @[BVH_memory.scala 16:26]
  `else
  assign mem_MPORT_1_data = mem_MPORT_1_addr >= 25'h140832c ? _RAND_2[31:0] : mem[mem_MPORT_1_addr]; // @[BVH_memory.scala 16:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_2_data = 32'h0;
  assign mem_MPORT_2_addr = 25'h0;
  assign mem_MPORT_2_mask = 1'h1;
  assign mem_MPORT_2_en = 1'h0;
  assign io_BVH_out = mem_MPORT_data; // @[BVH_memory.scala 18:16]
  assign io_BVH_out_2 = mem_MPORT_1_data; // @[BVH_memory.scala 19:18]
  always @(posedge clock) begin
    if(mem_MPORT_2_en & mem_MPORT_2_mask) begin
      mem[mem_MPORT_2_addr] <= mem_MPORT_2_data; // @[BVH_memory.scala 16:26]
    end
    mem_MPORT_addr_pipe_0 <= _T[24:0];
    mem_MPORT_1_addr_pipe_0 <= _T_2[24:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {1{`RANDOM}};
  _RAND_2 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 21005100; initvar = initvar+1)
    mem[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  mem_MPORT_addr_pipe_0 = _RAND_3[24:0];
  _RAND_4 = {1{`RANDOM}};
  mem_MPORT_1_addr_pipe_0 = _RAND_4[24:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BVH_memory_0(
  input         clock,
  input  [31:0] io_BVH_id,
  input  [31:0] io_BVH_id_2,
  output [31:0] io_BVH_out,
  output [31:0] io_BVH_out_2
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg /* sparse */ [31:0] mem [0:21005099]; // @[BVH_memory_0.scala 16:26]
  wire [31:0] mem_MPORT_data; // @[BVH_memory_0.scala 16:26]
  wire [24:0] mem_MPORT_addr; // @[BVH_memory_0.scala 16:26]
  wire [31:0] mem_MPORT_1_data; // @[BVH_memory_0.scala 16:26]
  wire [24:0] mem_MPORT_1_addr; // @[BVH_memory_0.scala 16:26]
  wire [31:0] mem_MPORT_2_data; // @[BVH_memory_0.scala 16:26]
  wire [24:0] mem_MPORT_2_addr; // @[BVH_memory_0.scala 16:26]
  wire  mem_MPORT_2_mask; // @[BVH_memory_0.scala 16:26]
  wire  mem_MPORT_2_en; // @[BVH_memory_0.scala 16:26]
  reg [24:0] mem_MPORT_addr_pipe_0;
  reg [24:0] mem_MPORT_1_addr_pipe_0;
  wire [31:0] _T = io_BVH_id; // @[BVH_memory_0.scala 18:38]
  wire [31:0] _T_2 = io_BVH_id_2; // @[BVH_memory_0.scala 19:42]
  assign mem_MPORT_addr = mem_MPORT_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_data = mem[mem_MPORT_addr]; // @[BVH_memory_0.scala 16:26]
  `else
  assign mem_MPORT_data = mem_MPORT_addr >= 25'h140832c ? _RAND_1[31:0] : mem[mem_MPORT_addr]; // @[BVH_memory_0.scala 16:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_1_addr = mem_MPORT_1_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_1_data = mem[mem_MPORT_1_addr]; // @[BVH_memory_0.scala 16:26]
  `else
  assign mem_MPORT_1_data = mem_MPORT_1_addr >= 25'h140832c ? _RAND_2[31:0] : mem[mem_MPORT_1_addr]; // @[BVH_memory_0.scala 16:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_2_data = 32'sh0;
  assign mem_MPORT_2_addr = 25'h0;
  assign mem_MPORT_2_mask = 1'h1;
  assign mem_MPORT_2_en = 1'h0;
  assign io_BVH_out = mem_MPORT_data; // @[BVH_memory_0.scala 18:16]
  assign io_BVH_out_2 = mem_MPORT_1_data; // @[BVH_memory_0.scala 19:18]
  always @(posedge clock) begin
    if(mem_MPORT_2_en & mem_MPORT_2_mask) begin
      mem[mem_MPORT_2_addr] <= mem_MPORT_2_data; // @[BVH_memory_0.scala 16:26]
    end
    mem_MPORT_addr_pipe_0 <= _T[24:0];
    mem_MPORT_1_addr_pipe_0 <= _T_2[24:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {1{`RANDOM}};
  _RAND_2 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 21005100; initvar = initvar+1)
    mem[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  mem_MPORT_addr_pipe_0 = _RAND_3[24:0];
  _RAND_4 = {1{`RANDOM}};
  mem_MPORT_1_addr_pipe_0 = _RAND_4[24:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Triangle_memory_valid(
  input         clock,
  input  [31:0] io_Triangle_id,
  output [31:0] io_v00_out,
  output [31:0] io_v11_out,
  output [31:0] io_v22_out,
  output [31:0] io_valid
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg /* sparse */ [31:0] mem [0:51005099]; // @[Triangle_memory_valid.scala 18:26]
  wire [31:0] mem_MPORT_data; // @[Triangle_memory_valid.scala 18:26]
  wire [25:0] mem_MPORT_addr; // @[Triangle_memory_valid.scala 18:26]
  wire [31:0] mem_MPORT_1_data; // @[Triangle_memory_valid.scala 18:26]
  wire [25:0] mem_MPORT_1_addr; // @[Triangle_memory_valid.scala 18:26]
  wire [31:0] mem_MPORT_2_data; // @[Triangle_memory_valid.scala 18:26]
  wire [25:0] mem_MPORT_2_addr; // @[Triangle_memory_valid.scala 18:26]
  wire [31:0] mem_MPORT_3_data; // @[Triangle_memory_valid.scala 18:26]
  wire [25:0] mem_MPORT_3_addr; // @[Triangle_memory_valid.scala 18:26]
  wire [31:0] mem_MPORT_4_data; // @[Triangle_memory_valid.scala 18:26]
  wire [25:0] mem_MPORT_4_addr; // @[Triangle_memory_valid.scala 18:26]
  wire  mem_MPORT_4_mask; // @[Triangle_memory_valid.scala 18:26]
  wire  mem_MPORT_4_en; // @[Triangle_memory_valid.scala 18:26]
  reg [25:0] mem_MPORT_addr_pipe_0;
  reg [25:0] mem_MPORT_1_addr_pipe_0;
  reg [25:0] mem_MPORT_2_addr_pipe_0;
  reg [25:0] mem_MPORT_3_addr_pipe_0;
  wire [31:0] _T = io_Triangle_id; // @[Triangle_memory_valid.scala 20:43]
  wire [31:0] _T_4 = io_Triangle_id + 32'h1; // @[Triangle_memory_valid.scala 21:49]
  wire [31:0] _T_8 = io_Triangle_id + 32'h2; // @[Triangle_memory_valid.scala 22:49]
  wire [31:0] _T_12 = io_Triangle_id + 32'h3; // @[Triangle_memory_valid.scala 23:47]
  assign mem_MPORT_addr = mem_MPORT_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_data = mem[mem_MPORT_addr]; // @[Triangle_memory_valid.scala 18:26]
  `else
  assign mem_MPORT_data = mem_MPORT_addr >= 26'h30a46ac ? _RAND_1[31:0] : mem[mem_MPORT_addr]; // @[Triangle_memory_valid.scala 18:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_1_addr = mem_MPORT_1_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_1_data = mem[mem_MPORT_1_addr]; // @[Triangle_memory_valid.scala 18:26]
  `else
  assign mem_MPORT_1_data = mem_MPORT_1_addr >= 26'h30a46ac ? _RAND_2[31:0] : mem[mem_MPORT_1_addr]; // @[Triangle_memory_valid.scala 18:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_2_addr = mem_MPORT_2_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_2_data = mem[mem_MPORT_2_addr]; // @[Triangle_memory_valid.scala 18:26]
  `else
  assign mem_MPORT_2_data = mem_MPORT_2_addr >= 26'h30a46ac ? _RAND_3[31:0] : mem[mem_MPORT_2_addr]; // @[Triangle_memory_valid.scala 18:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_3_addr = mem_MPORT_3_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_3_data = mem[mem_MPORT_3_addr]; // @[Triangle_memory_valid.scala 18:26]
  `else
  assign mem_MPORT_3_data = mem_MPORT_3_addr >= 26'h30a46ac ? _RAND_4[31:0] : mem[mem_MPORT_3_addr]; // @[Triangle_memory_valid.scala 18:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_4_data = 32'h0;
  assign mem_MPORT_4_addr = 26'h0;
  assign mem_MPORT_4_mask = 1'h1;
  assign mem_MPORT_4_en = 1'h0;
  assign io_v00_out = mem_MPORT_data; // @[Triangle_memory_valid.scala 20:16]
  assign io_v11_out = mem_MPORT_1_data; // @[Triangle_memory_valid.scala 21:16]
  assign io_v22_out = mem_MPORT_2_data; // @[Triangle_memory_valid.scala 22:16]
  assign io_valid = mem_MPORT_3_data; // @[Triangle_memory_valid.scala 23:14]
  always @(posedge clock) begin
    if(mem_MPORT_4_en & mem_MPORT_4_mask) begin
      mem[mem_MPORT_4_addr] <= mem_MPORT_4_data; // @[Triangle_memory_valid.scala 18:26]
    end
    mem_MPORT_addr_pipe_0 <= _T[25:0];
    mem_MPORT_1_addr_pipe_0 <= _T_4[25:0];
    mem_MPORT_2_addr_pipe_0 <= _T_8[25:0];
    mem_MPORT_3_addr_pipe_0 <= _T_12[25:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {1{`RANDOM}};
  _RAND_2 = {1{`RANDOM}};
  _RAND_3 = {1{`RANDOM}};
  _RAND_4 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 51005100; initvar = initvar+1)
    mem[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  mem_MPORT_addr_pipe_0 = _RAND_5[25:0];
  _RAND_6 = {1{`RANDOM}};
  mem_MPORT_1_addr_pipe_0 = _RAND_6[25:0];
  _RAND_7 = {1{`RANDOM}};
  mem_MPORT_2_addr_pipe_0 = _RAND_7[25:0];
  _RAND_8 = {1{`RANDOM}};
  mem_MPORT_3_addr_pipe_0 = _RAND_8[25:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Triangle_memory(
  input         clock,
  input  [31:0] io_Triangle_id,
  output [31:0] io_v00_out,
  output [31:0] io_v11_out,
  output [31:0] io_v22_out
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg /* sparse */ [31:0] mem [0:51005099]; // @[Triangle_memory.scala 16:26]
  wire [31:0] mem_MPORT_data; // @[Triangle_memory.scala 16:26]
  wire [25:0] mem_MPORT_addr; // @[Triangle_memory.scala 16:26]
  wire [31:0] mem_MPORT_1_data; // @[Triangle_memory.scala 16:26]
  wire [25:0] mem_MPORT_1_addr; // @[Triangle_memory.scala 16:26]
  wire [31:0] mem_MPORT_2_data; // @[Triangle_memory.scala 16:26]
  wire [25:0] mem_MPORT_2_addr; // @[Triangle_memory.scala 16:26]
  wire [31:0] mem_MPORT_3_data; // @[Triangle_memory.scala 16:26]
  wire [25:0] mem_MPORT_3_addr; // @[Triangle_memory.scala 16:26]
  wire  mem_MPORT_3_mask; // @[Triangle_memory.scala 16:26]
  wire  mem_MPORT_3_en; // @[Triangle_memory.scala 16:26]
  reg [25:0] mem_MPORT_addr_pipe_0;
  reg [25:0] mem_MPORT_1_addr_pipe_0;
  reg [25:0] mem_MPORT_2_addr_pipe_0;
  wire [31:0] _T = io_Triangle_id; // @[Triangle_memory.scala 18:43]
  wire [31:0] _T_4 = io_Triangle_id + 32'h1; // @[Triangle_memory.scala 19:49]
  wire [31:0] _T_8 = io_Triangle_id + 32'h2; // @[Triangle_memory.scala 20:49]
  assign mem_MPORT_addr = mem_MPORT_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_data = mem[mem_MPORT_addr]; // @[Triangle_memory.scala 16:26]
  `else
  assign mem_MPORT_data = mem_MPORT_addr >= 26'h30a46ac ? _RAND_1[31:0] : mem[mem_MPORT_addr]; // @[Triangle_memory.scala 16:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_1_addr = mem_MPORT_1_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_1_data = mem[mem_MPORT_1_addr]; // @[Triangle_memory.scala 16:26]
  `else
  assign mem_MPORT_1_data = mem_MPORT_1_addr >= 26'h30a46ac ? _RAND_2[31:0] : mem[mem_MPORT_1_addr]; // @[Triangle_memory.scala 16:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_2_addr = mem_MPORT_2_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_2_data = mem[mem_MPORT_2_addr]; // @[Triangle_memory.scala 16:26]
  `else
  assign mem_MPORT_2_data = mem_MPORT_2_addr >= 26'h30a46ac ? _RAND_3[31:0] : mem[mem_MPORT_2_addr]; // @[Triangle_memory.scala 16:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_3_data = 32'h0;
  assign mem_MPORT_3_addr = 26'h0;
  assign mem_MPORT_3_mask = 1'h1;
  assign mem_MPORT_3_en = 1'h0;
  assign io_v00_out = mem_MPORT_data; // @[Triangle_memory.scala 18:16]
  assign io_v11_out = mem_MPORT_1_data; // @[Triangle_memory.scala 19:16]
  assign io_v22_out = mem_MPORT_2_data; // @[Triangle_memory.scala 20:16]
  always @(posedge clock) begin
    if(mem_MPORT_3_en & mem_MPORT_3_mask) begin
      mem[mem_MPORT_3_addr] <= mem_MPORT_3_data; // @[Triangle_memory.scala 16:26]
    end
    mem_MPORT_addr_pipe_0 <= _T[25:0];
    mem_MPORT_1_addr_pipe_0 <= _T_4[25:0];
    mem_MPORT_2_addr_pipe_0 <= _T_8[25:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {1{`RANDOM}};
  _RAND_2 = {1{`RANDOM}};
  _RAND_3 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 51005100; initvar = initvar+1)
    mem[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  mem_MPORT_addr_pipe_0 = _RAND_4[25:0];
  _RAND_5 = {1{`RANDOM}};
  mem_MPORT_1_addr_pipe_0 = _RAND_5[25:0];
  _RAND_6 = {1{`RANDOM}};
  mem_MPORT_2_addr_pipe_0 = _RAND_6[25:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MulAddRecFNToRaw_preMul(
  input  [32:0] io_a,
  input  [32:0] io_b,
  input  [32:0] io_c,
  output [23:0] io_mulAddA,
  output [23:0] io_mulAddB,
  output [47:0] io_mulAddC,
  output        io_toPostMul_isSigNaNAny,
  output        io_toPostMul_isNaNAOrB,
  output        io_toPostMul_isInfA,
  output        io_toPostMul_isZeroA,
  output        io_toPostMul_isInfB,
  output        io_toPostMul_isZeroB,
  output        io_toPostMul_signProd,
  output        io_toPostMul_isNaNC,
  output        io_toPostMul_isInfC,
  output        io_toPostMul_isZeroC,
  output [9:0]  io_toPostMul_sExpSum,
  output        io_toPostMul_doSubMags,
  output        io_toPostMul_CIsDominant,
  output [4:0]  io_toPostMul_CDom_CAlignDist,
  output [25:0] io_toPostMul_highAlignedSigC,
  output        io_toPostMul_bit0AlignedSigC
);
  wire  rawA_isZero = io_a[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_4 = io_a[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawA_isNaN = _T_4 & io_a[29]; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawA_sign = io_a[32]; // @[rawFloatFromRecFN.scala 58:25]
  wire [9:0] rawA_sExp = {1'b0,$signed(io_a[31:23])}; // @[rawFloatFromRecFN.scala 59:27]
  wire  hi_lo = ~rawA_isZero; // @[rawFloatFromRecFN.scala 60:39]
  wire [22:0] lo = io_a[22:0]; // @[rawFloatFromRecFN.scala 60:51]
  wire [24:0] rawA_sig = {1'h0,hi_lo,lo}; // @[Cat.scala 30:58]
  wire  rawB_isZero = io_b[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_17 = io_b[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawB_isNaN = _T_17 & io_b[29]; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawB_sign = io_b[32]; // @[rawFloatFromRecFN.scala 58:25]
  wire [9:0] rawB_sExp = {1'b0,$signed(io_b[31:23])}; // @[rawFloatFromRecFN.scala 59:27]
  wire  hi_lo_1 = ~rawB_isZero; // @[rawFloatFromRecFN.scala 60:39]
  wire [22:0] lo_1 = io_b[22:0]; // @[rawFloatFromRecFN.scala 60:51]
  wire [24:0] rawB_sig = {1'h0,hi_lo_1,lo_1}; // @[Cat.scala 30:58]
  wire  rawC_isZero = io_c[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_30 = io_c[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawC_isNaN = _T_30 & io_c[29]; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawC_sign = io_c[32]; // @[rawFloatFromRecFN.scala 58:25]
  wire [9:0] rawC_sExp = {1'b0,$signed(io_c[31:23])}; // @[rawFloatFromRecFN.scala 59:27]
  wire  hi_lo_2 = ~rawC_isZero; // @[rawFloatFromRecFN.scala 60:39]
  wire [22:0] lo_2 = io_c[22:0]; // @[rawFloatFromRecFN.scala 60:51]
  wire [24:0] rawC_sig = {1'h0,hi_lo_2,lo_2}; // @[Cat.scala 30:58]
  wire  signProd = rawA_sign ^ rawB_sign; // @[MulAddRecFN.scala 98:30]
  wire [10:0] _T_41 = $signed(rawA_sExp) + $signed(rawB_sExp); // @[MulAddRecFN.scala 101:19]
  wire [10:0] sExpAlignedProd = $signed(_T_41) - 11'she5; // @[MulAddRecFN.scala 101:32]
  wire  doSubMags = signProd ^ rawC_sign; // @[MulAddRecFN.scala 103:30]
  wire [10:0] _GEN_0 = {{1{rawC_sExp[9]}},rawC_sExp}; // @[MulAddRecFN.scala 107:42]
  wire [10:0] sNatCAlignDist = $signed(sExpAlignedProd) - $signed(_GEN_0); // @[MulAddRecFN.scala 107:42]
  wire [9:0] posNatCAlignDist = sNatCAlignDist[9:0]; // @[MulAddRecFN.scala 108:42]
  wire  isMinCAlign = rawA_isZero | rawB_isZero | $signed(sNatCAlignDist) < 11'sh0; // @[MulAddRecFN.scala 109:50]
  wire  CIsDominant = hi_lo_2 & (isMinCAlign | posNatCAlignDist <= 10'h18); // @[MulAddRecFN.scala 111:23]
  wire [6:0] _T_55 = posNatCAlignDist < 10'h4a ? posNatCAlignDist[6:0] : 7'h4a; // @[MulAddRecFN.scala 115:16]
  wire [6:0] CAlignDist = isMinCAlign ? 7'h0 : _T_55; // @[MulAddRecFN.scala 113:12]
  wire [24:0] _T_56 = ~rawC_sig; // @[MulAddRecFN.scala 121:28]
  wire [24:0] hi_3 = doSubMags ? _T_56 : rawC_sig; // @[MulAddRecFN.scala 121:16]
  wire [52:0] lo_3 = doSubMags ? 53'h1fffffffffffff : 53'h0; // @[Bitwise.scala 72:12]
  wire [77:0] _T_59 = {hi_3,lo_3}; // @[MulAddRecFN.scala 123:11]
  wire [77:0] mainAlignedSigC = $signed(_T_59) >>> CAlignDist; // @[MulAddRecFN.scala 123:17]
  wire [26:0] _T_60 = {rawC_sig, 2'h0}; // @[MulAddRecFN.scala 125:30]
  wire  _T_62 = |_T_60[3:0]; // @[primitives.scala 121:54]
  wire  _T_64 = |_T_60[7:4]; // @[primitives.scala 121:54]
  wire  _T_66 = |_T_60[11:8]; // @[primitives.scala 121:54]
  wire  _T_68 = |_T_60[15:12]; // @[primitives.scala 121:54]
  wire  _T_70 = |_T_60[19:16]; // @[primitives.scala 121:54]
  wire  _T_72 = |_T_60[23:20]; // @[primitives.scala 121:54]
  wire  _T_74 = |_T_60[26:24]; // @[primitives.scala 124:57]
  wire [6:0] _T_75 = {_T_74,_T_72,_T_70,_T_68,_T_66,_T_64,_T_62}; // @[primitives.scala 125:20]
  wire [32:0] _T_77 = 33'sh100000000 >>> CAlignDist[6:2]; // @[primitives.scala 77:58]
  wire  hi_5 = _T_77[14]; // @[Bitwise.scala 109:18]
  wire  lo_5 = _T_77[15]; // @[Bitwise.scala 109:44]
  wire  hi_7 = _T_77[16]; // @[Bitwise.scala 109:18]
  wire  lo_6 = _T_77[17]; // @[Bitwise.scala 109:44]
  wire  hi_9 = _T_77[18]; // @[Bitwise.scala 109:18]
  wire  lo_8 = _T_77[19]; // @[Bitwise.scala 109:44]
  wire [5:0] _T_83 = {hi_5,lo_5,hi_7,lo_6,hi_9,lo_8}; // @[Cat.scala 30:58]
  wire [6:0] _GEN_1 = {{1'd0}, _T_83}; // @[MulAddRecFN.scala 125:68]
  wire [6:0] _T_84 = _T_75 & _GEN_1; // @[MulAddRecFN.scala 125:68]
  wire  reduced4CExtra = |_T_84; // @[MulAddRecFN.scala 133:11]
  wire  _T_89 = &mainAlignedSigC[2:0] & ~reduced4CExtra; // @[MulAddRecFN.scala 137:44]
  wire  _T_92 = |mainAlignedSigC[2:0] | reduced4CExtra; // @[MulAddRecFN.scala 138:44]
  wire  lo_10 = doSubMags ? _T_89 : _T_92; // @[MulAddRecFN.scala 136:16]
  wire [74:0] hi_10 = mainAlignedSigC[77:3]; // @[Cat.scala 30:58]
  wire [75:0] alignedSigC = {hi_10,lo_10}; // @[Cat.scala 30:58]
  wire  _T_96 = rawA_isNaN & ~rawA_sig[22]; // @[common.scala 81:46]
  wire  _T_99 = rawB_isNaN & ~rawB_sig[22]; // @[common.scala 81:46]
  wire  _T_103 = rawC_isNaN & ~rawC_sig[22]; // @[common.scala 81:46]
  wire [10:0] _T_108 = $signed(sExpAlignedProd) - 11'sh18; // @[MulAddRecFN.scala 161:53]
  wire [10:0] _T_109 = CIsDominant ? $signed({{1{rawC_sExp[9]}},rawC_sExp}) : $signed(_T_108); // @[MulAddRecFN.scala 161:12]
  assign io_mulAddA = rawA_sig[23:0]; // @[MulAddRecFN.scala 144:16]
  assign io_mulAddB = rawB_sig[23:0]; // @[MulAddRecFN.scala 145:16]
  assign io_mulAddC = alignedSigC[48:1]; // @[MulAddRecFN.scala 146:30]
  assign io_toPostMul_isSigNaNAny = _T_96 | _T_99 | _T_103; // @[MulAddRecFN.scala 149:58]
  assign io_toPostMul_isNaNAOrB = rawA_isNaN | rawB_isNaN; // @[MulAddRecFN.scala 151:42]
  assign io_toPostMul_isInfA = _T_4 & ~io_a[29]; // @[rawFloatFromRecFN.scala 56:33]
  assign io_toPostMul_isZeroA = io_a[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign io_toPostMul_isInfB = _T_17 & ~io_b[29]; // @[rawFloatFromRecFN.scala 56:33]
  assign io_toPostMul_isZeroB = io_b[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign io_toPostMul_signProd = rawA_sign ^ rawB_sign; // @[MulAddRecFN.scala 98:30]
  assign io_toPostMul_isNaNC = _T_30 & io_c[29]; // @[rawFloatFromRecFN.scala 55:33]
  assign io_toPostMul_isInfC = _T_30 & ~io_c[29]; // @[rawFloatFromRecFN.scala 56:33]
  assign io_toPostMul_isZeroC = io_c[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign io_toPostMul_sExpSum = _T_109[9:0]; // @[MulAddRecFN.scala 160:28]
  assign io_toPostMul_doSubMags = signProd ^ rawC_sign; // @[MulAddRecFN.scala 103:30]
  assign io_toPostMul_CIsDominant = hi_lo_2 & (isMinCAlign | posNatCAlignDist <= 10'h18); // @[MulAddRecFN.scala 111:23]
  assign io_toPostMul_CDom_CAlignDist = CAlignDist[4:0]; // @[MulAddRecFN.scala 164:47]
  assign io_toPostMul_highAlignedSigC = alignedSigC[74:49]; // @[MulAddRecFN.scala 166:20]
  assign io_toPostMul_bit0AlignedSigC = alignedSigC[0]; // @[MulAddRecFN.scala 167:48]
endmodule
module MulAddRecFNToRaw_postMul(
  input         io_fromPreMul_isSigNaNAny,
  input         io_fromPreMul_isNaNAOrB,
  input         io_fromPreMul_isInfA,
  input         io_fromPreMul_isZeroA,
  input         io_fromPreMul_isInfB,
  input         io_fromPreMul_isZeroB,
  input         io_fromPreMul_signProd,
  input         io_fromPreMul_isNaNC,
  input         io_fromPreMul_isInfC,
  input         io_fromPreMul_isZeroC,
  input  [9:0]  io_fromPreMul_sExpSum,
  input         io_fromPreMul_doSubMags,
  input         io_fromPreMul_CIsDominant,
  input  [4:0]  io_fromPreMul_CDom_CAlignDist,
  input  [25:0] io_fromPreMul_highAlignedSigC,
  input         io_fromPreMul_bit0AlignedSigC,
  input  [48:0] io_mulAddResult,
  output        io_invalidExc,
  output        io_rawOut_isNaN,
  output        io_rawOut_isInf,
  output        io_rawOut_isZero,
  output        io_rawOut_sign,
  output [9:0]  io_rawOut_sExp,
  output [26:0] io_rawOut_sig
);
  wire  CDom_sign = io_fromPreMul_signProd ^ io_fromPreMul_doSubMags; // @[MulAddRecFN.scala 192:42]
  wire [25:0] _T_2 = io_fromPreMul_highAlignedSigC + 26'h1; // @[MulAddRecFN.scala 195:47]
  wire [25:0] hi_hi = io_mulAddResult[48] ? _T_2 : io_fromPreMul_highAlignedSigC; // @[MulAddRecFN.scala 194:16]
  wire [47:0] hi_lo = io_mulAddResult[47:0]; // @[MulAddRecFN.scala 198:28]
  wire [74:0] sigSum = {hi_hi,hi_lo,io_fromPreMul_bit0AlignedSigC}; // @[Cat.scala 30:58]
  wire [1:0] _T_3 = {1'b0,$signed(io_fromPreMul_doSubMags)}; // @[MulAddRecFN.scala 205:69]
  wire [9:0] _GEN_0 = {{8{_T_3[1]}},_T_3}; // @[MulAddRecFN.scala 205:43]
  wire [9:0] CDom_sExp = $signed(io_fromPreMul_sExpSum) - $signed(_GEN_0); // @[MulAddRecFN.scala 205:43]
  wire [49:0] _T_7 = ~sigSum[74:25]; // @[MulAddRecFN.scala 208:13]
  wire [1:0] hi_lo_1 = io_fromPreMul_highAlignedSigC[25:24]; // @[MulAddRecFN.scala 211:46]
  wire [46:0] lo = sigSum[72:26]; // @[MulAddRecFN.scala 212:23]
  wire [49:0] _T_8 = {1'h0,hi_lo_1,lo}; // @[Cat.scala 30:58]
  wire [49:0] CDom_absSigSum = io_fromPreMul_doSubMags ? _T_7 : _T_8; // @[MulAddRecFN.scala 207:12]
  wire [23:0] _T_10 = ~sigSum[24:1]; // @[MulAddRecFN.scala 217:14]
  wire  _T_11 = |_T_10; // @[MulAddRecFN.scala 217:36]
  wire  _T_13 = |sigSum[25:1]; // @[MulAddRecFN.scala 218:37]
  wire  CDom_absSigSumExtra = io_fromPreMul_doSubMags ? _T_11 : _T_13; // @[MulAddRecFN.scala 216:12]
  wire [80:0] _GEN_1 = {{31'd0}, CDom_absSigSum}; // @[MulAddRecFN.scala 221:24]
  wire [80:0] _T_14 = _GEN_1 << io_fromPreMul_CDom_CAlignDist; // @[MulAddRecFN.scala 221:24]
  wire [28:0] CDom_mainSig = _T_14[49:21]; // @[MulAddRecFN.scala 221:56]
  wire [26:0] _T_16 = {CDom_absSigSum[23:0], 3'h0}; // @[MulAddRecFN.scala 224:53]
  wire  _T_18 = |_T_16[3:0]; // @[primitives.scala 121:54]
  wire  _T_20 = |_T_16[7:4]; // @[primitives.scala 121:54]
  wire  _T_22 = |_T_16[11:8]; // @[primitives.scala 121:54]
  wire  _T_24 = |_T_16[15:12]; // @[primitives.scala 121:54]
  wire  _T_26 = |_T_16[19:16]; // @[primitives.scala 121:54]
  wire  _T_28 = |_T_16[23:20]; // @[primitives.scala 121:54]
  wire  _T_30 = |_T_16[26:24]; // @[primitives.scala 124:57]
  wire [6:0] _T_31 = {_T_30,_T_28,_T_26,_T_24,_T_22,_T_20,_T_18}; // @[primitives.scala 125:20]
  wire [2:0] _T_33 = ~io_fromPreMul_CDom_CAlignDist[4:2]; // @[primitives.scala 51:21]
  wire [8:0] _T_34 = 9'sh100 >>> _T_33; // @[primitives.scala 77:58]
  wire  hi_3 = _T_34[1]; // @[Bitwise.scala 109:18]
  wire  lo_2 = _T_34[2]; // @[Bitwise.scala 109:44]
  wire  hi_5 = _T_34[3]; // @[Bitwise.scala 109:18]
  wire  lo_3 = _T_34[4]; // @[Bitwise.scala 109:44]
  wire  hi_7 = _T_34[5]; // @[Bitwise.scala 109:18]
  wire  lo_5 = _T_34[6]; // @[Bitwise.scala 109:44]
  wire [5:0] _T_40 = {hi_3,lo_2,hi_5,lo_3,hi_7,lo_5}; // @[Cat.scala 30:58]
  wire [6:0] _GEN_2 = {{1'd0}, _T_40}; // @[MulAddRecFN.scala 224:72]
  wire [6:0] _T_41 = _T_31 & _GEN_2; // @[MulAddRecFN.scala 224:72]
  wire  CDom_reduced4SigExtra = |_T_41; // @[MulAddRecFN.scala 225:73]
  wire [25:0] hi_8 = CDom_mainSig[28:3]; // @[MulAddRecFN.scala 227:25]
  wire  lo_7 = |CDom_mainSig[2:0] | CDom_reduced4SigExtra | CDom_absSigSumExtra; // @[MulAddRecFN.scala 228:61]
  wire [26:0] CDom_sig = {hi_8,lo_7}; // @[Cat.scala 30:58]
  wire  notCDom_signSigSum = sigSum[51]; // @[MulAddRecFN.scala 234:36]
  wire [50:0] _T_46 = ~sigSum[50:0]; // @[MulAddRecFN.scala 237:13]
  wire [50:0] _GEN_3 = {{50'd0}, io_fromPreMul_doSubMags}; // @[MulAddRecFN.scala 238:41]
  wire [50:0] _T_49 = sigSum[50:0] + _GEN_3; // @[MulAddRecFN.scala 238:41]
  wire [50:0] notCDom_absSigSum = notCDom_signSigSum ? _T_46 : _T_49; // @[MulAddRecFN.scala 236:12]
  wire  _T_51 = |notCDom_absSigSum[1:0]; // @[primitives.scala 104:54]
  wire  _T_53 = |notCDom_absSigSum[3:2]; // @[primitives.scala 104:54]
  wire  _T_55 = |notCDom_absSigSum[5:4]; // @[primitives.scala 104:54]
  wire  _T_57 = |notCDom_absSigSum[7:6]; // @[primitives.scala 104:54]
  wire  _T_59 = |notCDom_absSigSum[9:8]; // @[primitives.scala 104:54]
  wire  _T_61 = |notCDom_absSigSum[11:10]; // @[primitives.scala 104:54]
  wire  _T_63 = |notCDom_absSigSum[13:12]; // @[primitives.scala 104:54]
  wire  _T_65 = |notCDom_absSigSum[15:14]; // @[primitives.scala 104:54]
  wire  _T_67 = |notCDom_absSigSum[17:16]; // @[primitives.scala 104:54]
  wire  _T_69 = |notCDom_absSigSum[19:18]; // @[primitives.scala 104:54]
  wire  _T_71 = |notCDom_absSigSum[21:20]; // @[primitives.scala 104:54]
  wire  _T_73 = |notCDom_absSigSum[23:22]; // @[primitives.scala 104:54]
  wire  _T_75 = |notCDom_absSigSum[25:24]; // @[primitives.scala 104:54]
  wire  _T_77 = |notCDom_absSigSum[27:26]; // @[primitives.scala 104:54]
  wire  _T_79 = |notCDom_absSigSum[29:28]; // @[primitives.scala 104:54]
  wire  _T_81 = |notCDom_absSigSum[31:30]; // @[primitives.scala 104:54]
  wire  _T_83 = |notCDom_absSigSum[33:32]; // @[primitives.scala 104:54]
  wire  _T_85 = |notCDom_absSigSum[35:34]; // @[primitives.scala 104:54]
  wire  _T_87 = |notCDom_absSigSum[37:36]; // @[primitives.scala 104:54]
  wire  _T_89 = |notCDom_absSigSum[39:38]; // @[primitives.scala 104:54]
  wire  _T_91 = |notCDom_absSigSum[41:40]; // @[primitives.scala 104:54]
  wire  _T_93 = |notCDom_absSigSum[43:42]; // @[primitives.scala 104:54]
  wire  _T_95 = |notCDom_absSigSum[45:44]; // @[primitives.scala 104:54]
  wire  _T_97 = |notCDom_absSigSum[47:46]; // @[primitives.scala 104:54]
  wire  _T_99 = |notCDom_absSigSum[49:48]; // @[primitives.scala 104:54]
  wire  _T_101 = |notCDom_absSigSum[50]; // @[primitives.scala 107:57]
  wire [5:0] lo_lo = {_T_61,_T_59,_T_57,_T_55,_T_53,_T_51}; // @[primitives.scala 108:20]
  wire [12:0] lo_8 = {_T_75,_T_73,_T_71,_T_69,_T_67,_T_65,_T_63,lo_lo}; // @[primitives.scala 108:20]
  wire [5:0] hi_lo_3 = {_T_87,_T_85,_T_83,_T_81,_T_79,_T_77}; // @[primitives.scala 108:20]
  wire [25:0] notCDom_reduced2AbsSigSum = {_T_101,_T_99,_T_97,_T_95,_T_93,_T_91,_T_89,hi_lo_3,lo_8}; // @[primitives.scala 108:20]
  wire [4:0] _T_128 = notCDom_reduced2AbsSigSum[1] ? 5'h18 : 5'h19; // @[Mux.scala 47:69]
  wire [4:0] _T_129 = notCDom_reduced2AbsSigSum[2] ? 5'h17 : _T_128; // @[Mux.scala 47:69]
  wire [4:0] _T_130 = notCDom_reduced2AbsSigSum[3] ? 5'h16 : _T_129; // @[Mux.scala 47:69]
  wire [4:0] _T_131 = notCDom_reduced2AbsSigSum[4] ? 5'h15 : _T_130; // @[Mux.scala 47:69]
  wire [4:0] _T_132 = notCDom_reduced2AbsSigSum[5] ? 5'h14 : _T_131; // @[Mux.scala 47:69]
  wire [4:0] _T_133 = notCDom_reduced2AbsSigSum[6] ? 5'h13 : _T_132; // @[Mux.scala 47:69]
  wire [4:0] _T_134 = notCDom_reduced2AbsSigSum[7] ? 5'h12 : _T_133; // @[Mux.scala 47:69]
  wire [4:0] _T_135 = notCDom_reduced2AbsSigSum[8] ? 5'h11 : _T_134; // @[Mux.scala 47:69]
  wire [4:0] _T_136 = notCDom_reduced2AbsSigSum[9] ? 5'h10 : _T_135; // @[Mux.scala 47:69]
  wire [4:0] _T_137 = notCDom_reduced2AbsSigSum[10] ? 5'hf : _T_136; // @[Mux.scala 47:69]
  wire [4:0] _T_138 = notCDom_reduced2AbsSigSum[11] ? 5'he : _T_137; // @[Mux.scala 47:69]
  wire [4:0] _T_139 = notCDom_reduced2AbsSigSum[12] ? 5'hd : _T_138; // @[Mux.scala 47:69]
  wire [4:0] _T_140 = notCDom_reduced2AbsSigSum[13] ? 5'hc : _T_139; // @[Mux.scala 47:69]
  wire [4:0] _T_141 = notCDom_reduced2AbsSigSum[14] ? 5'hb : _T_140; // @[Mux.scala 47:69]
  wire [4:0] _T_142 = notCDom_reduced2AbsSigSum[15] ? 5'ha : _T_141; // @[Mux.scala 47:69]
  wire [4:0] _T_143 = notCDom_reduced2AbsSigSum[16] ? 5'h9 : _T_142; // @[Mux.scala 47:69]
  wire [4:0] _T_144 = notCDom_reduced2AbsSigSum[17] ? 5'h8 : _T_143; // @[Mux.scala 47:69]
  wire [4:0] _T_145 = notCDom_reduced2AbsSigSum[18] ? 5'h7 : _T_144; // @[Mux.scala 47:69]
  wire [4:0] _T_146 = notCDom_reduced2AbsSigSum[19] ? 5'h6 : _T_145; // @[Mux.scala 47:69]
  wire [4:0] _T_147 = notCDom_reduced2AbsSigSum[20] ? 5'h5 : _T_146; // @[Mux.scala 47:69]
  wire [4:0] _T_148 = notCDom_reduced2AbsSigSum[21] ? 5'h4 : _T_147; // @[Mux.scala 47:69]
  wire [4:0] _T_149 = notCDom_reduced2AbsSigSum[22] ? 5'h3 : _T_148; // @[Mux.scala 47:69]
  wire [4:0] _T_150 = notCDom_reduced2AbsSigSum[23] ? 5'h2 : _T_149; // @[Mux.scala 47:69]
  wire [4:0] _T_151 = notCDom_reduced2AbsSigSum[24] ? 5'h1 : _T_150; // @[Mux.scala 47:69]
  wire [4:0] notCDom_normDistReduced2 = notCDom_reduced2AbsSigSum[25] ? 5'h0 : _T_151; // @[Mux.scala 47:69]
  wire [5:0] notCDom_nearNormDist = {notCDom_normDistReduced2, 1'h0}; // @[MulAddRecFN.scala 242:56]
  wire [6:0] _T_152 = {1'b0,$signed(notCDom_nearNormDist)}; // @[MulAddRecFN.scala 243:69]
  wire [9:0] _GEN_4 = {{3{_T_152[6]}},_T_152}; // @[MulAddRecFN.scala 243:46]
  wire [9:0] notCDom_sExp = $signed(io_fromPreMul_sExpSum) - $signed(_GEN_4); // @[MulAddRecFN.scala 243:46]
  wire [113:0] _GEN_5 = {{63'd0}, notCDom_absSigSum}; // @[MulAddRecFN.scala 245:27]
  wire [113:0] _T_155 = _GEN_5 << notCDom_nearNormDist; // @[MulAddRecFN.scala 245:27]
  wire [28:0] notCDom_mainSig = _T_155[51:23]; // @[MulAddRecFN.scala 245:50]
  wire  _T_159 = |notCDom_reduced2AbsSigSum[1:0]; // @[primitives.scala 104:54]
  wire  _T_161 = |notCDom_reduced2AbsSigSum[3:2]; // @[primitives.scala 104:54]
  wire  _T_163 = |notCDom_reduced2AbsSigSum[5:4]; // @[primitives.scala 104:54]
  wire  _T_165 = |notCDom_reduced2AbsSigSum[7:6]; // @[primitives.scala 104:54]
  wire  _T_167 = |notCDom_reduced2AbsSigSum[9:8]; // @[primitives.scala 104:54]
  wire  _T_169 = |notCDom_reduced2AbsSigSum[11:10]; // @[primitives.scala 104:54]
  wire  _T_171 = |notCDom_reduced2AbsSigSum[12]; // @[primitives.scala 107:57]
  wire [6:0] _T_172 = {_T_171,_T_169,_T_167,_T_165,_T_163,_T_161,_T_159}; // @[primitives.scala 108:20]
  wire [3:0] _T_174 = ~notCDom_normDistReduced2[4:1]; // @[primitives.scala 51:21]
  wire [16:0] _T_175 = 17'sh10000 >>> _T_174; // @[primitives.scala 77:58]
  wire  hi_11 = _T_175[1]; // @[Bitwise.scala 109:18]
  wire  lo_10 = _T_175[2]; // @[Bitwise.scala 109:44]
  wire  hi_13 = _T_175[3]; // @[Bitwise.scala 109:18]
  wire  lo_11 = _T_175[4]; // @[Bitwise.scala 109:44]
  wire  hi_15 = _T_175[5]; // @[Bitwise.scala 109:18]
  wire  lo_13 = _T_175[6]; // @[Bitwise.scala 109:44]
  wire [5:0] _T_181 = {hi_11,lo_10,hi_13,lo_11,hi_15,lo_13}; // @[Cat.scala 30:58]
  wire [6:0] _GEN_6 = {{1'd0}, _T_181}; // @[MulAddRecFN.scala 249:78]
  wire [6:0] _T_182 = _T_172 & _GEN_6; // @[MulAddRecFN.scala 249:78]
  wire  notCDom_reduced4SigExtra = |_T_182; // @[MulAddRecFN.scala 251:11]
  wire [25:0] hi_16 = notCDom_mainSig[28:3]; // @[MulAddRecFN.scala 253:28]
  wire  lo_15 = |notCDom_mainSig[2:0] | notCDom_reduced4SigExtra; // @[MulAddRecFN.scala 254:39]
  wire [26:0] notCDom_sig = {hi_16,lo_15}; // @[Cat.scala 30:58]
  wire  notCDom_completeCancellation = notCDom_sig[26:25] == 2'h0; // @[MulAddRecFN.scala 257:50]
  wire  _T_186 = io_fromPreMul_signProd ^ notCDom_signSigSum; // @[MulAddRecFN.scala 261:36]
  wire  notCDom_sign = notCDom_completeCancellation ? 1'h0 : _T_186; // @[MulAddRecFN.scala 259:12]
  wire  notNaN_isInfProd = io_fromPreMul_isInfA | io_fromPreMul_isInfB; // @[MulAddRecFN.scala 266:49]
  wire  notNaN_isInfOut = notNaN_isInfProd | io_fromPreMul_isInfC; // @[MulAddRecFN.scala 267:44]
  wire  notNaN_addZeros = (io_fromPreMul_isZeroA | io_fromPreMul_isZeroB) & io_fromPreMul_isZeroC; // @[MulAddRecFN.scala 269:58]
  wire  _T_188 = io_fromPreMul_isInfA & io_fromPreMul_isZeroB; // @[MulAddRecFN.scala 274:31]
  wire  _T_189 = io_fromPreMul_isSigNaNAny | _T_188; // @[MulAddRecFN.scala 273:35]
  wire  _T_190 = io_fromPreMul_isZeroA & io_fromPreMul_isInfB; // @[MulAddRecFN.scala 275:32]
  wire  _T_191 = _T_189 | _T_190; // @[MulAddRecFN.scala 274:57]
  wire  _T_194 = ~io_fromPreMul_isNaNAOrB & notNaN_isInfProd; // @[MulAddRecFN.scala 276:36]
  wire  _T_195 = _T_194 & io_fromPreMul_isInfC; // @[MulAddRecFN.scala 277:61]
  wire  _T_196 = _T_195 & io_fromPreMul_doSubMags; // @[MulAddRecFN.scala 278:35]
  wire  _T_200 = ~io_fromPreMul_CIsDominant & notCDom_completeCancellation; // @[MulAddRecFN.scala 285:42]
  wire  _T_203 = io_fromPreMul_isInfC & CDom_sign; // @[MulAddRecFN.scala 288:31]
  wire  _T_204 = notNaN_isInfProd & io_fromPreMul_signProd | _T_203; // @[MulAddRecFN.scala 287:54]
  wire  _T_207 = notNaN_addZeros & io_fromPreMul_signProd; // @[MulAddRecFN.scala 289:48]
  wire  _T_208 = _T_207 & CDom_sign; // @[MulAddRecFN.scala 290:36]
  wire  _T_209 = _T_204 | _T_208; // @[MulAddRecFN.scala 288:43]
  wire  _T_217 = io_fromPreMul_CIsDominant ? CDom_sign : notCDom_sign; // @[MulAddRecFN.scala 294:17]
  wire  _T_218 = ~notNaN_isInfOut & ~notNaN_addZeros & _T_217; // @[MulAddRecFN.scala 293:49]
  assign io_invalidExc = _T_191 | _T_196; // @[MulAddRecFN.scala 275:57]
  assign io_rawOut_isNaN = io_fromPreMul_isNaNAOrB | io_fromPreMul_isNaNC; // @[MulAddRecFN.scala 280:48]
  assign io_rawOut_isInf = notNaN_isInfProd | io_fromPreMul_isInfC; // @[MulAddRecFN.scala 267:44]
  assign io_rawOut_isZero = notNaN_addZeros | _T_200; // @[MulAddRecFN.scala 284:25]
  assign io_rawOut_sign = _T_209 | _T_218; // @[MulAddRecFN.scala 292:50]
  assign io_rawOut_sExp = io_fromPreMul_CIsDominant ? $signed(CDom_sExp) : $signed(notCDom_sExp); // @[MulAddRecFN.scala 295:26]
  assign io_rawOut_sig = io_fromPreMul_CIsDominant ? CDom_sig : notCDom_sig; // @[MulAddRecFN.scala 296:25]
endmodule
module RoundAnyRawFNToRecFN(
  input         io_invalidExc,
  input         io_in_isNaN,
  input         io_in_isInf,
  input         io_in_isZero,
  input         io_in_sign,
  input  [9:0]  io_in_sExp,
  input  [26:0] io_in_sig,
  output [32:0] io_out
);
  wire  doShiftSigDown1 = io_in_sig[26]; // @[RoundAnyRawFNToRecFN.scala 118:61]
  wire [8:0] _T_4 = ~io_in_sExp[8:0]; // @[primitives.scala 51:21]
  wire [64:0] _T_11 = 65'sh10000000000000000 >>> _T_4[5:0]; // @[primitives.scala 77:58]
  wire [15:0] _T_17 = {{8'd0}, _T_11[57:50]}; // @[Bitwise.scala 103:31]
  wire [15:0] _T_19 = {_T_11[49:42], 8'h0}; // @[Bitwise.scala 103:65]
  wire [15:0] _T_21 = _T_19 & 16'hff00; // @[Bitwise.scala 103:75]
  wire [15:0] _T_22 = _T_17 | _T_21; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_0 = {{4'd0}, _T_22[15:4]}; // @[Bitwise.scala 103:31]
  wire [15:0] _T_27 = _GEN_0 & 16'hf0f; // @[Bitwise.scala 103:31]
  wire [15:0] _T_29 = {_T_22[11:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [15:0] _T_31 = _T_29 & 16'hf0f0; // @[Bitwise.scala 103:75]
  wire [15:0] _T_32 = _T_27 | _T_31; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_1 = {{2'd0}, _T_32[15:2]}; // @[Bitwise.scala 103:31]
  wire [15:0] _T_37 = _GEN_1 & 16'h3333; // @[Bitwise.scala 103:31]
  wire [15:0] _T_39 = {_T_32[13:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [15:0] _T_41 = _T_39 & 16'hcccc; // @[Bitwise.scala 103:75]
  wire [15:0] _T_42 = _T_37 | _T_41; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_2 = {{1'd0}, _T_42[15:1]}; // @[Bitwise.scala 103:31]
  wire [15:0] _T_47 = _GEN_2 & 16'h5555; // @[Bitwise.scala 103:31]
  wire [15:0] _T_49 = {_T_42[14:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [15:0] _T_51 = _T_49 & 16'haaaa; // @[Bitwise.scala 103:75]
  wire [15:0] hi = _T_47 | _T_51; // @[Bitwise.scala 103:39]
  wire  hi_1 = _T_11[58]; // @[Bitwise.scala 109:18]
  wire  lo = _T_11[59]; // @[Bitwise.scala 109:44]
  wire  hi_3 = _T_11[60]; // @[Bitwise.scala 109:18]
  wire  lo_1 = _T_11[61]; // @[Bitwise.scala 109:44]
  wire  hi_5 = _T_11[62]; // @[Bitwise.scala 109:18]
  wire  lo_3 = _T_11[63]; // @[Bitwise.scala 109:44]
  wire [21:0] _T_57 = {hi,hi_1,lo,hi_3,lo_1,hi_5,lo_3}; // @[Cat.scala 30:58]
  wire [21:0] _T_58 = ~_T_57; // @[primitives.scala 74:36]
  wire [21:0] _T_59 = _T_4[6] ? 22'h0 : _T_58; // @[primitives.scala 74:21]
  wire [21:0] hi_6 = ~_T_59; // @[primitives.scala 74:17]
  wire [24:0] _T_60 = {hi_6,3'h7}; // @[Cat.scala 30:58]
  wire  hi_7 = _T_11[0]; // @[Bitwise.scala 109:18]
  wire  lo_6 = _T_11[1]; // @[Bitwise.scala 109:44]
  wire  lo_7 = _T_11[2]; // @[Bitwise.scala 109:44]
  wire [2:0] _T_66 = {hi_7,lo_6,lo_7}; // @[Cat.scala 30:58]
  wire [2:0] _T_67 = _T_4[6] ? _T_66 : 3'h0; // @[primitives.scala 61:24]
  wire [24:0] _T_68 = _T_4[7] ? _T_60 : {{22'd0}, _T_67}; // @[primitives.scala 66:24]
  wire [24:0] _T_69 = _T_4[8] ? _T_68 : 25'h0; // @[primitives.scala 61:24]
  wire [24:0] _GEN_3 = {{24'd0}, doShiftSigDown1}; // @[RoundAnyRawFNToRecFN.scala 157:23]
  wire [24:0] hi_9 = _T_69 | _GEN_3; // @[RoundAnyRawFNToRecFN.scala 157:23]
  wire [26:0] _T_70 = {hi_9,2'h3}; // @[Cat.scala 30:58]
  wire [25:0] lo_8 = _T_70[26:1]; // @[RoundAnyRawFNToRecFN.scala 160:57]
  wire [26:0] _T_71 = {1'h0,lo_8}; // @[Cat.scala 30:58]
  wire [26:0] _T_72 = ~_T_71; // @[RoundAnyRawFNToRecFN.scala 161:28]
  wire [26:0] _T_73 = _T_72 & _T_70; // @[RoundAnyRawFNToRecFN.scala 161:46]
  wire [26:0] _T_74 = io_in_sig & _T_73; // @[RoundAnyRawFNToRecFN.scala 162:40]
  wire  _T_75 = |_T_74; // @[RoundAnyRawFNToRecFN.scala 162:56]
  wire [26:0] _T_76 = io_in_sig & _T_71; // @[RoundAnyRawFNToRecFN.scala 163:42]
  wire  _T_77 = |_T_76; // @[RoundAnyRawFNToRecFN.scala 163:62]
  wire [26:0] _T_83 = io_in_sig | _T_70; // @[RoundAnyRawFNToRecFN.scala 172:32]
  wire [25:0] _T_85 = _T_83[26:2] + 25'h1; // @[RoundAnyRawFNToRecFN.scala 172:49]
  wire  _T_87 = ~_T_77; // @[RoundAnyRawFNToRecFN.scala 174:30]
  wire [25:0] _T_90 = _T_75 & _T_87 ? lo_8 : 26'h0; // @[RoundAnyRawFNToRecFN.scala 173:25]
  wire [25:0] _T_91 = ~_T_90; // @[RoundAnyRawFNToRecFN.scala 173:21]
  wire [25:0] _T_92 = _T_85 & _T_91; // @[RoundAnyRawFNToRecFN.scala 172:61]
  wire [26:0] _T_93 = ~_T_70; // @[RoundAnyRawFNToRecFN.scala 178:32]
  wire [26:0] _T_94 = io_in_sig & _T_93; // @[RoundAnyRawFNToRecFN.scala 178:30]
  wire [25:0] _T_99 = {{1'd0}, _T_94[26:2]}; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [25:0] _T_100 = _T_75 ? _T_92 : _T_99; // @[RoundAnyRawFNToRecFN.scala 171:16]
  wire [2:0] _T_102 = {1'b0,$signed(_T_100[25:24])}; // @[RoundAnyRawFNToRecFN.scala 183:69]
  wire [9:0] _GEN_4 = {{7{_T_102[2]}},_T_102}; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [10:0] _T_103 = $signed(io_in_sExp) + $signed(_GEN_4); // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [8:0] common_expOut = _T_103[8:0]; // @[RoundAnyRawFNToRecFN.scala 185:37]
  wire [22:0] common_fractOut = doShiftSigDown1 ? _T_100[23:1] : _T_100[22:0]; // @[RoundAnyRawFNToRecFN.scala 187:16]
  wire [3:0] _T_108 = _T_103[10:7]; // @[RoundAnyRawFNToRecFN.scala 194:30]
  wire  common_overflow = $signed(_T_108) >= 4'sh3; // @[RoundAnyRawFNToRecFN.scala 194:50]
  wire  common_totalUnderflow = $signed(_T_103) < 11'sh6b; // @[RoundAnyRawFNToRecFN.scala 198:31]
  wire  isNaNOut = io_invalidExc | io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 233:34]
  wire  commonCase = ~isNaNOut & ~io_in_isInf & ~io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 235:61]
  wire  overflow = commonCase & common_overflow; // @[RoundAnyRawFNToRecFN.scala 236:32]
  wire  notNaN_isInfOut = io_in_isInf | overflow; // @[RoundAnyRawFNToRecFN.scala 246:32]
  wire  signOut = isNaNOut ? 1'h0 : io_in_sign; // @[RoundAnyRawFNToRecFN.scala 248:22]
  wire [8:0] _T_157 = io_in_isZero | common_totalUnderflow ? 9'h1c0 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 251:18]
  wire [8:0] _T_158 = ~_T_157; // @[RoundAnyRawFNToRecFN.scala 251:14]
  wire [8:0] _T_159 = common_expOut & _T_158; // @[RoundAnyRawFNToRecFN.scala 250:24]
  wire [8:0] _T_167 = notNaN_isInfOut ? 9'h40 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 263:18]
  wire [8:0] _T_168 = ~_T_167; // @[RoundAnyRawFNToRecFN.scala 263:14]
  wire [8:0] _T_169 = _T_159 & _T_168; // @[RoundAnyRawFNToRecFN.scala 262:17]
  wire [8:0] _T_174 = notNaN_isInfOut ? 9'h180 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 275:16]
  wire [8:0] _T_175 = _T_169 | _T_174; // @[RoundAnyRawFNToRecFN.scala 274:15]
  wire [8:0] _T_176 = isNaNOut ? 9'h1c0 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 276:16]
  wire [8:0] expOut = _T_175 | _T_176; // @[RoundAnyRawFNToRecFN.scala 275:77]
  wire [22:0] _T_179 = isNaNOut ? 23'h400000 : 23'h0; // @[RoundAnyRawFNToRecFN.scala 279:16]
  wire [22:0] fractOut = isNaNOut | io_in_isZero | common_totalUnderflow ? _T_179 : common_fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12]
  wire [9:0] hi_10 = {signOut,expOut}; // @[Cat.scala 30:58]
  assign io_out = {hi_10,fractOut}; // @[Cat.scala 30:58]
endmodule
module RoundRawFNToRecFN(
  input         io_invalidExc,
  input         io_in_isNaN,
  input         io_in_isInf,
  input         io_in_isZero,
  input         io_in_sign,
  input  [9:0]  io_in_sExp,
  input  [26:0] io_in_sig,
  output [32:0] io_out
);
  wire  roundAnyRawFNToRecFN_io_invalidExc; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_sign; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [9:0] roundAnyRawFNToRecFN_io_in_sExp; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [26:0] roundAnyRawFNToRecFN_io_in_sig; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [32:0] roundAnyRawFNToRecFN_io_out; // @[RoundAnyRawFNToRecFN.scala 307:15]
  RoundAnyRawFNToRecFN roundAnyRawFNToRecFN ( // @[RoundAnyRawFNToRecFN.scala 307:15]
    .io_invalidExc(roundAnyRawFNToRecFN_io_invalidExc),
    .io_in_isNaN(roundAnyRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundAnyRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundAnyRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundAnyRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundAnyRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundAnyRawFNToRecFN_io_in_sig),
    .io_out(roundAnyRawFNToRecFN_io_out)
  );
  assign io_out = roundAnyRawFNToRecFN_io_out; // @[RoundAnyRawFNToRecFN.scala 315:23]
  assign roundAnyRawFNToRecFN_io_invalidExc = io_invalidExc; // @[RoundAnyRawFNToRecFN.scala 310:44]
  assign roundAnyRawFNToRecFN_io_in_isNaN = io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_isInf = io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_isZero = io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_sign = io_in_sign; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_sExp = io_in_sExp; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_sig = io_in_sig; // @[RoundAnyRawFNToRecFN.scala 312:44]
endmodule
module MY_MULADD(
  input         clock,
  input         reset,
  input  [31:0] io_a,
  input  [31:0] io_b,
  input  [31:0] io_c,
  output [31:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_REG_INIT
  wire [32:0] mulAddRecFNToRaw_preMul_io_a; // @[FMULADD_1G_2.scala 36:15]
  wire [32:0] mulAddRecFNToRaw_preMul_io_b; // @[FMULADD_1G_2.scala 36:15]
  wire [32:0] mulAddRecFNToRaw_preMul_io_c; // @[FMULADD_1G_2.scala 36:15]
  wire [23:0] mulAddRecFNToRaw_preMul_io_mulAddA; // @[FMULADD_1G_2.scala 36:15]
  wire [23:0] mulAddRecFNToRaw_preMul_io_mulAddB; // @[FMULADD_1G_2.scala 36:15]
  wire [47:0] mulAddRecFNToRaw_preMul_io_mulAddC; // @[FMULADD_1G_2.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny; // @[FMULADD_1G_2.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB; // @[FMULADD_1G_2.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfA; // @[FMULADD_1G_2.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA; // @[FMULADD_1G_2.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfB; // @[FMULADD_1G_2.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB; // @[FMULADD_1G_2.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_signProd; // @[FMULADD_1G_2.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC; // @[FMULADD_1G_2.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfC; // @[FMULADD_1G_2.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC; // @[FMULADD_1G_2.scala 36:15]
  wire [9:0] mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum; // @[FMULADD_1G_2.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags; // @[FMULADD_1G_2.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant; // @[FMULADD_1G_2.scala 36:15]
  wire [4:0] mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist; // @[FMULADD_1G_2.scala 36:15]
  wire [25:0] mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC; // @[FMULADD_1G_2.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC; // @[FMULADD_1G_2.scala 36:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny; // @[FMULADD_1G_2.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB; // @[FMULADD_1G_2.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA; // @[FMULADD_1G_2.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA; // @[FMULADD_1G_2.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB; // @[FMULADD_1G_2.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB; // @[FMULADD_1G_2.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_signProd; // @[FMULADD_1G_2.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC; // @[FMULADD_1G_2.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC; // @[FMULADD_1G_2.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC; // @[FMULADD_1G_2.scala 116:15]
  wire [9:0] mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum; // @[FMULADD_1G_2.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags; // @[FMULADD_1G_2.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant; // @[FMULADD_1G_2.scala 116:15]
  wire [4:0] mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist; // @[FMULADD_1G_2.scala 116:15]
  wire [25:0] mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC; // @[FMULADD_1G_2.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC; // @[FMULADD_1G_2.scala 116:15]
  wire [48:0] mulAddRecFNToRaw_postMul_io_mulAddResult; // @[FMULADD_1G_2.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_invalidExc; // @[FMULADD_1G_2.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isNaN; // @[FMULADD_1G_2.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isInf; // @[FMULADD_1G_2.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isZero; // @[FMULADD_1G_2.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_sign; // @[FMULADD_1G_2.scala 116:15]
  wire [9:0] mulAddRecFNToRaw_postMul_io_rawOut_sExp; // @[FMULADD_1G_2.scala 116:15]
  wire [26:0] mulAddRecFNToRaw_postMul_io_rawOut_sig; // @[FMULADD_1G_2.scala 116:15]
  wire  roundRawFNToRecFN_io_invalidExc; // @[FMULADD_1G_2.scala 137:15]
  wire  roundRawFNToRecFN_io_in_isNaN; // @[FMULADD_1G_2.scala 137:15]
  wire  roundRawFNToRecFN_io_in_isInf; // @[FMULADD_1G_2.scala 137:15]
  wire  roundRawFNToRecFN_io_in_isZero; // @[FMULADD_1G_2.scala 137:15]
  wire  roundRawFNToRecFN_io_in_sign; // @[FMULADD_1G_2.scala 137:15]
  wire [9:0] roundRawFNToRecFN_io_in_sExp; // @[FMULADD_1G_2.scala 137:15]
  wire [26:0] roundRawFNToRecFN_io_in_sig; // @[FMULADD_1G_2.scala 137:15]
  wire [32:0] roundRawFNToRecFN_io_out; // @[FMULADD_1G_2.scala 137:15]
  reg [23:0] premul_a; // @[FMULADD_1G_2.scala 15:37]
  reg [23:0] premul_b; // @[FMULADD_1G_2.scala 16:37]
  reg [47:0] premul_c; // @[FMULADD_1G_2.scala 17:37]
  reg  isSigNaNAny; // @[FMULADD_1G_2.scala 18:33]
  reg  isNaNAOrB; // @[FMULADD_1G_2.scala 19:34]
  reg  isInfA; // @[FMULADD_1G_2.scala 20:43]
  reg  isZeroA; // @[FMULADD_1G_2.scala 21:40]
  reg  isInfB; // @[FMULADD_1G_2.scala 22:43]
  reg  isZeroB; // @[FMULADD_1G_2.scala 23:40]
  reg  signProd; // @[FMULADD_1G_2.scala 24:38]
  reg  isNaNC; // @[FMULADD_1G_2.scala 25:39]
  reg  isInfC; // @[FMULADD_1G_2.scala 26:42]
  reg  isZeroC; // @[FMULADD_1G_2.scala 27:39]
  reg [9:0] sExpSum; // @[FMULADD_1G_2.scala 28:36]
  reg  doSubMags; // @[FMULADD_1G_2.scala 29:33]
  reg  CIsDominant; // @[FMULADD_1G_2.scala 30:33]
  reg [4:0] CDom_CAlignDist; // @[FMULADD_1G_2.scala 31:34]
  reg [25:0] highAlignedSigC; // @[FMULADD_1G_2.scala 32:37]
  reg  bit0AlignedSigC; // @[FMULADD_1G_2.scala 33:38]
  wire  _T_3 = io_a[30:23] == 8'h0; // @[rawFloatFromFN.scala 50:34]
  wire  _T_4 = io_a[22:0] == 23'h0; // @[rawFloatFromFN.scala 51:38]
  wire [4:0] _T_28 = io_a[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:69]
  wire [4:0] _T_29 = io_a[2] ? 5'h14 : _T_28; // @[Mux.scala 47:69]
  wire [4:0] _T_30 = io_a[3] ? 5'h13 : _T_29; // @[Mux.scala 47:69]
  wire [4:0] _T_31 = io_a[4] ? 5'h12 : _T_30; // @[Mux.scala 47:69]
  wire [4:0] _T_32 = io_a[5] ? 5'h11 : _T_31; // @[Mux.scala 47:69]
  wire [4:0] _T_33 = io_a[6] ? 5'h10 : _T_32; // @[Mux.scala 47:69]
  wire [4:0] _T_34 = io_a[7] ? 5'hf : _T_33; // @[Mux.scala 47:69]
  wire [4:0] _T_35 = io_a[8] ? 5'he : _T_34; // @[Mux.scala 47:69]
  wire [4:0] _T_36 = io_a[9] ? 5'hd : _T_35; // @[Mux.scala 47:69]
  wire [4:0] _T_37 = io_a[10] ? 5'hc : _T_36; // @[Mux.scala 47:69]
  wire [4:0] _T_38 = io_a[11] ? 5'hb : _T_37; // @[Mux.scala 47:69]
  wire [4:0] _T_39 = io_a[12] ? 5'ha : _T_38; // @[Mux.scala 47:69]
  wire [4:0] _T_40 = io_a[13] ? 5'h9 : _T_39; // @[Mux.scala 47:69]
  wire [4:0] _T_41 = io_a[14] ? 5'h8 : _T_40; // @[Mux.scala 47:69]
  wire [4:0] _T_42 = io_a[15] ? 5'h7 : _T_41; // @[Mux.scala 47:69]
  wire [4:0] _T_43 = io_a[16] ? 5'h6 : _T_42; // @[Mux.scala 47:69]
  wire [4:0] _T_44 = io_a[17] ? 5'h5 : _T_43; // @[Mux.scala 47:69]
  wire [4:0] _T_45 = io_a[18] ? 5'h4 : _T_44; // @[Mux.scala 47:69]
  wire [4:0] _T_46 = io_a[19] ? 5'h3 : _T_45; // @[Mux.scala 47:69]
  wire [4:0] _T_47 = io_a[20] ? 5'h2 : _T_46; // @[Mux.scala 47:69]
  wire [4:0] _T_48 = io_a[21] ? 5'h1 : _T_47; // @[Mux.scala 47:69]
  wire [4:0] _T_49 = io_a[22] ? 5'h0 : _T_48; // @[Mux.scala 47:69]
  wire [53:0] _GEN_0 = {{31'd0}, io_a[22:0]}; // @[rawFloatFromFN.scala 54:36]
  wire [53:0] _T_50 = _GEN_0 << _T_49; // @[rawFloatFromFN.scala 54:36]
  wire [22:0] _T_52 = {_T_50[21:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  wire [8:0] _GEN_1 = {{4'd0}, _T_49}; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_53 = _GEN_1 ^ 9'h1ff; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_54 = _T_3 ? _T_53 : {{1'd0}, io_a[30:23]}; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_55 = _T_3 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  wire [7:0] _GEN_2 = {{6'd0}, _T_55}; // @[rawFloatFromFN.scala 60:22]
  wire [7:0] _T_56 = 8'h80 | _GEN_2; // @[rawFloatFromFN.scala 60:22]
  wire [8:0] _GEN_3 = {{1'd0}, _T_56}; // @[rawFloatFromFN.scala 59:15]
  wire [8:0] _T_58 = _T_54 + _GEN_3; // @[rawFloatFromFN.scala 59:15]
  wire  _T_59 = _T_3 & _T_4; // @[rawFloatFromFN.scala 62:34]
  wire  _T_61 = _T_58[8:7] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  wire  _T_63 = _T_61 & ~_T_4; // @[rawFloatFromFN.scala 66:33]
  wire [9:0] _T_66 = {1'b0,$signed(_T_58)}; // @[rawFloatFromFN.scala 70:48]
  wire  hi_lo = ~_T_59; // @[rawFloatFromFN.scala 72:29]
  wire [22:0] lo = _T_3 ? _T_52 : io_a[22:0]; // @[rawFloatFromFN.scala 72:42]
  wire [24:0] _T_67 = {1'h0,hi_lo,lo}; // @[Cat.scala 30:58]
  wire [2:0] _T_69 = _T_59 ? 3'h0 : _T_66[8:6]; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_4 = {{2'd0}, _T_63}; // @[recFNFromFN.scala 48:79]
  wire [2:0] hi_lo_1 = _T_69 | _GEN_4; // @[recFNFromFN.scala 48:79]
  wire [5:0] lo_hi = _T_66[5:0]; // @[recFNFromFN.scala 50:23]
  wire [22:0] lo_lo = _T_67[22:0]; // @[recFNFromFN.scala 51:22]
  wire [28:0] lo_1 = {lo_hi,lo_lo}; // @[Cat.scala 30:58]
  wire [3:0] hi_1 = {io_a[31],hi_lo_1}; // @[Cat.scala 30:58]
  wire  _T_75 = io_b[30:23] == 8'h0; // @[rawFloatFromFN.scala 50:34]
  wire  _T_76 = io_b[22:0] == 23'h0; // @[rawFloatFromFN.scala 51:38]
  wire [4:0] _T_100 = io_b[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:69]
  wire [4:0] _T_101 = io_b[2] ? 5'h14 : _T_100; // @[Mux.scala 47:69]
  wire [4:0] _T_102 = io_b[3] ? 5'h13 : _T_101; // @[Mux.scala 47:69]
  wire [4:0] _T_103 = io_b[4] ? 5'h12 : _T_102; // @[Mux.scala 47:69]
  wire [4:0] _T_104 = io_b[5] ? 5'h11 : _T_103; // @[Mux.scala 47:69]
  wire [4:0] _T_105 = io_b[6] ? 5'h10 : _T_104; // @[Mux.scala 47:69]
  wire [4:0] _T_106 = io_b[7] ? 5'hf : _T_105; // @[Mux.scala 47:69]
  wire [4:0] _T_107 = io_b[8] ? 5'he : _T_106; // @[Mux.scala 47:69]
  wire [4:0] _T_108 = io_b[9] ? 5'hd : _T_107; // @[Mux.scala 47:69]
  wire [4:0] _T_109 = io_b[10] ? 5'hc : _T_108; // @[Mux.scala 47:69]
  wire [4:0] _T_110 = io_b[11] ? 5'hb : _T_109; // @[Mux.scala 47:69]
  wire [4:0] _T_111 = io_b[12] ? 5'ha : _T_110; // @[Mux.scala 47:69]
  wire [4:0] _T_112 = io_b[13] ? 5'h9 : _T_111; // @[Mux.scala 47:69]
  wire [4:0] _T_113 = io_b[14] ? 5'h8 : _T_112; // @[Mux.scala 47:69]
  wire [4:0] _T_114 = io_b[15] ? 5'h7 : _T_113; // @[Mux.scala 47:69]
  wire [4:0] _T_115 = io_b[16] ? 5'h6 : _T_114; // @[Mux.scala 47:69]
  wire [4:0] _T_116 = io_b[17] ? 5'h5 : _T_115; // @[Mux.scala 47:69]
  wire [4:0] _T_117 = io_b[18] ? 5'h4 : _T_116; // @[Mux.scala 47:69]
  wire [4:0] _T_118 = io_b[19] ? 5'h3 : _T_117; // @[Mux.scala 47:69]
  wire [4:0] _T_119 = io_b[20] ? 5'h2 : _T_118; // @[Mux.scala 47:69]
  wire [4:0] _T_120 = io_b[21] ? 5'h1 : _T_119; // @[Mux.scala 47:69]
  wire [4:0] _T_121 = io_b[22] ? 5'h0 : _T_120; // @[Mux.scala 47:69]
  wire [53:0] _GEN_5 = {{31'd0}, io_b[22:0]}; // @[rawFloatFromFN.scala 54:36]
  wire [53:0] _T_122 = _GEN_5 << _T_121; // @[rawFloatFromFN.scala 54:36]
  wire [22:0] _T_124 = {_T_122[21:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  wire [8:0] _GEN_6 = {{4'd0}, _T_121}; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_125 = _GEN_6 ^ 9'h1ff; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_126 = _T_75 ? _T_125 : {{1'd0}, io_b[30:23]}; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_127 = _T_75 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  wire [7:0] _GEN_7 = {{6'd0}, _T_127}; // @[rawFloatFromFN.scala 60:22]
  wire [7:0] _T_128 = 8'h80 | _GEN_7; // @[rawFloatFromFN.scala 60:22]
  wire [8:0] _GEN_8 = {{1'd0}, _T_128}; // @[rawFloatFromFN.scala 59:15]
  wire [8:0] _T_130 = _T_126 + _GEN_8; // @[rawFloatFromFN.scala 59:15]
  wire  _T_131 = _T_75 & _T_76; // @[rawFloatFromFN.scala 62:34]
  wire  _T_133 = _T_130[8:7] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  wire  _T_135 = _T_133 & ~_T_76; // @[rawFloatFromFN.scala 66:33]
  wire [9:0] _T_138 = {1'b0,$signed(_T_130)}; // @[rawFloatFromFN.scala 70:48]
  wire  hi_lo_2 = ~_T_131; // @[rawFloatFromFN.scala 72:29]
  wire [22:0] lo_2 = _T_75 ? _T_124 : io_b[22:0]; // @[rawFloatFromFN.scala 72:42]
  wire [24:0] _T_139 = {1'h0,hi_lo_2,lo_2}; // @[Cat.scala 30:58]
  wire [2:0] _T_141 = _T_131 ? 3'h0 : _T_138[8:6]; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_9 = {{2'd0}, _T_135}; // @[recFNFromFN.scala 48:79]
  wire [2:0] hi_lo_3 = _T_141 | _GEN_9; // @[recFNFromFN.scala 48:79]
  wire [5:0] lo_hi_1 = _T_138[5:0]; // @[recFNFromFN.scala 50:23]
  wire [22:0] lo_lo_1 = _T_139[22:0]; // @[recFNFromFN.scala 51:22]
  wire [28:0] lo_3 = {lo_hi_1,lo_lo_1}; // @[Cat.scala 30:58]
  wire [3:0] hi_3 = {io_b[31],hi_lo_3}; // @[Cat.scala 30:58]
  wire  _T_147 = io_c[30:23] == 8'h0; // @[rawFloatFromFN.scala 50:34]
  wire  _T_148 = io_c[22:0] == 23'h0; // @[rawFloatFromFN.scala 51:38]
  wire [4:0] _T_172 = io_c[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:69]
  wire [4:0] _T_173 = io_c[2] ? 5'h14 : _T_172; // @[Mux.scala 47:69]
  wire [4:0] _T_174 = io_c[3] ? 5'h13 : _T_173; // @[Mux.scala 47:69]
  wire [4:0] _T_175 = io_c[4] ? 5'h12 : _T_174; // @[Mux.scala 47:69]
  wire [4:0] _T_176 = io_c[5] ? 5'h11 : _T_175; // @[Mux.scala 47:69]
  wire [4:0] _T_177 = io_c[6] ? 5'h10 : _T_176; // @[Mux.scala 47:69]
  wire [4:0] _T_178 = io_c[7] ? 5'hf : _T_177; // @[Mux.scala 47:69]
  wire [4:0] _T_179 = io_c[8] ? 5'he : _T_178; // @[Mux.scala 47:69]
  wire [4:0] _T_180 = io_c[9] ? 5'hd : _T_179; // @[Mux.scala 47:69]
  wire [4:0] _T_181 = io_c[10] ? 5'hc : _T_180; // @[Mux.scala 47:69]
  wire [4:0] _T_182 = io_c[11] ? 5'hb : _T_181; // @[Mux.scala 47:69]
  wire [4:0] _T_183 = io_c[12] ? 5'ha : _T_182; // @[Mux.scala 47:69]
  wire [4:0] _T_184 = io_c[13] ? 5'h9 : _T_183; // @[Mux.scala 47:69]
  wire [4:0] _T_185 = io_c[14] ? 5'h8 : _T_184; // @[Mux.scala 47:69]
  wire [4:0] _T_186 = io_c[15] ? 5'h7 : _T_185; // @[Mux.scala 47:69]
  wire [4:0] _T_187 = io_c[16] ? 5'h6 : _T_186; // @[Mux.scala 47:69]
  wire [4:0] _T_188 = io_c[17] ? 5'h5 : _T_187; // @[Mux.scala 47:69]
  wire [4:0] _T_189 = io_c[18] ? 5'h4 : _T_188; // @[Mux.scala 47:69]
  wire [4:0] _T_190 = io_c[19] ? 5'h3 : _T_189; // @[Mux.scala 47:69]
  wire [4:0] _T_191 = io_c[20] ? 5'h2 : _T_190; // @[Mux.scala 47:69]
  wire [4:0] _T_192 = io_c[21] ? 5'h1 : _T_191; // @[Mux.scala 47:69]
  wire [4:0] _T_193 = io_c[22] ? 5'h0 : _T_192; // @[Mux.scala 47:69]
  wire [53:0] _GEN_10 = {{31'd0}, io_c[22:0]}; // @[rawFloatFromFN.scala 54:36]
  wire [53:0] _T_194 = _GEN_10 << _T_193; // @[rawFloatFromFN.scala 54:36]
  wire [22:0] _T_196 = {_T_194[21:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  wire [8:0] _GEN_11 = {{4'd0}, _T_193}; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_197 = _GEN_11 ^ 9'h1ff; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_198 = _T_147 ? _T_197 : {{1'd0}, io_c[30:23]}; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_199 = _T_147 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  wire [7:0] _GEN_12 = {{6'd0}, _T_199}; // @[rawFloatFromFN.scala 60:22]
  wire [7:0] _T_200 = 8'h80 | _GEN_12; // @[rawFloatFromFN.scala 60:22]
  wire [8:0] _GEN_13 = {{1'd0}, _T_200}; // @[rawFloatFromFN.scala 59:15]
  wire [8:0] _T_202 = _T_198 + _GEN_13; // @[rawFloatFromFN.scala 59:15]
  wire  _T_203 = _T_147 & _T_148; // @[rawFloatFromFN.scala 62:34]
  wire  _T_205 = _T_202[8:7] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  wire  _T_207 = _T_205 & ~_T_148; // @[rawFloatFromFN.scala 66:33]
  wire [9:0] _T_210 = {1'b0,$signed(_T_202)}; // @[rawFloatFromFN.scala 70:48]
  wire  hi_lo_4 = ~_T_203; // @[rawFloatFromFN.scala 72:29]
  wire [22:0] lo_4 = _T_147 ? _T_196 : io_c[22:0]; // @[rawFloatFromFN.scala 72:42]
  wire [24:0] _T_211 = {1'h0,hi_lo_4,lo_4}; // @[Cat.scala 30:58]
  wire [2:0] _T_213 = _T_203 ? 3'h0 : _T_210[8:6]; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_14 = {{2'd0}, _T_207}; // @[recFNFromFN.scala 48:79]
  wire [2:0] hi_lo_5 = _T_213 | _GEN_14; // @[recFNFromFN.scala 48:79]
  wire [5:0] lo_hi_2 = _T_210[5:0]; // @[recFNFromFN.scala 50:23]
  wire [22:0] lo_lo_2 = _T_211[22:0]; // @[recFNFromFN.scala 51:22]
  wire [28:0] lo_5 = {lo_hi_2,lo_lo_2}; // @[Cat.scala 30:58]
  wire [3:0] hi_5 = {io_c[31],hi_lo_5}; // @[Cat.scala 30:58]
  wire [47:0] _T_216 = premul_a * premul_b; // @[FMULADD_1G_2.scala 113:19]
  wire  _T_219 = roundRawFNToRecFN_io_out[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_221 = roundRawFNToRecFN_io_out[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  wire  _T_223 = _T_221 & roundRawFNToRecFN_io_out[29]; // @[rawFloatFromRecFN.scala 55:33]
  wire  _T_226 = _T_221 & ~roundRawFNToRecFN_io_out[29]; // @[rawFloatFromRecFN.scala 56:33]
  wire [9:0] _T_228 = {1'b0,$signed(roundRawFNToRecFN_io_out[31:23])}; // @[rawFloatFromRecFN.scala 59:27]
  wire  hi_lo_6 = ~_T_219; // @[rawFloatFromRecFN.scala 60:39]
  wire [22:0] lo_6 = roundRawFNToRecFN_io_out[22:0]; // @[rawFloatFromRecFN.scala 60:51]
  wire [24:0] _T_229 = {1'h0,hi_lo_6,lo_6}; // @[Cat.scala 30:58]
  wire  _T_230 = $signed(_T_228) < 10'sh82; // @[fNFromRecFN.scala 50:39]
  wire [4:0] _T_233 = 5'h1 - _T_228[4:0]; // @[fNFromRecFN.scala 51:39]
  wire [23:0] _T_235 = _T_229[24:1] >> _T_233; // @[fNFromRecFN.scala 52:42]
  wire [7:0] _T_239 = _T_228[7:0] - 8'h81; // @[fNFromRecFN.scala 57:45]
  wire [7:0] _T_240 = _T_230 ? 8'h0 : _T_239; // @[fNFromRecFN.scala 55:16]
  wire  _T_241 = _T_223 | _T_226; // @[fNFromRecFN.scala 59:44]
  wire [7:0] _T_243 = _T_241 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] hi_lo_7 = _T_240 | _T_243; // @[fNFromRecFN.scala 59:15]
  wire [22:0] _T_245 = _T_226 ? 23'h0 : _T_229[22:0]; // @[fNFromRecFN.scala 63:20]
  wire [22:0] lo_7 = _T_230 ? _T_235[22:0] : _T_245; // @[fNFromRecFN.scala 61:16]
  wire [8:0] hi_7 = {roundRawFNToRecFN_io_out[32],hi_lo_7}; // @[Cat.scala 30:58]
  MulAddRecFNToRaw_preMul mulAddRecFNToRaw_preMul ( // @[FMULADD_1G_2.scala 36:15]
    .io_a(mulAddRecFNToRaw_preMul_io_a),
    .io_b(mulAddRecFNToRaw_preMul_io_b),
    .io_c(mulAddRecFNToRaw_preMul_io_c),
    .io_mulAddA(mulAddRecFNToRaw_preMul_io_mulAddA),
    .io_mulAddB(mulAddRecFNToRaw_preMul_io_mulAddB),
    .io_mulAddC(mulAddRecFNToRaw_preMul_io_mulAddC),
    .io_toPostMul_isSigNaNAny(mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny),
    .io_toPostMul_isNaNAOrB(mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB),
    .io_toPostMul_isInfA(mulAddRecFNToRaw_preMul_io_toPostMul_isInfA),
    .io_toPostMul_isZeroA(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA),
    .io_toPostMul_isInfB(mulAddRecFNToRaw_preMul_io_toPostMul_isInfB),
    .io_toPostMul_isZeroB(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB),
    .io_toPostMul_signProd(mulAddRecFNToRaw_preMul_io_toPostMul_signProd),
    .io_toPostMul_isNaNC(mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC),
    .io_toPostMul_isInfC(mulAddRecFNToRaw_preMul_io_toPostMul_isInfC),
    .io_toPostMul_isZeroC(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC),
    .io_toPostMul_sExpSum(mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum),
    .io_toPostMul_doSubMags(mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags),
    .io_toPostMul_CIsDominant(mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant),
    .io_toPostMul_CDom_CAlignDist(mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist),
    .io_toPostMul_highAlignedSigC(mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC),
    .io_toPostMul_bit0AlignedSigC(mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC)
  );
  MulAddRecFNToRaw_postMul mulAddRecFNToRaw_postMul ( // @[FMULADD_1G_2.scala 116:15]
    .io_fromPreMul_isSigNaNAny(mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny),
    .io_fromPreMul_isNaNAOrB(mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB),
    .io_fromPreMul_isInfA(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA),
    .io_fromPreMul_isZeroA(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA),
    .io_fromPreMul_isInfB(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB),
    .io_fromPreMul_isZeroB(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB),
    .io_fromPreMul_signProd(mulAddRecFNToRaw_postMul_io_fromPreMul_signProd),
    .io_fromPreMul_isNaNC(mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC),
    .io_fromPreMul_isInfC(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC),
    .io_fromPreMul_isZeroC(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC),
    .io_fromPreMul_sExpSum(mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum),
    .io_fromPreMul_doSubMags(mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags),
    .io_fromPreMul_CIsDominant(mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant),
    .io_fromPreMul_CDom_CAlignDist(mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist),
    .io_fromPreMul_highAlignedSigC(mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC),
    .io_fromPreMul_bit0AlignedSigC(mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC),
    .io_mulAddResult(mulAddRecFNToRaw_postMul_io_mulAddResult),
    .io_invalidExc(mulAddRecFNToRaw_postMul_io_invalidExc),
    .io_rawOut_isNaN(mulAddRecFNToRaw_postMul_io_rawOut_isNaN),
    .io_rawOut_isInf(mulAddRecFNToRaw_postMul_io_rawOut_isInf),
    .io_rawOut_isZero(mulAddRecFNToRaw_postMul_io_rawOut_isZero),
    .io_rawOut_sign(mulAddRecFNToRaw_postMul_io_rawOut_sign),
    .io_rawOut_sExp(mulAddRecFNToRaw_postMul_io_rawOut_sExp),
    .io_rawOut_sig(mulAddRecFNToRaw_postMul_io_rawOut_sig)
  );
  RoundRawFNToRecFN roundRawFNToRecFN ( // @[FMULADD_1G_2.scala 137:15]
    .io_invalidExc(roundRawFNToRecFN_io_invalidExc),
    .io_in_isNaN(roundRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundRawFNToRecFN_io_in_sig),
    .io_out(roundRawFNToRecFN_io_out)
  );
  assign io_out = {hi_7,lo_7}; // @[Cat.scala 30:58]
  assign mulAddRecFNToRaw_preMul_io_a = {hi_1,lo_1}; // @[Cat.scala 30:58]
  assign mulAddRecFNToRaw_preMul_io_b = {hi_3,lo_3}; // @[Cat.scala 30:58]
  assign mulAddRecFNToRaw_preMul_io_c = {hi_5,lo_5}; // @[Cat.scala 30:58]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny = isSigNaNAny; // @[FMULADD_1G_2.scala 119:84]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB = isNaNAOrB; // @[FMULADD_1G_2.scala 120:86]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA = isInfA; // @[FMULADD_1G_2.scala 121:94]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA = isZeroA; // @[FMULADD_1G_2.scala 122:91]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB = isInfB; // @[FMULADD_1G_2.scala 123:94]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB = isZeroB; // @[FMULADD_1G_2.scala 124:91]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_signProd = signProd; // @[FMULADD_1G_2.scala 125:89]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC = isNaNC; // @[FMULADD_1G_2.scala 126:90]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC = isInfC; // @[FMULADD_1G_2.scala 127:94]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC = isZeroC; // @[FMULADD_1G_2.scala 128:91]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum = sExpSum; // @[FMULADD_1G_2.scala 129:88]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags = doSubMags; // @[FMULADD_1G_2.scala 130:85]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant = CIsDominant; // @[FMULADD_1G_2.scala 131:84]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist = CDom_CAlignDist; // @[FMULADD_1G_2.scala 132:78]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC = highAlignedSigC; // @[FMULADD_1G_2.scala 133:80]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC = bit0AlignedSigC; // @[FMULADD_1G_2.scala 134:82]
  assign mulAddRecFNToRaw_postMul_io_mulAddResult = _T_216 + premul_c; // @[FMULADD_1G_2.scala 113:31]
  assign roundRawFNToRecFN_io_invalidExc = mulAddRecFNToRaw_postMul_io_invalidExc; // @[FMULADD_1G_2.scala 138:39]
  assign roundRawFNToRecFN_io_in_isNaN = mulAddRecFNToRaw_postMul_io_rawOut_isNaN; // @[FMULADD_1G_2.scala 140:39]
  assign roundRawFNToRecFN_io_in_isInf = mulAddRecFNToRaw_postMul_io_rawOut_isInf; // @[FMULADD_1G_2.scala 140:39]
  assign roundRawFNToRecFN_io_in_isZero = mulAddRecFNToRaw_postMul_io_rawOut_isZero; // @[FMULADD_1G_2.scala 140:39]
  assign roundRawFNToRecFN_io_in_sign = mulAddRecFNToRaw_postMul_io_rawOut_sign; // @[FMULADD_1G_2.scala 140:39]
  assign roundRawFNToRecFN_io_in_sExp = mulAddRecFNToRaw_postMul_io_rawOut_sExp; // @[FMULADD_1G_2.scala 140:39]
  assign roundRawFNToRecFN_io_in_sig = mulAddRecFNToRaw_postMul_io_rawOut_sig; // @[FMULADD_1G_2.scala 140:39]
  always @(posedge clock) begin
    if (reset) begin // @[FMULADD_1G_2.scala 15:37]
      premul_a <= 24'h0; // @[FMULADD_1G_2.scala 15:37]
    end else begin
      premul_a <= mulAddRecFNToRaw_preMul_io_mulAddA; // @[FMULADD_1G_2.scala 103:63]
    end
    if (reset) begin // @[FMULADD_1G_2.scala 16:37]
      premul_b <= 24'h0; // @[FMULADD_1G_2.scala 16:37]
    end else begin
      premul_b <= mulAddRecFNToRaw_preMul_io_mulAddB; // @[FMULADD_1G_2.scala 104:63]
    end
    if (reset) begin // @[FMULADD_1G_2.scala 17:37]
      premul_c <= 48'h0; // @[FMULADD_1G_2.scala 17:37]
    end else begin
      premul_c <= mulAddRecFNToRaw_preMul_io_mulAddC; // @[FMULADD_1G_2.scala 105:63]
    end
    if (reset) begin // @[FMULADD_1G_2.scala 18:33]
      isSigNaNAny <= 1'h0; // @[FMULADD_1G_2.scala 18:33]
    end else begin
      isSigNaNAny <= mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny; // @[FMULADD_1G_2.scala 43:61]
    end
    if (reset) begin // @[FMULADD_1G_2.scala 19:34]
      isNaNAOrB <= 1'h0; // @[FMULADD_1G_2.scala 19:34]
    end else begin
      isNaNAOrB <= mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB; // @[FMULADD_1G_2.scala 44:62]
    end
    if (reset) begin // @[FMULADD_1G_2.scala 20:43]
      isInfA <= 1'h0; // @[FMULADD_1G_2.scala 20:43]
    end else begin
      isInfA <= mulAddRecFNToRaw_preMul_io_toPostMul_isInfA; // @[FMULADD_1G_2.scala 45:70]
    end
    if (reset) begin // @[FMULADD_1G_2.scala 21:40]
      isZeroA <= 1'h0; // @[FMULADD_1G_2.scala 21:40]
    end else begin
      isZeroA <= mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA; // @[FMULADD_1G_2.scala 46:67]
    end
    if (reset) begin // @[FMULADD_1G_2.scala 22:43]
      isInfB <= 1'h0; // @[FMULADD_1G_2.scala 22:43]
    end else begin
      isInfB <= mulAddRecFNToRaw_preMul_io_toPostMul_isInfB; // @[FMULADD_1G_2.scala 47:70]
    end
    if (reset) begin // @[FMULADD_1G_2.scala 23:40]
      isZeroB <= 1'h0; // @[FMULADD_1G_2.scala 23:40]
    end else begin
      isZeroB <= mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB; // @[FMULADD_1G_2.scala 48:67]
    end
    if (reset) begin // @[FMULADD_1G_2.scala 24:38]
      signProd <= 1'h0; // @[FMULADD_1G_2.scala 24:38]
    end else begin
      signProd <= mulAddRecFNToRaw_preMul_io_toPostMul_signProd; // @[FMULADD_1G_2.scala 49:65]
    end
    if (reset) begin // @[FMULADD_1G_2.scala 25:39]
      isNaNC <= 1'h0; // @[FMULADD_1G_2.scala 25:39]
    end else begin
      isNaNC <= mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC; // @[FMULADD_1G_2.scala 50:66]
    end
    if (reset) begin // @[FMULADD_1G_2.scala 26:42]
      isInfC <= 1'h0; // @[FMULADD_1G_2.scala 26:42]
    end else begin
      isInfC <= mulAddRecFNToRaw_preMul_io_toPostMul_isInfC; // @[FMULADD_1G_2.scala 51:69]
    end
    if (reset) begin // @[FMULADD_1G_2.scala 27:39]
      isZeroC <= 1'h0; // @[FMULADD_1G_2.scala 27:39]
    end else begin
      isZeroC <= mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC; // @[FMULADD_1G_2.scala 52:66]
    end
    if (reset) begin // @[FMULADD_1G_2.scala 28:36]
      sExpSum <= 10'sh0; // @[FMULADD_1G_2.scala 28:36]
    end else begin
      sExpSum <= mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum; // @[FMULADD_1G_2.scala 53:63]
    end
    if (reset) begin // @[FMULADD_1G_2.scala 29:33]
      doSubMags <= 1'h0; // @[FMULADD_1G_2.scala 29:33]
    end else begin
      doSubMags <= mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags; // @[FMULADD_1G_2.scala 54:60]
    end
    if (reset) begin // @[FMULADD_1G_2.scala 30:33]
      CIsDominant <= 1'h0; // @[FMULADD_1G_2.scala 30:33]
    end else begin
      CIsDominant <= mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant; // @[FMULADD_1G_2.scala 55:59]
    end
    if (reset) begin // @[FMULADD_1G_2.scala 31:34]
      CDom_CAlignDist <= 5'h0; // @[FMULADD_1G_2.scala 31:34]
    end else begin
      CDom_CAlignDist <= mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist; // @[FMULADD_1G_2.scala 56:54]
    end
    if (reset) begin // @[FMULADD_1G_2.scala 32:37]
      highAlignedSigC <= 26'h0; // @[FMULADD_1G_2.scala 32:37]
    end else begin
      highAlignedSigC <= mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC; // @[FMULADD_1G_2.scala 57:56]
    end
    if (reset) begin // @[FMULADD_1G_2.scala 33:38]
      bit0AlignedSigC <= 1'h0; // @[FMULADD_1G_2.scala 33:38]
    end else begin
      bit0AlignedSigC <= mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC; // @[FMULADD_1G_2.scala 58:57]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  premul_a = _RAND_0[23:0];
  _RAND_1 = {1{`RANDOM}};
  premul_b = _RAND_1[23:0];
  _RAND_2 = {2{`RANDOM}};
  premul_c = _RAND_2[47:0];
  _RAND_3 = {1{`RANDOM}};
  isSigNaNAny = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  isNaNAOrB = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  isInfA = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  isZeroA = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  isInfB = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  isZeroB = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  signProd = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  isNaNC = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  isInfC = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  isZeroC = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  sExpSum = _RAND_13[9:0];
  _RAND_14 = {1{`RANDOM}};
  doSubMags = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  CIsDominant = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  CDom_CAlignDist = _RAND_16[4:0];
  _RAND_17 = {1{`RANDOM}};
  highAlignedSigC = _RAND_17[25:0];
  _RAND_18 = {1{`RANDOM}};
  bit0AlignedSigC = _RAND_18[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CompareRecFN(
  input  [32:0] io_a,
  input  [32:0] io_b,
  output        io_lt,
  output        io_eq
);
  wire  rawA_isZero = io_a[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_4 = io_a[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawA_isNaN = _T_4 & io_a[29]; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawA_isInf = _T_4 & ~io_a[29]; // @[rawFloatFromRecFN.scala 56:33]
  wire  rawA_sign = io_a[32]; // @[rawFloatFromRecFN.scala 58:25]
  wire [9:0] rawA_sExp = {1'b0,$signed(io_a[31:23])}; // @[rawFloatFromRecFN.scala 59:27]
  wire  hi_lo = ~rawA_isZero; // @[rawFloatFromRecFN.scala 60:39]
  wire [22:0] lo = io_a[22:0]; // @[rawFloatFromRecFN.scala 60:51]
  wire [24:0] rawA_sig = {1'h0,hi_lo,lo}; // @[Cat.scala 30:58]
  wire  rawB_isZero = io_b[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_17 = io_b[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawB_isNaN = _T_17 & io_b[29]; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawB_isInf = _T_17 & ~io_b[29]; // @[rawFloatFromRecFN.scala 56:33]
  wire  rawB_sign = io_b[32]; // @[rawFloatFromRecFN.scala 58:25]
  wire [9:0] rawB_sExp = {1'b0,$signed(io_b[31:23])}; // @[rawFloatFromRecFN.scala 59:27]
  wire  hi_lo_1 = ~rawB_isZero; // @[rawFloatFromRecFN.scala 60:39]
  wire [22:0] lo_1 = io_b[22:0]; // @[rawFloatFromRecFN.scala 60:51]
  wire [24:0] rawB_sig = {1'h0,hi_lo_1,lo_1}; // @[Cat.scala 30:58]
  wire  ordered = ~rawA_isNaN & ~rawB_isNaN; // @[CompareRecFN.scala 57:32]
  wire  bothInfs = rawA_isInf & rawB_isInf; // @[CompareRecFN.scala 58:33]
  wire  bothZeros = rawA_isZero & rawB_isZero; // @[CompareRecFN.scala 59:33]
  wire  eqExps = $signed(rawA_sExp) == $signed(rawB_sExp); // @[CompareRecFN.scala 60:29]
  wire  common_ltMags = $signed(rawA_sExp) < $signed(rawB_sExp) | eqExps & rawA_sig < rawB_sig; // @[CompareRecFN.scala 62:33]
  wire  common_eqMags = eqExps & rawA_sig == rawB_sig; // @[CompareRecFN.scala 63:32]
  wire  _T_33 = ~rawB_sign; // @[CompareRecFN.scala 67:28]
  wire  _T_41 = _T_33 & common_ltMags; // @[CompareRecFN.scala 70:41]
  wire  _T_42 = rawA_sign & ~common_ltMags & ~common_eqMags | _T_41; // @[CompareRecFN.scala 69:74]
  wire  _T_43 = ~bothInfs & _T_42; // @[CompareRecFN.scala 68:30]
  wire  _T_44 = rawA_sign & ~rawB_sign | _T_43; // @[CompareRecFN.scala 67:41]
  wire  ordered_lt = ~bothZeros & _T_44; // @[CompareRecFN.scala 66:21]
  wire  ordered_eq = bothZeros | rawA_sign == rawB_sign & (bothInfs | common_eqMags); // @[CompareRecFN.scala 72:19]
  assign io_lt = ordered & ordered_lt; // @[CompareRecFN.scala 78:22]
  assign io_eq = ordered & ordered_eq; // @[CompareRecFN.scala 79:22]
endmodule
module ValExec_CompareRecF32_le(
  input  [31:0] io_a,
  input  [31:0] io_b,
  output        io_actual_out
);
  wire [32:0] compareRecFN_io_a; // @[ValExec_CompareRecFN.scala 94:30]
  wire [32:0] compareRecFN_io_b; // @[ValExec_CompareRecFN.scala 94:30]
  wire  compareRecFN_io_lt; // @[ValExec_CompareRecFN.scala 94:30]
  wire  compareRecFN_io_eq; // @[ValExec_CompareRecFN.scala 94:30]
  wire  _T_3 = io_a[30:23] == 8'h0; // @[rawFloatFromFN.scala 50:34]
  wire  _T_4 = io_a[22:0] == 23'h0; // @[rawFloatFromFN.scala 51:38]
  wire [4:0] _T_28 = io_a[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:69]
  wire [4:0] _T_29 = io_a[2] ? 5'h14 : _T_28; // @[Mux.scala 47:69]
  wire [4:0] _T_30 = io_a[3] ? 5'h13 : _T_29; // @[Mux.scala 47:69]
  wire [4:0] _T_31 = io_a[4] ? 5'h12 : _T_30; // @[Mux.scala 47:69]
  wire [4:0] _T_32 = io_a[5] ? 5'h11 : _T_31; // @[Mux.scala 47:69]
  wire [4:0] _T_33 = io_a[6] ? 5'h10 : _T_32; // @[Mux.scala 47:69]
  wire [4:0] _T_34 = io_a[7] ? 5'hf : _T_33; // @[Mux.scala 47:69]
  wire [4:0] _T_35 = io_a[8] ? 5'he : _T_34; // @[Mux.scala 47:69]
  wire [4:0] _T_36 = io_a[9] ? 5'hd : _T_35; // @[Mux.scala 47:69]
  wire [4:0] _T_37 = io_a[10] ? 5'hc : _T_36; // @[Mux.scala 47:69]
  wire [4:0] _T_38 = io_a[11] ? 5'hb : _T_37; // @[Mux.scala 47:69]
  wire [4:0] _T_39 = io_a[12] ? 5'ha : _T_38; // @[Mux.scala 47:69]
  wire [4:0] _T_40 = io_a[13] ? 5'h9 : _T_39; // @[Mux.scala 47:69]
  wire [4:0] _T_41 = io_a[14] ? 5'h8 : _T_40; // @[Mux.scala 47:69]
  wire [4:0] _T_42 = io_a[15] ? 5'h7 : _T_41; // @[Mux.scala 47:69]
  wire [4:0] _T_43 = io_a[16] ? 5'h6 : _T_42; // @[Mux.scala 47:69]
  wire [4:0] _T_44 = io_a[17] ? 5'h5 : _T_43; // @[Mux.scala 47:69]
  wire [4:0] _T_45 = io_a[18] ? 5'h4 : _T_44; // @[Mux.scala 47:69]
  wire [4:0] _T_46 = io_a[19] ? 5'h3 : _T_45; // @[Mux.scala 47:69]
  wire [4:0] _T_47 = io_a[20] ? 5'h2 : _T_46; // @[Mux.scala 47:69]
  wire [4:0] _T_48 = io_a[21] ? 5'h1 : _T_47; // @[Mux.scala 47:69]
  wire [4:0] _T_49 = io_a[22] ? 5'h0 : _T_48; // @[Mux.scala 47:69]
  wire [53:0] _GEN_0 = {{31'd0}, io_a[22:0]}; // @[rawFloatFromFN.scala 54:36]
  wire [53:0] _T_50 = _GEN_0 << _T_49; // @[rawFloatFromFN.scala 54:36]
  wire [22:0] _T_52 = {_T_50[21:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  wire [8:0] _GEN_1 = {{4'd0}, _T_49}; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_53 = _GEN_1 ^ 9'h1ff; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_54 = _T_3 ? _T_53 : {{1'd0}, io_a[30:23]}; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_55 = _T_3 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  wire [7:0] _GEN_2 = {{6'd0}, _T_55}; // @[rawFloatFromFN.scala 60:22]
  wire [7:0] _T_56 = 8'h80 | _GEN_2; // @[rawFloatFromFN.scala 60:22]
  wire [8:0] _GEN_3 = {{1'd0}, _T_56}; // @[rawFloatFromFN.scala 59:15]
  wire [8:0] _T_58 = _T_54 + _GEN_3; // @[rawFloatFromFN.scala 59:15]
  wire  _T_59 = _T_3 & _T_4; // @[rawFloatFromFN.scala 62:34]
  wire  _T_61 = _T_58[8:7] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  wire  _T_63 = _T_61 & ~_T_4; // @[rawFloatFromFN.scala 66:33]
  wire [9:0] _T_66 = {1'b0,$signed(_T_58)}; // @[rawFloatFromFN.scala 70:48]
  wire  hi_lo = ~_T_59; // @[rawFloatFromFN.scala 72:29]
  wire [22:0] lo = _T_3 ? _T_52 : io_a[22:0]; // @[rawFloatFromFN.scala 72:42]
  wire [24:0] _T_67 = {1'h0,hi_lo,lo}; // @[Cat.scala 30:58]
  wire [2:0] _T_69 = _T_59 ? 3'h0 : _T_66[8:6]; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_4 = {{2'd0}, _T_63}; // @[recFNFromFN.scala 48:79]
  wire [2:0] hi_lo_1 = _T_69 | _GEN_4; // @[recFNFromFN.scala 48:79]
  wire [5:0] lo_hi = _T_66[5:0]; // @[recFNFromFN.scala 50:23]
  wire [22:0] lo_lo = _T_67[22:0]; // @[recFNFromFN.scala 51:22]
  wire [28:0] lo_1 = {lo_hi,lo_lo}; // @[Cat.scala 30:58]
  wire [3:0] hi_1 = {io_a[31],hi_lo_1}; // @[Cat.scala 30:58]
  wire  _T_75 = io_b[30:23] == 8'h0; // @[rawFloatFromFN.scala 50:34]
  wire  _T_76 = io_b[22:0] == 23'h0; // @[rawFloatFromFN.scala 51:38]
  wire [4:0] _T_100 = io_b[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:69]
  wire [4:0] _T_101 = io_b[2] ? 5'h14 : _T_100; // @[Mux.scala 47:69]
  wire [4:0] _T_102 = io_b[3] ? 5'h13 : _T_101; // @[Mux.scala 47:69]
  wire [4:0] _T_103 = io_b[4] ? 5'h12 : _T_102; // @[Mux.scala 47:69]
  wire [4:0] _T_104 = io_b[5] ? 5'h11 : _T_103; // @[Mux.scala 47:69]
  wire [4:0] _T_105 = io_b[6] ? 5'h10 : _T_104; // @[Mux.scala 47:69]
  wire [4:0] _T_106 = io_b[7] ? 5'hf : _T_105; // @[Mux.scala 47:69]
  wire [4:0] _T_107 = io_b[8] ? 5'he : _T_106; // @[Mux.scala 47:69]
  wire [4:0] _T_108 = io_b[9] ? 5'hd : _T_107; // @[Mux.scala 47:69]
  wire [4:0] _T_109 = io_b[10] ? 5'hc : _T_108; // @[Mux.scala 47:69]
  wire [4:0] _T_110 = io_b[11] ? 5'hb : _T_109; // @[Mux.scala 47:69]
  wire [4:0] _T_111 = io_b[12] ? 5'ha : _T_110; // @[Mux.scala 47:69]
  wire [4:0] _T_112 = io_b[13] ? 5'h9 : _T_111; // @[Mux.scala 47:69]
  wire [4:0] _T_113 = io_b[14] ? 5'h8 : _T_112; // @[Mux.scala 47:69]
  wire [4:0] _T_114 = io_b[15] ? 5'h7 : _T_113; // @[Mux.scala 47:69]
  wire [4:0] _T_115 = io_b[16] ? 5'h6 : _T_114; // @[Mux.scala 47:69]
  wire [4:0] _T_116 = io_b[17] ? 5'h5 : _T_115; // @[Mux.scala 47:69]
  wire [4:0] _T_117 = io_b[18] ? 5'h4 : _T_116; // @[Mux.scala 47:69]
  wire [4:0] _T_118 = io_b[19] ? 5'h3 : _T_117; // @[Mux.scala 47:69]
  wire [4:0] _T_119 = io_b[20] ? 5'h2 : _T_118; // @[Mux.scala 47:69]
  wire [4:0] _T_120 = io_b[21] ? 5'h1 : _T_119; // @[Mux.scala 47:69]
  wire [4:0] _T_121 = io_b[22] ? 5'h0 : _T_120; // @[Mux.scala 47:69]
  wire [53:0] _GEN_5 = {{31'd0}, io_b[22:0]}; // @[rawFloatFromFN.scala 54:36]
  wire [53:0] _T_122 = _GEN_5 << _T_121; // @[rawFloatFromFN.scala 54:36]
  wire [22:0] _T_124 = {_T_122[21:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  wire [8:0] _GEN_6 = {{4'd0}, _T_121}; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_125 = _GEN_6 ^ 9'h1ff; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_126 = _T_75 ? _T_125 : {{1'd0}, io_b[30:23]}; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_127 = _T_75 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  wire [7:0] _GEN_7 = {{6'd0}, _T_127}; // @[rawFloatFromFN.scala 60:22]
  wire [7:0] _T_128 = 8'h80 | _GEN_7; // @[rawFloatFromFN.scala 60:22]
  wire [8:0] _GEN_8 = {{1'd0}, _T_128}; // @[rawFloatFromFN.scala 59:15]
  wire [8:0] _T_130 = _T_126 + _GEN_8; // @[rawFloatFromFN.scala 59:15]
  wire  _T_131 = _T_75 & _T_76; // @[rawFloatFromFN.scala 62:34]
  wire  _T_133 = _T_130[8:7] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  wire  _T_135 = _T_133 & ~_T_76; // @[rawFloatFromFN.scala 66:33]
  wire [9:0] _T_138 = {1'b0,$signed(_T_130)}; // @[rawFloatFromFN.scala 70:48]
  wire  hi_lo_2 = ~_T_131; // @[rawFloatFromFN.scala 72:29]
  wire [22:0] lo_2 = _T_75 ? _T_124 : io_b[22:0]; // @[rawFloatFromFN.scala 72:42]
  wire [24:0] _T_139 = {1'h0,hi_lo_2,lo_2}; // @[Cat.scala 30:58]
  wire [2:0] _T_141 = _T_131 ? 3'h0 : _T_138[8:6]; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_9 = {{2'd0}, _T_135}; // @[recFNFromFN.scala 48:79]
  wire [2:0] hi_lo_3 = _T_141 | _GEN_9; // @[recFNFromFN.scala 48:79]
  wire [5:0] lo_hi_1 = _T_138[5:0]; // @[recFNFromFN.scala 50:23]
  wire [22:0] lo_lo_1 = _T_139[22:0]; // @[recFNFromFN.scala 51:22]
  wire [28:0] lo_3 = {lo_hi_1,lo_lo_1}; // @[Cat.scala 30:58]
  wire [3:0] hi_3 = {io_b[31],hi_lo_3}; // @[Cat.scala 30:58]
  CompareRecFN compareRecFN ( // @[ValExec_CompareRecFN.scala 94:30]
    .io_a(compareRecFN_io_a),
    .io_b(compareRecFN_io_b),
    .io_lt(compareRecFN_io_lt),
    .io_eq(compareRecFN_io_eq)
  );
  assign io_actual_out = compareRecFN_io_lt | compareRecFN_io_eq; // @[ValExec_CompareRecFN.scala 99:41]
  assign compareRecFN_io_a = {hi_1,lo_1}; // @[Cat.scala 30:58]
  assign compareRecFN_io_b = {hi_3,lo_3}; // @[Cat.scala 30:58]
endmodule
module ValExec_CompareRecF32_lt(
  input  [31:0] io_a,
  input  [31:0] io_b,
  output        io_actual_out
);
  wire [32:0] compareRecFN_io_a; // @[ValExec_CompareRecFN.scala 59:30]
  wire [32:0] compareRecFN_io_b; // @[ValExec_CompareRecFN.scala 59:30]
  wire  compareRecFN_io_lt; // @[ValExec_CompareRecFN.scala 59:30]
  wire  compareRecFN_io_eq; // @[ValExec_CompareRecFN.scala 59:30]
  wire  _T_3 = io_a[30:23] == 8'h0; // @[rawFloatFromFN.scala 50:34]
  wire  _T_4 = io_a[22:0] == 23'h0; // @[rawFloatFromFN.scala 51:38]
  wire [4:0] _T_28 = io_a[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:69]
  wire [4:0] _T_29 = io_a[2] ? 5'h14 : _T_28; // @[Mux.scala 47:69]
  wire [4:0] _T_30 = io_a[3] ? 5'h13 : _T_29; // @[Mux.scala 47:69]
  wire [4:0] _T_31 = io_a[4] ? 5'h12 : _T_30; // @[Mux.scala 47:69]
  wire [4:0] _T_32 = io_a[5] ? 5'h11 : _T_31; // @[Mux.scala 47:69]
  wire [4:0] _T_33 = io_a[6] ? 5'h10 : _T_32; // @[Mux.scala 47:69]
  wire [4:0] _T_34 = io_a[7] ? 5'hf : _T_33; // @[Mux.scala 47:69]
  wire [4:0] _T_35 = io_a[8] ? 5'he : _T_34; // @[Mux.scala 47:69]
  wire [4:0] _T_36 = io_a[9] ? 5'hd : _T_35; // @[Mux.scala 47:69]
  wire [4:0] _T_37 = io_a[10] ? 5'hc : _T_36; // @[Mux.scala 47:69]
  wire [4:0] _T_38 = io_a[11] ? 5'hb : _T_37; // @[Mux.scala 47:69]
  wire [4:0] _T_39 = io_a[12] ? 5'ha : _T_38; // @[Mux.scala 47:69]
  wire [4:0] _T_40 = io_a[13] ? 5'h9 : _T_39; // @[Mux.scala 47:69]
  wire [4:0] _T_41 = io_a[14] ? 5'h8 : _T_40; // @[Mux.scala 47:69]
  wire [4:0] _T_42 = io_a[15] ? 5'h7 : _T_41; // @[Mux.scala 47:69]
  wire [4:0] _T_43 = io_a[16] ? 5'h6 : _T_42; // @[Mux.scala 47:69]
  wire [4:0] _T_44 = io_a[17] ? 5'h5 : _T_43; // @[Mux.scala 47:69]
  wire [4:0] _T_45 = io_a[18] ? 5'h4 : _T_44; // @[Mux.scala 47:69]
  wire [4:0] _T_46 = io_a[19] ? 5'h3 : _T_45; // @[Mux.scala 47:69]
  wire [4:0] _T_47 = io_a[20] ? 5'h2 : _T_46; // @[Mux.scala 47:69]
  wire [4:0] _T_48 = io_a[21] ? 5'h1 : _T_47; // @[Mux.scala 47:69]
  wire [4:0] _T_49 = io_a[22] ? 5'h0 : _T_48; // @[Mux.scala 47:69]
  wire [53:0] _GEN_0 = {{31'd0}, io_a[22:0]}; // @[rawFloatFromFN.scala 54:36]
  wire [53:0] _T_50 = _GEN_0 << _T_49; // @[rawFloatFromFN.scala 54:36]
  wire [22:0] _T_52 = {_T_50[21:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  wire [8:0] _GEN_1 = {{4'd0}, _T_49}; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_53 = _GEN_1 ^ 9'h1ff; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_54 = _T_3 ? _T_53 : {{1'd0}, io_a[30:23]}; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_55 = _T_3 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  wire [7:0] _GEN_2 = {{6'd0}, _T_55}; // @[rawFloatFromFN.scala 60:22]
  wire [7:0] _T_56 = 8'h80 | _GEN_2; // @[rawFloatFromFN.scala 60:22]
  wire [8:0] _GEN_3 = {{1'd0}, _T_56}; // @[rawFloatFromFN.scala 59:15]
  wire [8:0] _T_58 = _T_54 + _GEN_3; // @[rawFloatFromFN.scala 59:15]
  wire  _T_59 = _T_3 & _T_4; // @[rawFloatFromFN.scala 62:34]
  wire  _T_61 = _T_58[8:7] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  wire  _T_63 = _T_61 & ~_T_4; // @[rawFloatFromFN.scala 66:33]
  wire [9:0] _T_66 = {1'b0,$signed(_T_58)}; // @[rawFloatFromFN.scala 70:48]
  wire  hi_lo = ~_T_59; // @[rawFloatFromFN.scala 72:29]
  wire [22:0] lo = _T_3 ? _T_52 : io_a[22:0]; // @[rawFloatFromFN.scala 72:42]
  wire [24:0] _T_67 = {1'h0,hi_lo,lo}; // @[Cat.scala 30:58]
  wire [2:0] _T_69 = _T_59 ? 3'h0 : _T_66[8:6]; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_4 = {{2'd0}, _T_63}; // @[recFNFromFN.scala 48:79]
  wire [2:0] hi_lo_1 = _T_69 | _GEN_4; // @[recFNFromFN.scala 48:79]
  wire [5:0] lo_hi = _T_66[5:0]; // @[recFNFromFN.scala 50:23]
  wire [22:0] lo_lo = _T_67[22:0]; // @[recFNFromFN.scala 51:22]
  wire [28:0] lo_1 = {lo_hi,lo_lo}; // @[Cat.scala 30:58]
  wire [3:0] hi_1 = {io_a[31],hi_lo_1}; // @[Cat.scala 30:58]
  wire  _T_75 = io_b[30:23] == 8'h0; // @[rawFloatFromFN.scala 50:34]
  wire  _T_76 = io_b[22:0] == 23'h0; // @[rawFloatFromFN.scala 51:38]
  wire [4:0] _T_100 = io_b[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:69]
  wire [4:0] _T_101 = io_b[2] ? 5'h14 : _T_100; // @[Mux.scala 47:69]
  wire [4:0] _T_102 = io_b[3] ? 5'h13 : _T_101; // @[Mux.scala 47:69]
  wire [4:0] _T_103 = io_b[4] ? 5'h12 : _T_102; // @[Mux.scala 47:69]
  wire [4:0] _T_104 = io_b[5] ? 5'h11 : _T_103; // @[Mux.scala 47:69]
  wire [4:0] _T_105 = io_b[6] ? 5'h10 : _T_104; // @[Mux.scala 47:69]
  wire [4:0] _T_106 = io_b[7] ? 5'hf : _T_105; // @[Mux.scala 47:69]
  wire [4:0] _T_107 = io_b[8] ? 5'he : _T_106; // @[Mux.scala 47:69]
  wire [4:0] _T_108 = io_b[9] ? 5'hd : _T_107; // @[Mux.scala 47:69]
  wire [4:0] _T_109 = io_b[10] ? 5'hc : _T_108; // @[Mux.scala 47:69]
  wire [4:0] _T_110 = io_b[11] ? 5'hb : _T_109; // @[Mux.scala 47:69]
  wire [4:0] _T_111 = io_b[12] ? 5'ha : _T_110; // @[Mux.scala 47:69]
  wire [4:0] _T_112 = io_b[13] ? 5'h9 : _T_111; // @[Mux.scala 47:69]
  wire [4:0] _T_113 = io_b[14] ? 5'h8 : _T_112; // @[Mux.scala 47:69]
  wire [4:0] _T_114 = io_b[15] ? 5'h7 : _T_113; // @[Mux.scala 47:69]
  wire [4:0] _T_115 = io_b[16] ? 5'h6 : _T_114; // @[Mux.scala 47:69]
  wire [4:0] _T_116 = io_b[17] ? 5'h5 : _T_115; // @[Mux.scala 47:69]
  wire [4:0] _T_117 = io_b[18] ? 5'h4 : _T_116; // @[Mux.scala 47:69]
  wire [4:0] _T_118 = io_b[19] ? 5'h3 : _T_117; // @[Mux.scala 47:69]
  wire [4:0] _T_119 = io_b[20] ? 5'h2 : _T_118; // @[Mux.scala 47:69]
  wire [4:0] _T_120 = io_b[21] ? 5'h1 : _T_119; // @[Mux.scala 47:69]
  wire [4:0] _T_121 = io_b[22] ? 5'h0 : _T_120; // @[Mux.scala 47:69]
  wire [53:0] _GEN_5 = {{31'd0}, io_b[22:0]}; // @[rawFloatFromFN.scala 54:36]
  wire [53:0] _T_122 = _GEN_5 << _T_121; // @[rawFloatFromFN.scala 54:36]
  wire [22:0] _T_124 = {_T_122[21:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  wire [8:0] _GEN_6 = {{4'd0}, _T_121}; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_125 = _GEN_6 ^ 9'h1ff; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_126 = _T_75 ? _T_125 : {{1'd0}, io_b[30:23]}; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_127 = _T_75 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  wire [7:0] _GEN_7 = {{6'd0}, _T_127}; // @[rawFloatFromFN.scala 60:22]
  wire [7:0] _T_128 = 8'h80 | _GEN_7; // @[rawFloatFromFN.scala 60:22]
  wire [8:0] _GEN_8 = {{1'd0}, _T_128}; // @[rawFloatFromFN.scala 59:15]
  wire [8:0] _T_130 = _T_126 + _GEN_8; // @[rawFloatFromFN.scala 59:15]
  wire  _T_131 = _T_75 & _T_76; // @[rawFloatFromFN.scala 62:34]
  wire  _T_133 = _T_130[8:7] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  wire  _T_135 = _T_133 & ~_T_76; // @[rawFloatFromFN.scala 66:33]
  wire [9:0] _T_138 = {1'b0,$signed(_T_130)}; // @[rawFloatFromFN.scala 70:48]
  wire  hi_lo_2 = ~_T_131; // @[rawFloatFromFN.scala 72:29]
  wire [22:0] lo_2 = _T_75 ? _T_124 : io_b[22:0]; // @[rawFloatFromFN.scala 72:42]
  wire [24:0] _T_139 = {1'h0,hi_lo_2,lo_2}; // @[Cat.scala 30:58]
  wire [2:0] _T_141 = _T_131 ? 3'h0 : _T_138[8:6]; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_9 = {{2'd0}, _T_135}; // @[recFNFromFN.scala 48:79]
  wire [2:0] hi_lo_3 = _T_141 | _GEN_9; // @[recFNFromFN.scala 48:79]
  wire [5:0] lo_hi_1 = _T_138[5:0]; // @[recFNFromFN.scala 50:23]
  wire [22:0] lo_lo_1 = _T_139[22:0]; // @[recFNFromFN.scala 51:22]
  wire [28:0] lo_3 = {lo_hi_1,lo_lo_1}; // @[Cat.scala 30:58]
  wire [3:0] hi_3 = {io_b[31],hi_lo_3}; // @[Cat.scala 30:58]
  CompareRecFN compareRecFN ( // @[ValExec_CompareRecFN.scala 59:30]
    .io_a(compareRecFN_io_a),
    .io_b(compareRecFN_io_b),
    .io_lt(compareRecFN_io_lt),
    .io_eq(compareRecFN_io_eq)
  );
  assign io_actual_out = compareRecFN_io_lt; // @[ValExec_CompareRecFN.scala 64:19]
  assign compareRecFN_io_a = {hi_1,lo_1}; // @[Cat.scala 30:58]
  assign compareRecFN_io_b = {hi_3,lo_3}; // @[Cat.scala 30:58]
endmodule
module ray_AABB_1(
  input         clock,
  input         reset,
  input  [31:0] io_ray_idir_x,
  input  [31:0] io_ray_idir_y,
  input  [31:0] io_ray_idir_z,
  input  [31:0] io_ray_ood_x,
  input  [31:0] io_ray_ood_y,
  input  [31:0] io_ray_ood_z,
  input  [31:0] io_ray_hitT,
  input  [31:0] io_bvh_n0xy_x,
  input  [31:0] io_bvh_n0xy_y,
  input  [31:0] io_bvh_n0xy_z,
  input  [31:0] io_bvh_n0xy_w,
  input  [31:0] io_bvh_n1xy_x,
  input  [31:0] io_bvh_n1xy_y,
  input  [31:0] io_bvh_n1xy_z,
  input  [31:0] io_bvh_n1xy_w,
  input  [31:0] io_bvh_nz_x,
  input  [31:0] io_bvh_nz_y,
  input  [31:0] io_bvh_nz_z,
  input  [31:0] io_bvh_nz_w,
  input  [31:0] io_bvh_temp_x,
  input  [31:0] io_bvh_temp_y,
  input  [31:0] io_rayid,
  input         io_valid_en,
  output [31:0] io_rayid_out,
  output [31:0] io_nodeIdx_0,
  output [31:0] io_nodeIdx_1,
  output [31:0] io_nodeIdx_2,
  output        io_push,
  output        io_pop,
  output        io_leaf,
  output        io_back,
  output [31:0] io_hitT_out,
  output        io_valid_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
`endif // RANDOMIZE_REG_INIT
  wire  FADD_MUL_1_clock; // @[Ray_AABB_1.scala 80:33]
  wire  FADD_MUL_1_reset; // @[Ray_AABB_1.scala 80:33]
  wire [31:0] FADD_MUL_1_io_a; // @[Ray_AABB_1.scala 80:33]
  wire [31:0] FADD_MUL_1_io_b; // @[Ray_AABB_1.scala 80:33]
  wire [31:0] FADD_MUL_1_io_c; // @[Ray_AABB_1.scala 80:33]
  wire [31:0] FADD_MUL_1_io_out; // @[Ray_AABB_1.scala 80:33]
  wire  FADD_MUL_2_clock; // @[Ray_AABB_1.scala 90:33]
  wire  FADD_MUL_2_reset; // @[Ray_AABB_1.scala 90:33]
  wire [31:0] FADD_MUL_2_io_a; // @[Ray_AABB_1.scala 90:33]
  wire [31:0] FADD_MUL_2_io_b; // @[Ray_AABB_1.scala 90:33]
  wire [31:0] FADD_MUL_2_io_c; // @[Ray_AABB_1.scala 90:33]
  wire [31:0] FADD_MUL_2_io_out; // @[Ray_AABB_1.scala 90:33]
  wire  FADD_MUL_3_clock; // @[Ray_AABB_1.scala 100:33]
  wire  FADD_MUL_3_reset; // @[Ray_AABB_1.scala 100:33]
  wire [31:0] FADD_MUL_3_io_a; // @[Ray_AABB_1.scala 100:33]
  wire [31:0] FADD_MUL_3_io_b; // @[Ray_AABB_1.scala 100:33]
  wire [31:0] FADD_MUL_3_io_c; // @[Ray_AABB_1.scala 100:33]
  wire [31:0] FADD_MUL_3_io_out; // @[Ray_AABB_1.scala 100:33]
  wire  FADD_MUL_4_clock; // @[Ray_AABB_1.scala 110:33]
  wire  FADD_MUL_4_reset; // @[Ray_AABB_1.scala 110:33]
  wire [31:0] FADD_MUL_4_io_a; // @[Ray_AABB_1.scala 110:33]
  wire [31:0] FADD_MUL_4_io_b; // @[Ray_AABB_1.scala 110:33]
  wire [31:0] FADD_MUL_4_io_c; // @[Ray_AABB_1.scala 110:33]
  wire [31:0] FADD_MUL_4_io_out; // @[Ray_AABB_1.scala 110:33]
  wire  FADD_MUL_5_clock; // @[Ray_AABB_1.scala 120:33]
  wire  FADD_MUL_5_reset; // @[Ray_AABB_1.scala 120:33]
  wire [31:0] FADD_MUL_5_io_a; // @[Ray_AABB_1.scala 120:33]
  wire [31:0] FADD_MUL_5_io_b; // @[Ray_AABB_1.scala 120:33]
  wire [31:0] FADD_MUL_5_io_c; // @[Ray_AABB_1.scala 120:33]
  wire [31:0] FADD_MUL_5_io_out; // @[Ray_AABB_1.scala 120:33]
  wire  FADD_MUL_6_clock; // @[Ray_AABB_1.scala 130:33]
  wire  FADD_MUL_6_reset; // @[Ray_AABB_1.scala 130:33]
  wire [31:0] FADD_MUL_6_io_a; // @[Ray_AABB_1.scala 130:33]
  wire [31:0] FADD_MUL_6_io_b; // @[Ray_AABB_1.scala 130:33]
  wire [31:0] FADD_MUL_6_io_c; // @[Ray_AABB_1.scala 130:33]
  wire [31:0] FADD_MUL_6_io_out; // @[Ray_AABB_1.scala 130:33]
  wire  FADD_MUL_7_clock; // @[Ray_AABB_1.scala 140:33]
  wire  FADD_MUL_7_reset; // @[Ray_AABB_1.scala 140:33]
  wire [31:0] FADD_MUL_7_io_a; // @[Ray_AABB_1.scala 140:33]
  wire [31:0] FADD_MUL_7_io_b; // @[Ray_AABB_1.scala 140:33]
  wire [31:0] FADD_MUL_7_io_c; // @[Ray_AABB_1.scala 140:33]
  wire [31:0] FADD_MUL_7_io_out; // @[Ray_AABB_1.scala 140:33]
  wire  FADD_MUL_8_clock; // @[Ray_AABB_1.scala 150:33]
  wire  FADD_MUL_8_reset; // @[Ray_AABB_1.scala 150:33]
  wire [31:0] FADD_MUL_8_io_a; // @[Ray_AABB_1.scala 150:33]
  wire [31:0] FADD_MUL_8_io_b; // @[Ray_AABB_1.scala 150:33]
  wire [31:0] FADD_MUL_8_io_c; // @[Ray_AABB_1.scala 150:33]
  wire [31:0] FADD_MUL_8_io_out; // @[Ray_AABB_1.scala 150:33]
  wire  FADD_MUL_9_clock; // @[Ray_AABB_1.scala 160:33]
  wire  FADD_MUL_9_reset; // @[Ray_AABB_1.scala 160:33]
  wire [31:0] FADD_MUL_9_io_a; // @[Ray_AABB_1.scala 160:33]
  wire [31:0] FADD_MUL_9_io_b; // @[Ray_AABB_1.scala 160:33]
  wire [31:0] FADD_MUL_9_io_c; // @[Ray_AABB_1.scala 160:33]
  wire [31:0] FADD_MUL_9_io_out; // @[Ray_AABB_1.scala 160:33]
  wire  FADD_MUL_10_clock; // @[Ray_AABB_1.scala 170:33]
  wire  FADD_MUL_10_reset; // @[Ray_AABB_1.scala 170:33]
  wire [31:0] FADD_MUL_10_io_a; // @[Ray_AABB_1.scala 170:33]
  wire [31:0] FADD_MUL_10_io_b; // @[Ray_AABB_1.scala 170:33]
  wire [31:0] FADD_MUL_10_io_c; // @[Ray_AABB_1.scala 170:33]
  wire [31:0] FADD_MUL_10_io_out; // @[Ray_AABB_1.scala 170:33]
  wire  FADD_MUL_11_clock; // @[Ray_AABB_1.scala 180:33]
  wire  FADD_MUL_11_reset; // @[Ray_AABB_1.scala 180:33]
  wire [31:0] FADD_MUL_11_io_a; // @[Ray_AABB_1.scala 180:33]
  wire [31:0] FADD_MUL_11_io_b; // @[Ray_AABB_1.scala 180:33]
  wire [31:0] FADD_MUL_11_io_c; // @[Ray_AABB_1.scala 180:33]
  wire [31:0] FADD_MUL_11_io_out; // @[Ray_AABB_1.scala 180:33]
  wire  FADD_MUL_12_clock; // @[Ray_AABB_1.scala 190:33]
  wire  FADD_MUL_12_reset; // @[Ray_AABB_1.scala 190:33]
  wire [31:0] FADD_MUL_12_io_a; // @[Ray_AABB_1.scala 190:33]
  wire [31:0] FADD_MUL_12_io_b; // @[Ray_AABB_1.scala 190:33]
  wire [31:0] FADD_MUL_12_io_c; // @[Ray_AABB_1.scala 190:33]
  wire [31:0] FADD_MUL_12_io_out; // @[Ray_AABB_1.scala 190:33]
  wire [31:0] FCMP_1_io_a; // @[Ray_AABB_1.scala 238:24]
  wire [31:0] FCMP_1_io_b; // @[Ray_AABB_1.scala 238:24]
  wire  FCMP_1_io_actual_out; // @[Ray_AABB_1.scala 238:24]
  wire [31:0] FCMP_2_io_a; // @[Ray_AABB_1.scala 253:24]
  wire [31:0] FCMP_2_io_b; // @[Ray_AABB_1.scala 253:24]
  wire  FCMP_2_io_actual_out; // @[Ray_AABB_1.scala 253:24]
  wire [31:0] FCMP_3_io_a; // @[Ray_AABB_1.scala 266:24]
  wire [31:0] FCMP_3_io_b; // @[Ray_AABB_1.scala 266:24]
  wire  FCMP_3_io_actual_out; // @[Ray_AABB_1.scala 266:24]
  wire [31:0] FCMP_4_io_a; // @[Ray_AABB_1.scala 279:24]
  wire [31:0] FCMP_4_io_b; // @[Ray_AABB_1.scala 279:24]
  wire  FCMP_4_io_actual_out; // @[Ray_AABB_1.scala 279:24]
  wire [31:0] FCMP_5_io_a; // @[Ray_AABB_1.scala 292:25]
  wire [31:0] FCMP_5_io_b; // @[Ray_AABB_1.scala 292:25]
  wire  FCMP_5_io_actual_out; // @[Ray_AABB_1.scala 292:25]
  wire [31:0] FCMP_6_io_a; // @[Ray_AABB_1.scala 305:24]
  wire [31:0] FCMP_6_io_b; // @[Ray_AABB_1.scala 305:24]
  wire  FCMP_6_io_actual_out; // @[Ray_AABB_1.scala 305:24]
  wire [31:0] FCMP_7_io_a; // @[Ray_AABB_1.scala 350:24]
  wire [31:0] FCMP_7_io_b; // @[Ray_AABB_1.scala 350:24]
  wire  FCMP_7_io_actual_out; // @[Ray_AABB_1.scala 350:24]
  wire [31:0] FCMP_8_io_a; // @[Ray_AABB_1.scala 361:24]
  wire [31:0] FCMP_8_io_b; // @[Ray_AABB_1.scala 361:24]
  wire  FCMP_8_io_actual_out; // @[Ray_AABB_1.scala 361:24]
  wire [31:0] FCMP_9_io_a; // @[Ray_AABB_1.scala 372:24]
  wire [31:0] FCMP_9_io_b; // @[Ray_AABB_1.scala 372:24]
  wire  FCMP_9_io_actual_out; // @[Ray_AABB_1.scala 372:24]
  wire [31:0] FCMP_10_io_a; // @[Ray_AABB_1.scala 383:25]
  wire [31:0] FCMP_10_io_b; // @[Ray_AABB_1.scala 383:25]
  wire  FCMP_10_io_actual_out; // @[Ray_AABB_1.scala 383:25]
  wire [31:0] FCMP_11_io_a; // @[Ray_AABB_1.scala 394:25]
  wire [31:0] FCMP_11_io_b; // @[Ray_AABB_1.scala 394:25]
  wire  FCMP_11_io_actual_out; // @[Ray_AABB_1.scala 394:25]
  wire [31:0] FCMP_12_io_a; // @[Ray_AABB_1.scala 405:25]
  wire [31:0] FCMP_12_io_b; // @[Ray_AABB_1.scala 405:25]
  wire  FCMP_12_io_actual_out; // @[Ray_AABB_1.scala 405:25]
  wire [31:0] FCMP_13_io_a; // @[Ray_AABB_1.scala 416:25]
  wire [31:0] FCMP_13_io_b; // @[Ray_AABB_1.scala 416:25]
  wire  FCMP_13_io_actual_out; // @[Ray_AABB_1.scala 416:25]
  wire [31:0] FCMP_14_io_a; // @[Ray_AABB_1.scala 427:25]
  wire [31:0] FCMP_14_io_b; // @[Ray_AABB_1.scala 427:25]
  wire  FCMP_14_io_actual_out; // @[Ray_AABB_1.scala 427:25]
  wire [31:0] FCMP_15_io_a; // @[Ray_AABB_1.scala 465:25]
  wire [31:0] FCMP_15_io_b; // @[Ray_AABB_1.scala 465:25]
  wire  FCMP_15_io_actual_out; // @[Ray_AABB_1.scala 465:25]
  wire [31:0] FCMP_16_io_a; // @[Ray_AABB_1.scala 476:25]
  wire [31:0] FCMP_16_io_b; // @[Ray_AABB_1.scala 476:25]
  wire  FCMP_16_io_actual_out; // @[Ray_AABB_1.scala 476:25]
  wire [31:0] FCMP_17_io_a; // @[Ray_AABB_1.scala 487:25]
  wire [31:0] FCMP_17_io_b; // @[Ray_AABB_1.scala 487:25]
  wire  FCMP_17_io_actual_out; // @[Ray_AABB_1.scala 487:25]
  wire [31:0] FCMP_18_io_a; // @[Ray_AABB_1.scala 498:25]
  wire [31:0] FCMP_18_io_b; // @[Ray_AABB_1.scala 498:25]
  wire  FCMP_18_io_actual_out; // @[Ray_AABB_1.scala 498:25]
  wire [31:0] FCMP_19_io_a; // @[Ray_AABB_1.scala 541:25]
  wire [31:0] FCMP_19_io_b; // @[Ray_AABB_1.scala 541:25]
  wire  FCMP_19_io_actual_out; // @[Ray_AABB_1.scala 541:25]
  wire [31:0] FCMP_20_io_a; // @[Ray_AABB_1.scala 554:25]
  wire [31:0] FCMP_20_io_b; // @[Ray_AABB_1.scala 554:25]
  wire  FCMP_20_io_actual_out; // @[Ray_AABB_1.scala 554:25]
  wire [31:0] FCMP_21_io_a; // @[Ray_AABB_1.scala 567:25]
  wire [31:0] FCMP_21_io_b; // @[Ray_AABB_1.scala 567:25]
  wire  FCMP_21_io_actual_out; // @[Ray_AABB_1.scala 567:25]
  reg  traverseChild0; // @[Ray_AABB_1.scala 32:33]
  reg  traverseChild1; // @[Ray_AABB_1.scala 33:33]
  reg [31:0] c0lox; // @[Ray_AABB_1.scala 35:34]
  reg [31:0] c0hix; // @[Ray_AABB_1.scala 36:34]
  reg [31:0] c0loy; // @[Ray_AABB_1.scala 37:34]
  reg [31:0] c0hiy; // @[Ray_AABB_1.scala 38:33]
  reg [31:0] c0loz; // @[Ray_AABB_1.scala 39:34]
  reg [31:0] c0hiz; // @[Ray_AABB_1.scala 40:34]
  reg [31:0] c1lox; // @[Ray_AABB_1.scala 42:34]
  reg [31:0] c1hix; // @[Ray_AABB_1.scala 43:34]
  reg [31:0] c1loy; // @[Ray_AABB_1.scala 44:34]
  reg [31:0] c1hiy; // @[Ray_AABB_1.scala 45:34]
  reg [31:0] c1loz; // @[Ray_AABB_1.scala 46:34]
  reg [31:0] c1hiz; // @[Ray_AABB_1.scala 47:34]
  reg [31:0] rayid_1; // @[Ray_AABB_1.scala 49:32]
  reg [31:0] hitT_1; // @[Ray_AABB_1.scala 50:33]
  reg [31:0] valid_1; // @[Ray_AABB_1.scala 52:32]
  reg [31:0] cidx_0_1; // @[Ray_AABB_1.scala 53:45]
  reg [31:0] cidx_1_1; // @[Ray_AABB_1.scala 54:45]
  reg [31:0] rayid_temp; // @[Ray_AABB_1.scala 62:35]
  reg [31:0] hitT_temp; // @[Ray_AABB_1.scala 63:36]
  reg [31:0] valid_temp; // @[Ray_AABB_1.scala 65:35]
  reg [31:0] cidx_0_temp; // @[Ray_AABB_1.scala 72:48]
  reg [31:0] cidx_1_temp; // @[Ray_AABB_1.scala 73:48]
  wire  hi = ~io_ray_ood_x[31]; // @[common.scala 90:20]
  wire [30:0] lo = io_ray_ood_x[30:0]; // @[common.scala 90:30]
  wire  hi_2 = ~io_ray_ood_y[31]; // @[common.scala 90:20]
  wire [30:0] lo_2 = io_ray_ood_y[30:0]; // @[common.scala 90:30]
  wire  hi_4 = ~io_ray_ood_z[31]; // @[common.scala 90:20]
  wire [30:0] lo_4 = io_ray_ood_z[30:0]; // @[common.scala 90:30]
  reg [31:0] cidx_0_2; // @[Ray_AABB_1.scala 201:45]
  reg [31:0] cidx_1_2; // @[Ray_AABB_1.scala 202:45]
  reg [31:0] rayid_2; // @[Ray_AABB_1.scala 215:32]
  reg [31:0] hitT_2; // @[Ray_AABB_1.scala 216:33]
  reg [31:0] valid_2; // @[Ray_AABB_1.scala 218:32]
  reg [31:0] cmpMin0_1; // @[Ray_AABB_1.scala 225:28]
  reg [31:0] cmpMin0_2; // @[Ray_AABB_1.scala 226:28]
  reg [31:0] cmpMin0_3; // @[Ray_AABB_1.scala 227:28]
  reg [31:0] cmpMax0_1; // @[Ray_AABB_1.scala 228:28]
  reg [31:0] cmpMax0_2; // @[Ray_AABB_1.scala 229:28]
  reg [31:0] cmpMax0_3; // @[Ray_AABB_1.scala 230:28]
  reg [31:0] cmpMin1_1; // @[Ray_AABB_1.scala 231:28]
  reg [31:0] cmpMin1_2; // @[Ray_AABB_1.scala 232:28]
  reg [31:0] cmpMin1_3; // @[Ray_AABB_1.scala 233:28]
  reg [31:0] cmpMax1_1; // @[Ray_AABB_1.scala 234:28]
  reg [31:0] cmpMax1_2; // @[Ray_AABB_1.scala 235:28]
  reg [31:0] cmpMax1_3; // @[Ray_AABB_1.scala 236:28]
  wire  _T_24 = FCMP_1_io_actual_out; // @[Ray_AABB_1.scala 243:47]
  reg [31:0] c0Min_temp_1; // @[Ray_AABB_1.scala 319:31]
  reg [31:0] c0Min_temp_2; // @[Ray_AABB_1.scala 320:31]
  reg [31:0] c0Max_temp_1; // @[Ray_AABB_1.scala 321:31]
  reg [31:0] c0Max_temp_2; // @[Ray_AABB_1.scala 322:31]
  reg [31:0] c1Min_temp_1; // @[Ray_AABB_1.scala 323:31]
  reg [31:0] c1Min_temp_2; // @[Ray_AABB_1.scala 324:31]
  reg [31:0] c1Max_temp_1; // @[Ray_AABB_1.scala 325:31]
  reg [31:0] c1Max_temp_2; // @[Ray_AABB_1.scala 326:31]
  reg [31:0] cidx_0_3; // @[Ray_AABB_1.scala 328:45]
  reg [31:0] cidx_1_3; // @[Ray_AABB_1.scala 329:45]
  reg [31:0] hitT_3; // @[Ray_AABB_1.scala 343:49]
  reg [31:0] rayid_3; // @[Ray_AABB_1.scala 345:48]
  reg  valid_3; // @[Ray_AABB_1.scala 347:49]
  reg [31:0] c0Min; // @[Ray_AABB_1.scala 438:24]
  reg [31:0] c0Max; // @[Ray_AABB_1.scala 439:24]
  reg [31:0] c1Min; // @[Ray_AABB_1.scala 440:24]
  reg [31:0] c1Max; // @[Ray_AABB_1.scala 441:24]
  reg [31:0] cidx_0_4; // @[Ray_AABB_1.scala 443:45]
  reg [31:0] cidx_1_4; // @[Ray_AABB_1.scala 444:45]
  reg [31:0] hitT_4; // @[Ray_AABB_1.scala 458:49]
  reg [31:0] rayid_4; // @[Ray_AABB_1.scala 460:48]
  reg  valid_4; // @[Ray_AABB_1.scala 462:49]
  reg [31:0] rayid_5; // @[Ray_AABB_1.scala 510:48]
  reg [31:0] hitT_5; // @[Ray_AABB_1.scala 512:49]
  reg  valid_5; // @[Ray_AABB_1.scala 514:49]
  reg [31:0] cidx_0_5; // @[Ray_AABB_1.scala 519:45]
  reg [31:0] cidx_1_5; // @[Ray_AABB_1.scala 520:45]
  reg  swp; // @[Ray_AABB_1.scala 526:49]
  wire  _T_47 = FCMP_21_io_actual_out > 1'h0; // @[Ray_AABB_1.scala 572:36]
  wire  _T_48 = ~traverseChild0; // @[Ray_AABB_1.scala 580:10]
  wire  _T_49 = ~traverseChild1; // @[Ray_AABB_1.scala 580:29]
  wire  _T_60 = ~cidx_1_5[31]; // @[common.scala 100:25]
  wire  _T_62 = ~_T_60; // @[Ray_AABB_1.scala 600:32]
  wire [31:0] _GEN_28 = _T_60 ? $signed(cidx_1_5) : $signed(32'sh0); // @[Ray_AABB_1.scala 609:45 Ray_AABB_1.scala 615:29 Ray_AABB_1.scala 624:29]
  wire  _GEN_31 = ~_T_60 ? 1'h0 : _T_60; // @[Ray_AABB_1.scala 600:39 Ray_AABB_1.scala 604:37]
  wire [31:0] _GEN_33 = ~_T_60 ? $signed(32'sh0) : $signed(_GEN_28); // @[Ray_AABB_1.scala 600:39 Ray_AABB_1.scala 606:30]
  wire [31:0] _GEN_34 = ~_T_60 ? $signed(cidx_1_5) : $signed(32'sh0); // @[Ray_AABB_1.scala 600:39 Ray_AABB_1.scala 607:30]
  wire  _GEN_35 = ~_T_60 | _T_60; // @[Ray_AABB_1.scala 600:39 Ray_AABB_1.scala 608:32]
  wire  _T_73 = ~cidx_0_5[31]; // @[common.scala 100:25]
  wire  _T_75 = ~_T_73; // @[Ray_AABB_1.scala 639:32]
  wire [31:0] _GEN_39 = _T_73 ? $signed(cidx_0_5) : $signed(32'sh0); // @[Ray_AABB_1.scala 648:45 Ray_AABB_1.scala 654:33 Ray_AABB_1.scala 663:33]
  wire  _GEN_42 = ~_T_73 ? 1'h0 : _T_73; // @[Ray_AABB_1.scala 639:39 Ray_AABB_1.scala 643:41]
  wire [31:0] _GEN_44 = ~_T_73 ? $signed(32'sh0) : $signed(_GEN_39); // @[Ray_AABB_1.scala 639:39 Ray_AABB_1.scala 645:34]
  wire [31:0] _GEN_45 = ~_T_73 ? $signed(cidx_0_5) : $signed(32'sh0); // @[Ray_AABB_1.scala 639:39 Ray_AABB_1.scala 646:34]
  wire  _GEN_46 = ~_T_73 | _T_73; // @[Ray_AABB_1.scala 639:39 Ray_AABB_1.scala 647:36]
  wire [31:0] _GEN_49 = _T_60 ? $signed(cidx_0_5) : $signed(32'sh0); // @[Ray_AABB_1.scala 678:49 Ray_AABB_1.scala 683:32 Ray_AABB_1.scala 692:32]
  wire [31:0] _GEN_56 = _T_62 ? $signed(cidx_0_5) : $signed(_GEN_49); // @[Ray_AABB_1.scala 669:43 Ray_AABB_1.scala 674:32]
  wire [31:0] _GEN_61 = _T_73 ? $signed(cidx_1_5) : $signed(32'sh0); // @[Ray_AABB_1.scala 707:49 Ray_AABB_1.scala 712:32 Ray_AABB_1.scala 721:32]
  wire [31:0] _GEN_68 = _T_75 ? $signed(cidx_1_5) : $signed(_GEN_61); // @[Ray_AABB_1.scala 698:43 Ray_AABB_1.scala 703:32]
  wire  _GEN_71 = ~swp & valid_5 & _GEN_46; // @[Ray_AABB_1.scala 697:49 Ray_AABB_1.scala 746:38]
  wire  _GEN_73 = ~swp & valid_5 & _T_75; // @[Ray_AABB_1.scala 697:49 Ray_AABB_1.scala 748:41]
  wire  _GEN_74 = ~swp & valid_5 & _GEN_42; // @[Ray_AABB_1.scala 697:49 Ray_AABB_1.scala 749:39]
  wire [31:0] _GEN_75 = ~swp & valid_5 ? $signed(_GEN_68) : $signed(32'sh0); // @[Ray_AABB_1.scala 697:49 Ray_AABB_1.scala 750:32]
  wire [31:0] _GEN_76 = ~swp & valid_5 ? $signed(_GEN_44) : $signed(32'sh0); // @[Ray_AABB_1.scala 697:49 Ray_AABB_1.scala 751:32]
  wire [31:0] _GEN_77 = ~swp & valid_5 ? $signed(_GEN_45) : $signed(32'sh0); // @[Ray_AABB_1.scala 697:49 Ray_AABB_1.scala 752:32]
  wire  _GEN_78 = swp & valid_5 ? _GEN_35 : _GEN_71; // @[Ray_AABB_1.scala 668:43]
  wire  _GEN_80 = swp & valid_5 ? _T_62 : _GEN_73; // @[Ray_AABB_1.scala 668:43]
  wire  _GEN_81 = swp & valid_5 ? _GEN_31 : _GEN_74; // @[Ray_AABB_1.scala 668:43]
  wire [31:0] _GEN_82 = swp & valid_5 ? $signed(_GEN_56) : $signed(_GEN_75); // @[Ray_AABB_1.scala 668:43]
  wire [31:0] _GEN_83 = swp & valid_5 ? $signed(_GEN_33) : $signed(_GEN_76); // @[Ray_AABB_1.scala 668:43]
  wire [31:0] _GEN_84 = swp & valid_5 ? $signed(_GEN_34) : $signed(_GEN_77); // @[Ray_AABB_1.scala 668:43]
  wire  _GEN_85 = traverseChild0 & traverseChild1 & valid_5 & _GEN_78; // @[Ray_AABB_1.scala 667:84 Ray_AABB_1.scala 756:30]
  wire  _GEN_87 = traverseChild0 & traverseChild1 & valid_5 & _GEN_80; // @[Ray_AABB_1.scala 667:84 Ray_AABB_1.scala 758:33]
  wire  _GEN_88 = traverseChild0 & traverseChild1 & valid_5 & _GEN_81; // @[Ray_AABB_1.scala 667:84 Ray_AABB_1.scala 759:31]
  wire [31:0] _GEN_89 = traverseChild0 & traverseChild1 & valid_5 ? $signed(_GEN_82) : $signed(32'sh0); // @[Ray_AABB_1.scala 667:84 Ray_AABB_1.scala 760:24]
  wire [31:0] _GEN_90 = traverseChild0 & traverseChild1 & valid_5 ? $signed(_GEN_83) : $signed(32'sh0); // @[Ray_AABB_1.scala 667:84 Ray_AABB_1.scala 761:24]
  wire [31:0] _GEN_91 = traverseChild0 & traverseChild1 & valid_5 ? $signed(_GEN_84) : $signed(32'sh0); // @[Ray_AABB_1.scala 667:84 Ray_AABB_1.scala 762:24]
  wire  _GEN_92 = traverseChild0 & _T_49 & valid_5 ? _T_75 : _GEN_87; // @[Ray_AABB_1.scala 628:78]
  wire  _GEN_94 = traverseChild0 & _T_49 & valid_5 ? 1'h0 : _GEN_85; // @[Ray_AABB_1.scala 628:78]
  wire  _GEN_95 = traverseChild0 & _T_49 & valid_5 ? _GEN_42 : _GEN_88; // @[Ray_AABB_1.scala 628:78]
  wire [31:0] _GEN_96 = traverseChild0 & _T_49 & valid_5 ? $signed(32'sh0) : $signed(_GEN_89); // @[Ray_AABB_1.scala 628:78]
  wire [31:0] _GEN_97 = traverseChild0 & _T_49 & valid_5 ? $signed(_GEN_44) : $signed(_GEN_90); // @[Ray_AABB_1.scala 628:78]
  wire [31:0] _GEN_98 = traverseChild0 & _T_49 & valid_5 ? $signed(_GEN_45) : $signed(_GEN_91); // @[Ray_AABB_1.scala 628:78]
  wire  _GEN_99 = traverseChild0 & _T_49 & valid_5 ? _GEN_46 : _GEN_85; // @[Ray_AABB_1.scala 628:78]
  wire  _GEN_100 = _T_48 & traverseChild1 & valid_5 ? _T_62 : _GEN_92; // @[Ray_AABB_1.scala 589:74]
  wire  _GEN_102 = _T_48 & traverseChild1 & valid_5 ? 1'h0 : _GEN_94; // @[Ray_AABB_1.scala 589:74]
  wire  _GEN_103 = _T_48 & traverseChild1 & valid_5 ? _GEN_31 : _GEN_95; // @[Ray_AABB_1.scala 589:74]
  wire [31:0] _GEN_104 = _T_48 & traverseChild1 & valid_5 ? $signed(32'sh0) : $signed(_GEN_96); // @[Ray_AABB_1.scala 589:74]
  wire [31:0] _GEN_105 = _T_48 & traverseChild1 & valid_5 ? $signed(_GEN_33) : $signed(_GEN_97); // @[Ray_AABB_1.scala 589:74]
  wire [31:0] _GEN_106 = _T_48 & traverseChild1 & valid_5 ? $signed(_GEN_34) : $signed(_GEN_98); // @[Ray_AABB_1.scala 589:74]
  wire  _GEN_107 = _T_48 & traverseChild1 & valid_5 ? _GEN_35 : _GEN_99; // @[Ray_AABB_1.scala 589:74]
  MY_MULADD FADD_MUL_1 ( // @[Ray_AABB_1.scala 80:33]
    .clock(FADD_MUL_1_clock),
    .reset(FADD_MUL_1_reset),
    .io_a(FADD_MUL_1_io_a),
    .io_b(FADD_MUL_1_io_b),
    .io_c(FADD_MUL_1_io_c),
    .io_out(FADD_MUL_1_io_out)
  );
  MY_MULADD FADD_MUL_2 ( // @[Ray_AABB_1.scala 90:33]
    .clock(FADD_MUL_2_clock),
    .reset(FADD_MUL_2_reset),
    .io_a(FADD_MUL_2_io_a),
    .io_b(FADD_MUL_2_io_b),
    .io_c(FADD_MUL_2_io_c),
    .io_out(FADD_MUL_2_io_out)
  );
  MY_MULADD FADD_MUL_3 ( // @[Ray_AABB_1.scala 100:33]
    .clock(FADD_MUL_3_clock),
    .reset(FADD_MUL_3_reset),
    .io_a(FADD_MUL_3_io_a),
    .io_b(FADD_MUL_3_io_b),
    .io_c(FADD_MUL_3_io_c),
    .io_out(FADD_MUL_3_io_out)
  );
  MY_MULADD FADD_MUL_4 ( // @[Ray_AABB_1.scala 110:33]
    .clock(FADD_MUL_4_clock),
    .reset(FADD_MUL_4_reset),
    .io_a(FADD_MUL_4_io_a),
    .io_b(FADD_MUL_4_io_b),
    .io_c(FADD_MUL_4_io_c),
    .io_out(FADD_MUL_4_io_out)
  );
  MY_MULADD FADD_MUL_5 ( // @[Ray_AABB_1.scala 120:33]
    .clock(FADD_MUL_5_clock),
    .reset(FADD_MUL_5_reset),
    .io_a(FADD_MUL_5_io_a),
    .io_b(FADD_MUL_5_io_b),
    .io_c(FADD_MUL_5_io_c),
    .io_out(FADD_MUL_5_io_out)
  );
  MY_MULADD FADD_MUL_6 ( // @[Ray_AABB_1.scala 130:33]
    .clock(FADD_MUL_6_clock),
    .reset(FADD_MUL_6_reset),
    .io_a(FADD_MUL_6_io_a),
    .io_b(FADD_MUL_6_io_b),
    .io_c(FADD_MUL_6_io_c),
    .io_out(FADD_MUL_6_io_out)
  );
  MY_MULADD FADD_MUL_7 ( // @[Ray_AABB_1.scala 140:33]
    .clock(FADD_MUL_7_clock),
    .reset(FADD_MUL_7_reset),
    .io_a(FADD_MUL_7_io_a),
    .io_b(FADD_MUL_7_io_b),
    .io_c(FADD_MUL_7_io_c),
    .io_out(FADD_MUL_7_io_out)
  );
  MY_MULADD FADD_MUL_8 ( // @[Ray_AABB_1.scala 150:33]
    .clock(FADD_MUL_8_clock),
    .reset(FADD_MUL_8_reset),
    .io_a(FADD_MUL_8_io_a),
    .io_b(FADD_MUL_8_io_b),
    .io_c(FADD_MUL_8_io_c),
    .io_out(FADD_MUL_8_io_out)
  );
  MY_MULADD FADD_MUL_9 ( // @[Ray_AABB_1.scala 160:33]
    .clock(FADD_MUL_9_clock),
    .reset(FADD_MUL_9_reset),
    .io_a(FADD_MUL_9_io_a),
    .io_b(FADD_MUL_9_io_b),
    .io_c(FADD_MUL_9_io_c),
    .io_out(FADD_MUL_9_io_out)
  );
  MY_MULADD FADD_MUL_10 ( // @[Ray_AABB_1.scala 170:33]
    .clock(FADD_MUL_10_clock),
    .reset(FADD_MUL_10_reset),
    .io_a(FADD_MUL_10_io_a),
    .io_b(FADD_MUL_10_io_b),
    .io_c(FADD_MUL_10_io_c),
    .io_out(FADD_MUL_10_io_out)
  );
  MY_MULADD FADD_MUL_11 ( // @[Ray_AABB_1.scala 180:33]
    .clock(FADD_MUL_11_clock),
    .reset(FADD_MUL_11_reset),
    .io_a(FADD_MUL_11_io_a),
    .io_b(FADD_MUL_11_io_b),
    .io_c(FADD_MUL_11_io_c),
    .io_out(FADD_MUL_11_io_out)
  );
  MY_MULADD FADD_MUL_12 ( // @[Ray_AABB_1.scala 190:33]
    .clock(FADD_MUL_12_clock),
    .reset(FADD_MUL_12_reset),
    .io_a(FADD_MUL_12_io_a),
    .io_b(FADD_MUL_12_io_b),
    .io_c(FADD_MUL_12_io_c),
    .io_out(FADD_MUL_12_io_out)
  );
  ValExec_CompareRecF32_le FCMP_1 ( // @[Ray_AABB_1.scala 238:24]
    .io_a(FCMP_1_io_a),
    .io_b(FCMP_1_io_b),
    .io_actual_out(FCMP_1_io_actual_out)
  );
  ValExec_CompareRecF32_le FCMP_2 ( // @[Ray_AABB_1.scala 253:24]
    .io_a(FCMP_2_io_a),
    .io_b(FCMP_2_io_b),
    .io_actual_out(FCMP_2_io_actual_out)
  );
  ValExec_CompareRecF32_le FCMP_3 ( // @[Ray_AABB_1.scala 266:24]
    .io_a(FCMP_3_io_a),
    .io_b(FCMP_3_io_b),
    .io_actual_out(FCMP_3_io_actual_out)
  );
  ValExec_CompareRecF32_le FCMP_4 ( // @[Ray_AABB_1.scala 279:24]
    .io_a(FCMP_4_io_a),
    .io_b(FCMP_4_io_b),
    .io_actual_out(FCMP_4_io_actual_out)
  );
  ValExec_CompareRecF32_le FCMP_5 ( // @[Ray_AABB_1.scala 292:25]
    .io_a(FCMP_5_io_a),
    .io_b(FCMP_5_io_b),
    .io_actual_out(FCMP_5_io_actual_out)
  );
  ValExec_CompareRecF32_le FCMP_6 ( // @[Ray_AABB_1.scala 305:24]
    .io_a(FCMP_6_io_a),
    .io_b(FCMP_6_io_b),
    .io_actual_out(FCMP_6_io_actual_out)
  );
  ValExec_CompareRecF32_le FCMP_7 ( // @[Ray_AABB_1.scala 350:24]
    .io_a(FCMP_7_io_a),
    .io_b(FCMP_7_io_b),
    .io_actual_out(FCMP_7_io_actual_out)
  );
  ValExec_CompareRecF32_le FCMP_8 ( // @[Ray_AABB_1.scala 361:24]
    .io_a(FCMP_8_io_a),
    .io_b(FCMP_8_io_b),
    .io_actual_out(FCMP_8_io_actual_out)
  );
  ValExec_CompareRecF32_le FCMP_9 ( // @[Ray_AABB_1.scala 372:24]
    .io_a(FCMP_9_io_a),
    .io_b(FCMP_9_io_b),
    .io_actual_out(FCMP_9_io_actual_out)
  );
  ValExec_CompareRecF32_le FCMP_10 ( // @[Ray_AABB_1.scala 383:25]
    .io_a(FCMP_10_io_a),
    .io_b(FCMP_10_io_b),
    .io_actual_out(FCMP_10_io_actual_out)
  );
  ValExec_CompareRecF32_le FCMP_11 ( // @[Ray_AABB_1.scala 394:25]
    .io_a(FCMP_11_io_a),
    .io_b(FCMP_11_io_b),
    .io_actual_out(FCMP_11_io_actual_out)
  );
  ValExec_CompareRecF32_le FCMP_12 ( // @[Ray_AABB_1.scala 405:25]
    .io_a(FCMP_12_io_a),
    .io_b(FCMP_12_io_b),
    .io_actual_out(FCMP_12_io_actual_out)
  );
  ValExec_CompareRecF32_le FCMP_13 ( // @[Ray_AABB_1.scala 416:25]
    .io_a(FCMP_13_io_a),
    .io_b(FCMP_13_io_b),
    .io_actual_out(FCMP_13_io_actual_out)
  );
  ValExec_CompareRecF32_le FCMP_14 ( // @[Ray_AABB_1.scala 427:25]
    .io_a(FCMP_14_io_a),
    .io_b(FCMP_14_io_b),
    .io_actual_out(FCMP_14_io_actual_out)
  );
  ValExec_CompareRecF32_le FCMP_15 ( // @[Ray_AABB_1.scala 465:25]
    .io_a(FCMP_15_io_a),
    .io_b(FCMP_15_io_b),
    .io_actual_out(FCMP_15_io_actual_out)
  );
  ValExec_CompareRecF32_le FCMP_16 ( // @[Ray_AABB_1.scala 476:25]
    .io_a(FCMP_16_io_a),
    .io_b(FCMP_16_io_b),
    .io_actual_out(FCMP_16_io_actual_out)
  );
  ValExec_CompareRecF32_le FCMP_17 ( // @[Ray_AABB_1.scala 487:25]
    .io_a(FCMP_17_io_a),
    .io_b(FCMP_17_io_b),
    .io_actual_out(FCMP_17_io_actual_out)
  );
  ValExec_CompareRecF32_le FCMP_18 ( // @[Ray_AABB_1.scala 498:25]
    .io_a(FCMP_18_io_a),
    .io_b(FCMP_18_io_b),
    .io_actual_out(FCMP_18_io_actual_out)
  );
  ValExec_CompareRecF32_lt FCMP_19 ( // @[Ray_AABB_1.scala 541:25]
    .io_a(FCMP_19_io_a),
    .io_b(FCMP_19_io_b),
    .io_actual_out(FCMP_19_io_actual_out)
  );
  ValExec_CompareRecF32_lt FCMP_20 ( // @[Ray_AABB_1.scala 554:25]
    .io_a(FCMP_20_io_a),
    .io_b(FCMP_20_io_b),
    .io_actual_out(FCMP_20_io_actual_out)
  );
  ValExec_CompareRecF32_lt FCMP_21 ( // @[Ray_AABB_1.scala 567:25]
    .io_a(FCMP_21_io_a),
    .io_b(FCMP_21_io_b),
    .io_actual_out(FCMP_21_io_actual_out)
  );
  assign io_rayid_out = rayid_5; // @[Ray_AABB_1.scala 578:47]
  assign io_nodeIdx_0 = ~traverseChild0 & ~traverseChild1 & valid_5 ? $signed(32'sh0) : $signed(_GEN_104); // @[Ray_AABB_1.scala 580:69 Ray_AABB_1.scala 585:26]
  assign io_nodeIdx_1 = ~traverseChild0 & ~traverseChild1 & valid_5 ? $signed(32'sh0) : $signed(_GEN_105); // @[Ray_AABB_1.scala 580:69 Ray_AABB_1.scala 586:26]
  assign io_nodeIdx_2 = ~traverseChild0 & ~traverseChild1 & valid_5 ? $signed(32'sh0) : $signed(_GEN_106); // @[Ray_AABB_1.scala 580:69 Ray_AABB_1.scala 587:26]
  assign io_push = ~traverseChild0 & ~traverseChild1 & valid_5 ? 1'h0 : _GEN_102; // @[Ray_AABB_1.scala 580:69 Ray_AABB_1.scala 582:32]
  assign io_pop = ~traverseChild0 & ~traverseChild1 & valid_5; // @[Ray_AABB_1.scala 580:51]
  assign io_leaf = ~traverseChild0 & ~traverseChild1 & valid_5 ? 1'h0 : _GEN_100; // @[Ray_AABB_1.scala 580:69 Ray_AABB_1.scala 583:35]
  assign io_back = ~traverseChild0 & ~traverseChild1 & valid_5 ? 1'h0 : _GEN_103; // @[Ray_AABB_1.scala 580:69 Ray_AABB_1.scala 584:33]
  assign io_hitT_out = hitT_5; // @[Ray_AABB_1.scala 579:48]
  assign io_valid_out = ~traverseChild0 & ~traverseChild1 & valid_5 | _GEN_107; // @[Ray_AABB_1.scala 580:69 Ray_AABB_1.scala 588:28]
  assign FADD_MUL_1_clock = clock;
  assign FADD_MUL_1_reset = reset;
  assign FADD_MUL_1_io_a = io_bvh_n0xy_x; // @[Ray_AABB_1.scala 81:21]
  assign FADD_MUL_1_io_b = io_ray_idir_x; // @[Ray_AABB_1.scala 82:21]
  assign FADD_MUL_1_io_c = {hi,lo}; // @[Cat.scala 30:58]
  assign FADD_MUL_2_clock = clock;
  assign FADD_MUL_2_reset = reset;
  assign FADD_MUL_2_io_a = io_bvh_n0xy_y; // @[Ray_AABB_1.scala 91:21]
  assign FADD_MUL_2_io_b = io_ray_idir_x; // @[Ray_AABB_1.scala 92:21]
  assign FADD_MUL_2_io_c = {hi,lo}; // @[Cat.scala 30:58]
  assign FADD_MUL_3_clock = clock;
  assign FADD_MUL_3_reset = reset;
  assign FADD_MUL_3_io_a = io_bvh_n0xy_z; // @[Ray_AABB_1.scala 101:21]
  assign FADD_MUL_3_io_b = io_ray_idir_y; // @[Ray_AABB_1.scala 102:21]
  assign FADD_MUL_3_io_c = {hi_2,lo_2}; // @[Cat.scala 30:58]
  assign FADD_MUL_4_clock = clock;
  assign FADD_MUL_4_reset = reset;
  assign FADD_MUL_4_io_a = io_bvh_n0xy_w; // @[Ray_AABB_1.scala 111:21]
  assign FADD_MUL_4_io_b = io_ray_idir_y; // @[Ray_AABB_1.scala 112:21]
  assign FADD_MUL_4_io_c = {hi_2,lo_2}; // @[Cat.scala 30:58]
  assign FADD_MUL_5_clock = clock;
  assign FADD_MUL_5_reset = reset;
  assign FADD_MUL_5_io_a = io_bvh_nz_x; // @[Ray_AABB_1.scala 121:21]
  assign FADD_MUL_5_io_b = io_ray_idir_z; // @[Ray_AABB_1.scala 122:21]
  assign FADD_MUL_5_io_c = {hi_4,lo_4}; // @[Cat.scala 30:58]
  assign FADD_MUL_6_clock = clock;
  assign FADD_MUL_6_reset = reset;
  assign FADD_MUL_6_io_a = io_bvh_nz_y; // @[Ray_AABB_1.scala 131:21]
  assign FADD_MUL_6_io_b = io_ray_idir_z; // @[Ray_AABB_1.scala 132:21]
  assign FADD_MUL_6_io_c = {hi_4,lo_4}; // @[Cat.scala 30:58]
  assign FADD_MUL_7_clock = clock;
  assign FADD_MUL_7_reset = reset;
  assign FADD_MUL_7_io_a = io_bvh_n1xy_x; // @[Ray_AABB_1.scala 141:21]
  assign FADD_MUL_7_io_b = io_ray_idir_x; // @[Ray_AABB_1.scala 142:21]
  assign FADD_MUL_7_io_c = {hi,lo}; // @[Cat.scala 30:58]
  assign FADD_MUL_8_clock = clock;
  assign FADD_MUL_8_reset = reset;
  assign FADD_MUL_8_io_a = io_bvh_n1xy_y; // @[Ray_AABB_1.scala 151:21]
  assign FADD_MUL_8_io_b = io_ray_idir_x; // @[Ray_AABB_1.scala 152:21]
  assign FADD_MUL_8_io_c = {hi,lo}; // @[Cat.scala 30:58]
  assign FADD_MUL_9_clock = clock;
  assign FADD_MUL_9_reset = reset;
  assign FADD_MUL_9_io_a = io_bvh_n1xy_z; // @[Ray_AABB_1.scala 161:21]
  assign FADD_MUL_9_io_b = io_ray_idir_y; // @[Ray_AABB_1.scala 162:21]
  assign FADD_MUL_9_io_c = {hi_2,lo_2}; // @[Cat.scala 30:58]
  assign FADD_MUL_10_clock = clock;
  assign FADD_MUL_10_reset = reset;
  assign FADD_MUL_10_io_a = io_bvh_n1xy_w; // @[Ray_AABB_1.scala 171:22]
  assign FADD_MUL_10_io_b = io_ray_idir_y; // @[Ray_AABB_1.scala 172:22]
  assign FADD_MUL_10_io_c = {hi_2,lo_2}; // @[Cat.scala 30:58]
  assign FADD_MUL_11_clock = clock;
  assign FADD_MUL_11_reset = reset;
  assign FADD_MUL_11_io_a = io_bvh_nz_z; // @[Ray_AABB_1.scala 181:22]
  assign FADD_MUL_11_io_b = io_ray_idir_z; // @[Ray_AABB_1.scala 182:22]
  assign FADD_MUL_11_io_c = {hi_4,lo_4}; // @[Cat.scala 30:58]
  assign FADD_MUL_12_clock = clock;
  assign FADD_MUL_12_reset = reset;
  assign FADD_MUL_12_io_a = io_bvh_nz_w; // @[Ray_AABB_1.scala 191:22]
  assign FADD_MUL_12_io_b = io_ray_idir_z; // @[Ray_AABB_1.scala 192:22]
  assign FADD_MUL_12_io_c = {hi_4,lo_4}; // @[Cat.scala 30:58]
  assign FCMP_1_io_a = c0lox; // @[Ray_AABB_1.scala 239:21]
  assign FCMP_1_io_b = c0hix; // @[Ray_AABB_1.scala 240:21]
  assign FCMP_2_io_a = c0loy; // @[Ray_AABB_1.scala 254:21]
  assign FCMP_2_io_b = c0hiy; // @[Ray_AABB_1.scala 255:21]
  assign FCMP_3_io_a = c0loz; // @[Ray_AABB_1.scala 267:21]
  assign FCMP_3_io_b = c0hiz; // @[Ray_AABB_1.scala 268:21]
  assign FCMP_4_io_a = c1lox; // @[Ray_AABB_1.scala 280:21]
  assign FCMP_4_io_b = c1hix; // @[Ray_AABB_1.scala 281:21]
  assign FCMP_5_io_a = c1loy; // @[Ray_AABB_1.scala 293:21]
  assign FCMP_5_io_b = c1hiy; // @[Ray_AABB_1.scala 294:21]
  assign FCMP_6_io_a = c1loz; // @[Ray_AABB_1.scala 306:21]
  assign FCMP_6_io_b = c1hiz; // @[Ray_AABB_1.scala 307:21]
  assign FCMP_7_io_a = cmpMin0_1; // @[Ray_AABB_1.scala 351:21]
  assign FCMP_7_io_b = cmpMin0_2; // @[Ray_AABB_1.scala 352:21]
  assign FCMP_8_io_a = cmpMin0_3; // @[Ray_AABB_1.scala 362:21]
  assign FCMP_8_io_b = 32'h0; // @[Ray_AABB_1.scala 363:21]
  assign FCMP_9_io_a = cmpMax0_1; // @[Ray_AABB_1.scala 373:21]
  assign FCMP_9_io_b = cmpMax0_2; // @[Ray_AABB_1.scala 374:21]
  assign FCMP_10_io_a = cmpMax0_3; // @[Ray_AABB_1.scala 384:22]
  assign FCMP_10_io_b = hitT_2; // @[Ray_AABB_1.scala 385:22]
  assign FCMP_11_io_a = cmpMin1_1; // @[Ray_AABB_1.scala 395:22]
  assign FCMP_11_io_b = cmpMin1_2; // @[Ray_AABB_1.scala 396:22]
  assign FCMP_12_io_a = cmpMin1_3; // @[Ray_AABB_1.scala 406:22]
  assign FCMP_12_io_b = 32'h0; // @[Ray_AABB_1.scala 407:22]
  assign FCMP_13_io_a = cmpMax1_1; // @[Ray_AABB_1.scala 417:22]
  assign FCMP_13_io_b = cmpMax1_2; // @[Ray_AABB_1.scala 418:22]
  assign FCMP_14_io_a = cmpMax1_3; // @[Ray_AABB_1.scala 428:22]
  assign FCMP_14_io_b = hitT_2; // @[Ray_AABB_1.scala 429:22]
  assign FCMP_15_io_a = c0Min_temp_1; // @[Ray_AABB_1.scala 466:22]
  assign FCMP_15_io_b = c0Min_temp_2; // @[Ray_AABB_1.scala 467:22]
  assign FCMP_16_io_a = c0Max_temp_1; // @[Ray_AABB_1.scala 477:22]
  assign FCMP_16_io_b = c0Max_temp_2; // @[Ray_AABB_1.scala 478:22]
  assign FCMP_17_io_a = c1Min_temp_1; // @[Ray_AABB_1.scala 488:22]
  assign FCMP_17_io_b = c1Min_temp_2; // @[Ray_AABB_1.scala 489:22]
  assign FCMP_18_io_a = c1Max_temp_1; // @[Ray_AABB_1.scala 499:22]
  assign FCMP_18_io_b = c1Max_temp_2; // @[Ray_AABB_1.scala 500:22]
  assign FCMP_19_io_a = c0Max; // @[Ray_AABB_1.scala 542:22]
  assign FCMP_19_io_b = c0Min; // @[Ray_AABB_1.scala 543:22]
  assign FCMP_20_io_a = c1Max; // @[Ray_AABB_1.scala 555:22]
  assign FCMP_20_io_b = c1Min; // @[Ray_AABB_1.scala 556:22]
  assign FCMP_21_io_a = c1Min; // @[Ray_AABB_1.scala 568:22]
  assign FCMP_21_io_b = c0Min; // @[Ray_AABB_1.scala 569:22]
  always @(posedge clock) begin
    if (reset) begin // @[Ray_AABB_1.scala 32:33]
      traverseChild0 <= 1'h0; // @[Ray_AABB_1.scala 32:33]
    end else if (FCMP_19_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 546:42]
      traverseChild0 <= 1'h0; // @[Ray_AABB_1.scala 547:28]
    end else begin
      traverseChild0 <= 1'h1; // @[Ray_AABB_1.scala 549:28]
    end
    if (reset) begin // @[Ray_AABB_1.scala 33:33]
      traverseChild1 <= 1'h0; // @[Ray_AABB_1.scala 33:33]
    end else if (FCMP_20_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 559:42]
      traverseChild1 <= 1'h0; // @[Ray_AABB_1.scala 560:28]
    end else begin
      traverseChild1 <= 1'h1; // @[Ray_AABB_1.scala 562:28]
    end
    if (reset) begin // @[Ray_AABB_1.scala 35:34]
      c0lox <= 32'h0; // @[Ray_AABB_1.scala 35:34]
    end else begin
      c0lox <= FADD_MUL_1_io_out; // @[Ray_AABB_1.scala 88:37]
    end
    if (reset) begin // @[Ray_AABB_1.scala 36:34]
      c0hix <= 32'h0; // @[Ray_AABB_1.scala 36:34]
    end else begin
      c0hix <= FADD_MUL_2_io_out; // @[Ray_AABB_1.scala 98:37]
    end
    if (reset) begin // @[Ray_AABB_1.scala 37:34]
      c0loy <= 32'h0; // @[Ray_AABB_1.scala 37:34]
    end else begin
      c0loy <= FADD_MUL_3_io_out; // @[Ray_AABB_1.scala 108:37]
    end
    if (reset) begin // @[Ray_AABB_1.scala 38:33]
      c0hiy <= 32'h0; // @[Ray_AABB_1.scala 38:33]
    end else begin
      c0hiy <= FADD_MUL_4_io_out; // @[Ray_AABB_1.scala 118:37]
    end
    if (reset) begin // @[Ray_AABB_1.scala 39:34]
      c0loz <= 32'h0; // @[Ray_AABB_1.scala 39:34]
    end else begin
      c0loz <= FADD_MUL_5_io_out; // @[Ray_AABB_1.scala 128:37]
    end
    if (reset) begin // @[Ray_AABB_1.scala 40:34]
      c0hiz <= 32'h0; // @[Ray_AABB_1.scala 40:34]
    end else begin
      c0hiz <= FADD_MUL_6_io_out; // @[Ray_AABB_1.scala 138:37]
    end
    if (reset) begin // @[Ray_AABB_1.scala 42:34]
      c1lox <= 32'h0; // @[Ray_AABB_1.scala 42:34]
    end else begin
      c1lox <= FADD_MUL_7_io_out; // @[Ray_AABB_1.scala 148:37]
    end
    if (reset) begin // @[Ray_AABB_1.scala 43:34]
      c1hix <= 32'h0; // @[Ray_AABB_1.scala 43:34]
    end else begin
      c1hix <= FADD_MUL_8_io_out; // @[Ray_AABB_1.scala 158:37]
    end
    if (reset) begin // @[Ray_AABB_1.scala 44:34]
      c1loy <= 32'h0; // @[Ray_AABB_1.scala 44:34]
    end else begin
      c1loy <= FADD_MUL_9_io_out; // @[Ray_AABB_1.scala 168:37]
    end
    if (reset) begin // @[Ray_AABB_1.scala 45:34]
      c1hiy <= 32'h0; // @[Ray_AABB_1.scala 45:34]
    end else begin
      c1hiy <= FADD_MUL_10_io_out; // @[Ray_AABB_1.scala 178:37]
    end
    if (reset) begin // @[Ray_AABB_1.scala 46:34]
      c1loz <= 32'h0; // @[Ray_AABB_1.scala 46:34]
    end else begin
      c1loz <= FADD_MUL_11_io_out; // @[Ray_AABB_1.scala 188:37]
    end
    if (reset) begin // @[Ray_AABB_1.scala 47:34]
      c1hiz <= 32'h0; // @[Ray_AABB_1.scala 47:34]
    end else begin
      c1hiz <= FADD_MUL_12_io_out; // @[Ray_AABB_1.scala 198:37]
    end
    if (reset) begin // @[Ray_AABB_1.scala 49:32]
      rayid_1 <= 32'h0; // @[Ray_AABB_1.scala 49:32]
    end else begin
      rayid_1 <= io_rayid; // @[Ray_AABB_1.scala 55:41]
    end
    if (reset) begin // @[Ray_AABB_1.scala 50:33]
      hitT_1 <= 32'h0; // @[Ray_AABB_1.scala 50:33]
    end else begin
      hitT_1 <= io_ray_hitT; // @[Ray_AABB_1.scala 57:43]
    end
    if (reset) begin // @[Ray_AABB_1.scala 52:32]
      valid_1 <= 32'h0; // @[Ray_AABB_1.scala 52:32]
    end else begin
      valid_1 <= {{31'd0}, io_valid_en}; // @[Ray_AABB_1.scala 58:42]
    end
    if (reset) begin // @[Ray_AABB_1.scala 53:45]
      cidx_0_1 <= 32'sh0; // @[Ray_AABB_1.scala 53:45]
    end else begin
      cidx_0_1 <= io_bvh_temp_x; // @[Ray_AABB_1.scala 59:44]
    end
    if (reset) begin // @[Ray_AABB_1.scala 54:45]
      cidx_1_1 <= 32'sh0; // @[Ray_AABB_1.scala 54:45]
    end else begin
      cidx_1_1 <= io_bvh_temp_y; // @[Ray_AABB_1.scala 60:44]
    end
    if (reset) begin // @[Ray_AABB_1.scala 62:35]
      rayid_temp <= 32'h0; // @[Ray_AABB_1.scala 62:35]
    end else begin
      rayid_temp <= rayid_1; // @[Ray_AABB_1.scala 69:31]
    end
    if (reset) begin // @[Ray_AABB_1.scala 63:36]
      hitT_temp <= 32'h0; // @[Ray_AABB_1.scala 63:36]
    end else begin
      hitT_temp <= hitT_1; // @[Ray_AABB_1.scala 67:32]
    end
    if (reset) begin // @[Ray_AABB_1.scala 65:35]
      valid_temp <= 32'h0; // @[Ray_AABB_1.scala 65:35]
    end else begin
      valid_temp <= valid_1; // @[Ray_AABB_1.scala 70:32]
    end
    if (reset) begin // @[Ray_AABB_1.scala 72:48]
      cidx_0_temp <= 32'sh0; // @[Ray_AABB_1.scala 72:48]
    end else begin
      cidx_0_temp <= cidx_0_1; // @[Ray_AABB_1.scala 76:41]
    end
    if (reset) begin // @[Ray_AABB_1.scala 73:48]
      cidx_1_temp <= 32'sh0; // @[Ray_AABB_1.scala 73:48]
    end else begin
      cidx_1_temp <= cidx_1_1; // @[Ray_AABB_1.scala 77:41]
    end
    if (reset) begin // @[Ray_AABB_1.scala 201:45]
      cidx_0_2 <= 32'sh0; // @[Ray_AABB_1.scala 201:45]
    end else begin
      cidx_0_2 <= cidx_0_temp; // @[Ray_AABB_1.scala 208:38]
    end
    if (reset) begin // @[Ray_AABB_1.scala 202:45]
      cidx_1_2 <= 32'sh0; // @[Ray_AABB_1.scala 202:45]
    end else begin
      cidx_1_2 <= cidx_1_temp; // @[Ray_AABB_1.scala 209:38]
    end
    if (reset) begin // @[Ray_AABB_1.scala 215:32]
      rayid_2 <= 32'h0; // @[Ray_AABB_1.scala 215:32]
    end else begin
      rayid_2 <= rayid_temp; // @[Ray_AABB_1.scala 222:28]
    end
    if (reset) begin // @[Ray_AABB_1.scala 216:33]
      hitT_2 <= 32'h0; // @[Ray_AABB_1.scala 216:33]
    end else begin
      hitT_2 <= hitT_temp; // @[Ray_AABB_1.scala 220:29]
    end
    if (reset) begin // @[Ray_AABB_1.scala 218:32]
      valid_2 <= 32'h0; // @[Ray_AABB_1.scala 218:32]
    end else begin
      valid_2 <= valid_temp; // @[Ray_AABB_1.scala 223:29]
    end
    if (reset) begin // @[Ray_AABB_1.scala 225:28]
      cmpMin0_1 <= 32'h0; // @[Ray_AABB_1.scala 225:28]
    end else if (FCMP_1_io_actual_out) begin // @[Ray_AABB_1.scala 243:25]
      cmpMin0_1 <= c0lox;
    end else begin
      cmpMin0_1 <= c0hix;
    end
    if (reset) begin // @[Ray_AABB_1.scala 226:28]
      cmpMin0_2 <= 32'h0; // @[Ray_AABB_1.scala 226:28]
    end else if (FCMP_2_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 258:41]
      cmpMin0_2 <= c0loy; // @[Ray_AABB_1.scala 259:23]
    end else begin
      cmpMin0_2 <= c0hiy; // @[Ray_AABB_1.scala 262:23]
    end
    if (reset) begin // @[Ray_AABB_1.scala 227:28]
      cmpMin0_3 <= 32'h0; // @[Ray_AABB_1.scala 227:28]
    end else if (FCMP_3_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 271:41]
      cmpMin0_3 <= c0loz; // @[Ray_AABB_1.scala 272:23]
    end else begin
      cmpMin0_3 <= c0hiz; // @[Ray_AABB_1.scala 275:23]
    end
    if (reset) begin // @[Ray_AABB_1.scala 228:28]
      cmpMax0_1 <= 32'h0; // @[Ray_AABB_1.scala 228:28]
    end else if (_T_24) begin // @[Ray_AABB_1.scala 244:25]
      cmpMax0_1 <= c0hix;
    end else begin
      cmpMax0_1 <= c0lox;
    end
    if (reset) begin // @[Ray_AABB_1.scala 229:28]
      cmpMax0_2 <= 32'h0; // @[Ray_AABB_1.scala 229:28]
    end else if (FCMP_2_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 258:41]
      cmpMax0_2 <= c0hiy; // @[Ray_AABB_1.scala 260:23]
    end else begin
      cmpMax0_2 <= c0loy; // @[Ray_AABB_1.scala 263:23]
    end
    if (reset) begin // @[Ray_AABB_1.scala 230:28]
      cmpMax0_3 <= 32'h0; // @[Ray_AABB_1.scala 230:28]
    end else if (FCMP_3_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 271:41]
      cmpMax0_3 <= c0hiz; // @[Ray_AABB_1.scala 273:23]
    end else begin
      cmpMax0_3 <= c0loz; // @[Ray_AABB_1.scala 276:23]
    end
    if (reset) begin // @[Ray_AABB_1.scala 231:28]
      cmpMin1_1 <= 32'h0; // @[Ray_AABB_1.scala 231:28]
    end else if (FCMP_4_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 284:41]
      cmpMin1_1 <= c1lox; // @[Ray_AABB_1.scala 285:23]
    end else begin
      cmpMin1_1 <= c1hix; // @[Ray_AABB_1.scala 288:23]
    end
    if (reset) begin // @[Ray_AABB_1.scala 232:28]
      cmpMin1_2 <= 32'h0; // @[Ray_AABB_1.scala 232:28]
    end else if (FCMP_5_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 297:41]
      cmpMin1_2 <= c1loy; // @[Ray_AABB_1.scala 298:23]
    end else begin
      cmpMin1_2 <= c1hiy; // @[Ray_AABB_1.scala 301:23]
    end
    if (reset) begin // @[Ray_AABB_1.scala 233:28]
      cmpMin1_3 <= 32'h0; // @[Ray_AABB_1.scala 233:28]
    end else if (FCMP_6_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 310:41]
      cmpMin1_3 <= c1loz; // @[Ray_AABB_1.scala 311:23]
    end else begin
      cmpMin1_3 <= c1hiz; // @[Ray_AABB_1.scala 314:23]
    end
    if (reset) begin // @[Ray_AABB_1.scala 234:28]
      cmpMax1_1 <= 32'h0; // @[Ray_AABB_1.scala 234:28]
    end else if (FCMP_4_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 284:41]
      cmpMax1_1 <= c1hix; // @[Ray_AABB_1.scala 286:23]
    end else begin
      cmpMax1_1 <= c1lox; // @[Ray_AABB_1.scala 289:23]
    end
    if (reset) begin // @[Ray_AABB_1.scala 235:28]
      cmpMax1_2 <= 32'h0; // @[Ray_AABB_1.scala 235:28]
    end else if (FCMP_5_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 297:41]
      cmpMax1_2 <= c1hiy; // @[Ray_AABB_1.scala 299:23]
    end else begin
      cmpMax1_2 <= c1loy; // @[Ray_AABB_1.scala 302:23]
    end
    if (reset) begin // @[Ray_AABB_1.scala 236:28]
      cmpMax1_3 <= 32'h0; // @[Ray_AABB_1.scala 236:28]
    end else if (FCMP_6_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 310:41]
      cmpMax1_3 <= c1hiz; // @[Ray_AABB_1.scala 312:23]
    end else begin
      cmpMax1_3 <= c1loz; // @[Ray_AABB_1.scala 315:23]
    end
    if (reset) begin // @[Ray_AABB_1.scala 319:31]
      c0Min_temp_1 <= 32'h0; // @[Ray_AABB_1.scala 319:31]
    end else if (FCMP_7_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 355:41]
      c0Min_temp_1 <= cmpMin0_2; // @[Ray_AABB_1.scala 356:26]
    end else begin
      c0Min_temp_1 <= cmpMin0_1; // @[Ray_AABB_1.scala 358:26]
    end
    if (reset) begin // @[Ray_AABB_1.scala 320:31]
      c0Min_temp_2 <= 32'h0; // @[Ray_AABB_1.scala 320:31]
    end else if (FCMP_8_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 366:41]
      c0Min_temp_2 <= 32'h0; // @[Ray_AABB_1.scala 367:26]
    end else begin
      c0Min_temp_2 <= cmpMin0_3; // @[Ray_AABB_1.scala 369:26]
    end
    if (reset) begin // @[Ray_AABB_1.scala 321:31]
      c0Max_temp_1 <= 32'h0; // @[Ray_AABB_1.scala 321:31]
    end else if (FCMP_9_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 377:41]
      c0Max_temp_1 <= cmpMax0_1; // @[Ray_AABB_1.scala 378:26]
    end else begin
      c0Max_temp_1 <= cmpMax0_2; // @[Ray_AABB_1.scala 380:26]
    end
    if (reset) begin // @[Ray_AABB_1.scala 322:31]
      c0Max_temp_2 <= 32'h0; // @[Ray_AABB_1.scala 322:31]
    end else if (FCMP_10_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 388:42]
      c0Max_temp_2 <= cmpMax0_3; // @[Ray_AABB_1.scala 389:26]
    end else begin
      c0Max_temp_2 <= hitT_2; // @[Ray_AABB_1.scala 391:26]
    end
    if (reset) begin // @[Ray_AABB_1.scala 323:31]
      c1Min_temp_1 <= 32'h0; // @[Ray_AABB_1.scala 323:31]
    end else if (FCMP_11_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 399:42]
      c1Min_temp_1 <= cmpMin1_2; // @[Ray_AABB_1.scala 400:26]
    end else begin
      c1Min_temp_1 <= cmpMin1_1; // @[Ray_AABB_1.scala 402:26]
    end
    if (reset) begin // @[Ray_AABB_1.scala 324:31]
      c1Min_temp_2 <= 32'h0; // @[Ray_AABB_1.scala 324:31]
    end else if (FCMP_12_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 410:42]
      c1Min_temp_2 <= 32'h0; // @[Ray_AABB_1.scala 411:26]
    end else begin
      c1Min_temp_2 <= cmpMin1_3; // @[Ray_AABB_1.scala 413:26]
    end
    if (reset) begin // @[Ray_AABB_1.scala 325:31]
      c1Max_temp_1 <= 32'h0; // @[Ray_AABB_1.scala 325:31]
    end else if (FCMP_13_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 421:42]
      c1Max_temp_1 <= cmpMax1_1; // @[Ray_AABB_1.scala 422:26]
    end else begin
      c1Max_temp_1 <= cmpMax1_2; // @[Ray_AABB_1.scala 424:26]
    end
    if (reset) begin // @[Ray_AABB_1.scala 326:31]
      c1Max_temp_2 <= 32'h0; // @[Ray_AABB_1.scala 326:31]
    end else if (FCMP_14_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 432:42]
      c1Max_temp_2 <= cmpMax1_3; // @[Ray_AABB_1.scala 433:26]
    end else begin
      c1Max_temp_2 <= hitT_2; // @[Ray_AABB_1.scala 435:26]
    end
    if (reset) begin // @[Ray_AABB_1.scala 328:45]
      cidx_0_3 <= 32'sh0; // @[Ray_AABB_1.scala 328:45]
    end else begin
      cidx_0_3 <= cidx_0_2; // @[Ray_AABB_1.scala 336:38]
    end
    if (reset) begin // @[Ray_AABB_1.scala 329:45]
      cidx_1_3 <= 32'sh0; // @[Ray_AABB_1.scala 329:45]
    end else begin
      cidx_1_3 <= cidx_1_2; // @[Ray_AABB_1.scala 337:38]
    end
    if (reset) begin // @[Ray_AABB_1.scala 343:49]
      hitT_3 <= 32'h0; // @[Ray_AABB_1.scala 343:49]
    end else begin
      hitT_3 <= hitT_2; // @[Ray_AABB_1.scala 344:42]
    end
    if (reset) begin // @[Ray_AABB_1.scala 345:48]
      rayid_3 <= 32'h0; // @[Ray_AABB_1.scala 345:48]
    end else begin
      rayid_3 <= rayid_2; // @[Ray_AABB_1.scala 346:41]
    end
    if (reset) begin // @[Ray_AABB_1.scala 347:49]
      valid_3 <= 1'h0; // @[Ray_AABB_1.scala 347:49]
    end else begin
      valid_3 <= valid_2[0]; // @[Ray_AABB_1.scala 348:41]
    end
    if (reset) begin // @[Ray_AABB_1.scala 438:24]
      c0Min <= 32'h0; // @[Ray_AABB_1.scala 438:24]
    end else if (FCMP_15_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 470:42]
      c0Min <= c0Min_temp_2; // @[Ray_AABB_1.scala 471:19]
    end else begin
      c0Min <= c0Min_temp_1; // @[Ray_AABB_1.scala 473:19]
    end
    if (reset) begin // @[Ray_AABB_1.scala 439:24]
      c0Max <= 32'h0; // @[Ray_AABB_1.scala 439:24]
    end else if (FCMP_16_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 481:42]
      c0Max <= c0Max_temp_1; // @[Ray_AABB_1.scala 482:19]
    end else begin
      c0Max <= c0Max_temp_2; // @[Ray_AABB_1.scala 484:19]
    end
    if (reset) begin // @[Ray_AABB_1.scala 440:24]
      c1Min <= 32'h0; // @[Ray_AABB_1.scala 440:24]
    end else if (FCMP_17_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 492:42]
      c1Min <= c1Min_temp_2; // @[Ray_AABB_1.scala 493:19]
    end else begin
      c1Min <= c1Min_temp_1; // @[Ray_AABB_1.scala 495:19]
    end
    if (reset) begin // @[Ray_AABB_1.scala 441:24]
      c1Max <= 32'h0; // @[Ray_AABB_1.scala 441:24]
    end else if (FCMP_18_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 503:42]
      c1Max <= c1Max_temp_1; // @[Ray_AABB_1.scala 504:19]
    end else begin
      c1Max <= c1Max_temp_2; // @[Ray_AABB_1.scala 506:19]
    end
    if (reset) begin // @[Ray_AABB_1.scala 443:45]
      cidx_0_4 <= 32'sh0; // @[Ray_AABB_1.scala 443:45]
    end else begin
      cidx_0_4 <= cidx_0_3; // @[Ray_AABB_1.scala 451:38]
    end
    if (reset) begin // @[Ray_AABB_1.scala 444:45]
      cidx_1_4 <= 32'sh0; // @[Ray_AABB_1.scala 444:45]
    end else begin
      cidx_1_4 <= cidx_1_3; // @[Ray_AABB_1.scala 452:38]
    end
    if (reset) begin // @[Ray_AABB_1.scala 458:49]
      hitT_4 <= 32'h0; // @[Ray_AABB_1.scala 458:49]
    end else begin
      hitT_4 <= hitT_3; // @[Ray_AABB_1.scala 459:43]
    end
    if (reset) begin // @[Ray_AABB_1.scala 460:48]
      rayid_4 <= 32'h0; // @[Ray_AABB_1.scala 460:48]
    end else begin
      rayid_4 <= rayid_3; // @[Ray_AABB_1.scala 461:42]
    end
    if (reset) begin // @[Ray_AABB_1.scala 462:49]
      valid_4 <= 1'h0; // @[Ray_AABB_1.scala 462:49]
    end else begin
      valid_4 <= valid_3; // @[Ray_AABB_1.scala 463:41]
    end
    if (reset) begin // @[Ray_AABB_1.scala 510:48]
      rayid_5 <= 32'h0; // @[Ray_AABB_1.scala 510:48]
    end else begin
      rayid_5 <= rayid_4; // @[Ray_AABB_1.scala 511:42]
    end
    if (reset) begin // @[Ray_AABB_1.scala 512:49]
      hitT_5 <= 32'h0; // @[Ray_AABB_1.scala 512:49]
    end else begin
      hitT_5 <= hitT_4; // @[Ray_AABB_1.scala 513:42]
    end
    if (reset) begin // @[Ray_AABB_1.scala 514:49]
      valid_5 <= 1'h0; // @[Ray_AABB_1.scala 514:49]
    end else begin
      valid_5 <= valid_4; // @[Ray_AABB_1.scala 515:41]
    end
    if (reset) begin // @[Ray_AABB_1.scala 519:45]
      cidx_0_5 <= 32'sh0; // @[Ray_AABB_1.scala 519:45]
    end else begin
      cidx_0_5 <= cidx_0_4; // @[Ray_AABB_1.scala 531:38]
    end
    if (reset) begin // @[Ray_AABB_1.scala 520:45]
      cidx_1_5 <= 32'sh0; // @[Ray_AABB_1.scala 520:45]
    end else begin
      cidx_1_5 <= cidx_1_4; // @[Ray_AABB_1.scala 532:38]
    end
    if (reset) begin // @[Ray_AABB_1.scala 526:49]
      swp <= 1'h0; // @[Ray_AABB_1.scala 526:49]
    end else begin
      swp <= _T_47;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  traverseChild0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  traverseChild1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  c0lox = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  c0hix = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  c0loy = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  c0hiy = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  c0loz = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  c0hiz = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  c1lox = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  c1hix = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  c1loy = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  c1hiy = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  c1loz = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  c1hiz = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  rayid_1 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  hitT_1 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  valid_1 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  cidx_0_1 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  cidx_1_1 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  rayid_temp = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  hitT_temp = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  valid_temp = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  cidx_0_temp = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  cidx_1_temp = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  cidx_0_2 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  cidx_1_2 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  rayid_2 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  hitT_2 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  valid_2 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  cmpMin0_1 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  cmpMin0_2 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  cmpMin0_3 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  cmpMax0_1 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  cmpMax0_2 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  cmpMax0_3 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  cmpMin1_1 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  cmpMin1_2 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  cmpMin1_3 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  cmpMax1_1 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  cmpMax1_2 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  cmpMax1_3 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  c0Min_temp_1 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  c0Min_temp_2 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  c0Max_temp_1 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  c0Max_temp_2 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  c1Min_temp_1 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  c1Min_temp_2 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  c1Max_temp_1 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  c1Max_temp_2 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  cidx_0_3 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  cidx_1_3 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  hitT_3 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  rayid_3 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  valid_3 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  c0Min = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  c0Max = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  c1Min = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  c1Max = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  cidx_0_4 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  cidx_1_4 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  hitT_4 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  rayid_4 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  valid_4 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  rayid_5 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  hitT_5 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  valid_5 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  cidx_0_5 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  cidx_1_5 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  swp = _RAND_68[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FIFO(
  input         clock,
  input         reset,
  input  [31:0] io_datain,
  output [31:0] io_dataout,
  input         io_wr,
  input         io_rd,
  output        io_empty
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] mem [0:34]; // @[FIFO.scala 23:16]
  wire [31:0] mem_MPORT_data; // @[FIFO.scala 23:16]
  wire [5:0] mem_MPORT_addr; // @[FIFO.scala 23:16]
  wire [31:0] mem_MPORT_3_data; // @[FIFO.scala 23:16]
  wire [5:0] mem_MPORT_3_addr; // @[FIFO.scala 23:16]
  wire [31:0] mem_MPORT_1_data; // @[FIFO.scala 23:16]
  wire [5:0] mem_MPORT_1_addr; // @[FIFO.scala 23:16]
  wire  mem_MPORT_1_mask; // @[FIFO.scala 23:16]
  wire  mem_MPORT_1_en; // @[FIFO.scala 23:16]
  wire [31:0] mem_MPORT_2_data; // @[FIFO.scala 23:16]
  wire [5:0] mem_MPORT_2_addr; // @[FIFO.scala 23:16]
  wire  mem_MPORT_2_mask; // @[FIFO.scala 23:16]
  wire  mem_MPORT_2_en; // @[FIFO.scala 23:16]
  reg [31:0] count; // @[FIFO.scala 22:22]
  reg [31:0] wPointer; // @[FIFO.scala 24:25]
  reg [31:0] rPointer; // @[FIFO.scala 25:25]
  reg [31:0] dataout; // @[FIFO.scala 26:24]
  wire  _T_2 = io_wr & io_rd; // @[FIFO.scala 34:25]
  wire [31:0] _T_7 = rPointer + 32'h1; // @[FIFO.scala 31:46]
  wire [31:0] _T_8 = rPointer == 32'h22 ? 32'h0 : _T_7; // @[FIFO.scala 31:10]
  wire [31:0] _T_12 = wPointer + 32'h1; // @[FIFO.scala 31:46]
  wire [31:0] _T_13 = wPointer == 32'h22 ? 32'h0 : _T_12; // @[FIFO.scala 31:10]
  wire  _GEN_4 = count == 32'h0 ? 1'h0 : 1'h1; // @[FIFO.scala 35:25 FIFO.scala 23:16 FIFO.scala 39:21]
  wire  _T_17 = count < 32'h23; // @[FIFO.scala 48:16]
  wire [31:0] _T_24 = count + 32'h1; // @[FIFO.scala 51:22]
  wire  _T_28 = count > 32'h0; // @[FIFO.scala 55:16]
  wire [31:0] _T_35 = count - 32'h1; // @[FIFO.scala 59:22]
  wire [31:0] _GEN_21 = count > 32'h0 ? $signed(mem_MPORT_3_data) : $signed(32'sh0); // @[FIFO.scala 55:23 FIFO.scala 56:15 FIFO.scala 61:15]
  wire [31:0] _GEN_22 = count > 32'h0 ? _T_8 : rPointer; // @[FIFO.scala 55:23 FIFO.scala 57:16 FIFO.scala 25:25]
  wire [31:0] _GEN_23 = count > 32'h0 ? _T_35 : count; // @[FIFO.scala 55:23 FIFO.scala 59:13 FIFO.scala 22:22]
  wire  _GEN_26 = ~io_wr & io_rd & _T_28; // @[FIFO.scala 54:55 FIFO.scala 23:16]
  wire  _GEN_31 = io_wr & ~io_rd ? 1'h0 : _GEN_26; // @[FIFO.scala 45:55]
  wire  _GEN_34 = io_wr & ~io_rd & _T_17; // @[FIFO.scala 45:55 FIFO.scala 23:16]
  assign mem_MPORT_addr = rPointer[5:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_data = mem[mem_MPORT_addr]; // @[FIFO.scala 23:16]
  `else
  assign mem_MPORT_data = mem_MPORT_addr >= 6'h23 ? _RAND_1[31:0] : mem[mem_MPORT_addr]; // @[FIFO.scala 23:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_3_addr = rPointer[5:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_3_data = mem[mem_MPORT_3_addr]; // @[FIFO.scala 23:16]
  `else
  assign mem_MPORT_3_data = mem_MPORT_3_addr >= 6'h23 ? _RAND_2[31:0] : mem[mem_MPORT_3_addr]; // @[FIFO.scala 23:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_1_data = io_datain;
  assign mem_MPORT_1_addr = wPointer[5:0];
  assign mem_MPORT_1_mask = 1'h1;
  assign mem_MPORT_1_en = _T_2 & _GEN_4;
  assign mem_MPORT_2_data = io_datain;
  assign mem_MPORT_2_addr = wPointer[5:0];
  assign mem_MPORT_2_mask = 1'h1;
  assign mem_MPORT_2_en = _T_2 ? 1'h0 : _GEN_34;
  assign io_dataout = dataout; // @[FIFO.scala 69:14]
  assign io_empty = count == 32'h0; // @[FIFO.scala 71:22]
  always @(posedge clock) begin
    if(mem_MPORT_1_en & mem_MPORT_1_mask) begin
      mem[mem_MPORT_1_addr] <= mem_MPORT_1_data; // @[FIFO.scala 23:16]
    end
    if(mem_MPORT_2_en & mem_MPORT_2_mask) begin
      mem[mem_MPORT_2_addr] <= mem_MPORT_2_data; // @[FIFO.scala 23:16]
    end
    if (reset) begin // @[FIFO.scala 22:22]
      count <= 32'h0; // @[FIFO.scala 22:22]
    end else if (!(io_wr & io_rd)) begin // @[FIFO.scala 34:46]
      if (io_wr & ~io_rd) begin // @[FIFO.scala 45:55]
        if (count < 32'h23) begin // @[FIFO.scala 48:26]
          count <= _T_24; // @[FIFO.scala 51:13]
        end
      end else if (~io_wr & io_rd) begin // @[FIFO.scala 54:55]
        count <= _GEN_23;
      end
    end
    if (reset) begin // @[FIFO.scala 24:25]
      wPointer <= 32'h0; // @[FIFO.scala 24:25]
    end else if (io_wr & io_rd) begin // @[FIFO.scala 34:46]
      if (!(count == 32'h0)) begin // @[FIFO.scala 35:25]
        wPointer <= _T_13; // @[FIFO.scala 43:16]
      end
    end else if (io_wr & ~io_rd) begin // @[FIFO.scala 45:55]
      if (count < 32'h23) begin // @[FIFO.scala 48:26]
        wPointer <= _T_13; // @[FIFO.scala 50:16]
      end
    end
    if (reset) begin // @[FIFO.scala 25:25]
      rPointer <= 32'h0; // @[FIFO.scala 25:25]
    end else if (io_wr & io_rd) begin // @[FIFO.scala 34:46]
      if (!(count == 32'h0)) begin // @[FIFO.scala 35:25]
        if (rPointer == 32'h22) begin // @[FIFO.scala 31:10]
          rPointer <= 32'h0;
        end else begin
          rPointer <= _T_7;
        end
      end
    end else if (!(io_wr & ~io_rd)) begin // @[FIFO.scala 45:55]
      if (~io_wr & io_rd) begin // @[FIFO.scala 54:55]
        rPointer <= _GEN_22;
      end
    end
    if (reset) begin // @[FIFO.scala 26:24]
      dataout <= 32'sh0; // @[FIFO.scala 26:24]
    end else if (io_wr & io_rd) begin // @[FIFO.scala 34:46]
      if (count == 32'h0) begin // @[FIFO.scala 35:25]
        dataout <= io_datain; // @[FIFO.scala 36:17]
      end else begin
        dataout <= mem_MPORT_data; // @[FIFO.scala 39:15]
      end
    end else if (io_wr & ~io_rd) begin // @[FIFO.scala 45:55]
      dataout <= 32'sh0; // @[FIFO.scala 46:13]
    end else if (~io_wr & io_rd) begin // @[FIFO.scala 54:55]
      dataout <= _GEN_21;
    end else begin
      dataout <= 32'sh0; // @[FIFO.scala 65:13]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {1{`RANDOM}};
  _RAND_2 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 35; initvar = initvar+1)
    mem[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  count = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  wPointer = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  rPointer = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  dataout = _RAND_6[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FIFO_0(
  input         clock,
  input         reset,
  input  [31:0] io_datain,
  output [31:0] io_dataout,
  input         io_wr,
  input         io_rd,
  output        io_empty
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] mem [0:34]; // @[FIFO_0.scala 23:16]
  wire [31:0] mem_MPORT_data; // @[FIFO_0.scala 23:16]
  wire [5:0] mem_MPORT_addr; // @[FIFO_0.scala 23:16]
  wire [31:0] mem_MPORT_3_data; // @[FIFO_0.scala 23:16]
  wire [5:0] mem_MPORT_3_addr; // @[FIFO_0.scala 23:16]
  wire [31:0] mem_MPORT_1_data; // @[FIFO_0.scala 23:16]
  wire [5:0] mem_MPORT_1_addr; // @[FIFO_0.scala 23:16]
  wire  mem_MPORT_1_mask; // @[FIFO_0.scala 23:16]
  wire  mem_MPORT_1_en; // @[FIFO_0.scala 23:16]
  wire [31:0] mem_MPORT_2_data; // @[FIFO_0.scala 23:16]
  wire [5:0] mem_MPORT_2_addr; // @[FIFO_0.scala 23:16]
  wire  mem_MPORT_2_mask; // @[FIFO_0.scala 23:16]
  wire  mem_MPORT_2_en; // @[FIFO_0.scala 23:16]
  reg [31:0] count; // @[FIFO_0.scala 22:22]
  reg [31:0] wPointer; // @[FIFO_0.scala 24:25]
  reg [31:0] rPointer; // @[FIFO_0.scala 25:25]
  reg [31:0] dataout; // @[FIFO_0.scala 26:24]
  wire  _T_2 = io_wr & io_rd; // @[FIFO_0.scala 33:25]
  wire [31:0] _T_7 = rPointer + 32'h1; // @[FIFO_0.scala 30:46]
  wire [31:0] _T_8 = rPointer == 32'h22 ? 32'h0 : _T_7; // @[FIFO_0.scala 30:10]
  wire [31:0] _T_12 = wPointer + 32'h1; // @[FIFO_0.scala 30:46]
  wire [31:0] _T_13 = wPointer == 32'h22 ? 32'h0 : _T_12; // @[FIFO_0.scala 30:10]
  wire  _GEN_4 = count == 32'h0 ? 1'h0 : 1'h1; // @[FIFO_0.scala 34:25 FIFO_0.scala 23:16 FIFO_0.scala 38:21]
  wire  _T_17 = count < 32'h23; // @[FIFO_0.scala 47:16]
  wire [31:0] _T_24 = count + 32'h1; // @[FIFO_0.scala 50:22]
  wire  _T_28 = count > 32'h0; // @[FIFO_0.scala 54:16]
  wire [31:0] _T_35 = count - 32'h1; // @[FIFO_0.scala 58:22]
  wire [31:0] _GEN_21 = count > 32'h0 ? mem_MPORT_3_data : 32'h0; // @[FIFO_0.scala 54:23 FIFO_0.scala 55:15 FIFO_0.scala 60:15]
  wire [31:0] _GEN_22 = count > 32'h0 ? _T_8 : rPointer; // @[FIFO_0.scala 54:23 FIFO_0.scala 56:16 FIFO_0.scala 25:25]
  wire [31:0] _GEN_23 = count > 32'h0 ? _T_35 : count; // @[FIFO_0.scala 54:23 FIFO_0.scala 58:13 FIFO_0.scala 22:22]
  wire  _GEN_26 = ~io_wr & io_rd & _T_28; // @[FIFO_0.scala 53:55 FIFO_0.scala 23:16]
  wire  _GEN_31 = io_wr & ~io_rd ? 1'h0 : _GEN_26; // @[FIFO_0.scala 44:55]
  wire  _GEN_34 = io_wr & ~io_rd & _T_17; // @[FIFO_0.scala 44:55 FIFO_0.scala 23:16]
  assign mem_MPORT_addr = rPointer[5:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_data = mem[mem_MPORT_addr]; // @[FIFO_0.scala 23:16]
  `else
  assign mem_MPORT_data = mem_MPORT_addr >= 6'h23 ? _RAND_1[31:0] : mem[mem_MPORT_addr]; // @[FIFO_0.scala 23:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_3_addr = rPointer[5:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_3_data = mem[mem_MPORT_3_addr]; // @[FIFO_0.scala 23:16]
  `else
  assign mem_MPORT_3_data = mem_MPORT_3_addr >= 6'h23 ? _RAND_2[31:0] : mem[mem_MPORT_3_addr]; // @[FIFO_0.scala 23:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_1_data = io_datain;
  assign mem_MPORT_1_addr = wPointer[5:0];
  assign mem_MPORT_1_mask = 1'h1;
  assign mem_MPORT_1_en = _T_2 & _GEN_4;
  assign mem_MPORT_2_data = io_datain;
  assign mem_MPORT_2_addr = wPointer[5:0];
  assign mem_MPORT_2_mask = 1'h1;
  assign mem_MPORT_2_en = _T_2 ? 1'h0 : _GEN_34;
  assign io_dataout = dataout; // @[FIFO_0.scala 68:14]
  assign io_empty = count == 32'h0; // @[FIFO_0.scala 70:22]
  always @(posedge clock) begin
    if(mem_MPORT_1_en & mem_MPORT_1_mask) begin
      mem[mem_MPORT_1_addr] <= mem_MPORT_1_data; // @[FIFO_0.scala 23:16]
    end
    if(mem_MPORT_2_en & mem_MPORT_2_mask) begin
      mem[mem_MPORT_2_addr] <= mem_MPORT_2_data; // @[FIFO_0.scala 23:16]
    end
    if (reset) begin // @[FIFO_0.scala 22:22]
      count <= 32'h0; // @[FIFO_0.scala 22:22]
    end else if (!(io_wr & io_rd)) begin // @[FIFO_0.scala 33:46]
      if (io_wr & ~io_rd) begin // @[FIFO_0.scala 44:55]
        if (count < 32'h23) begin // @[FIFO_0.scala 47:26]
          count <= _T_24; // @[FIFO_0.scala 50:13]
        end
      end else if (~io_wr & io_rd) begin // @[FIFO_0.scala 53:55]
        count <= _GEN_23;
      end
    end
    if (reset) begin // @[FIFO_0.scala 24:25]
      wPointer <= 32'h0; // @[FIFO_0.scala 24:25]
    end else if (io_wr & io_rd) begin // @[FIFO_0.scala 33:46]
      if (!(count == 32'h0)) begin // @[FIFO_0.scala 34:25]
        wPointer <= _T_13; // @[FIFO_0.scala 42:16]
      end
    end else if (io_wr & ~io_rd) begin // @[FIFO_0.scala 44:55]
      if (count < 32'h23) begin // @[FIFO_0.scala 47:26]
        wPointer <= _T_13; // @[FIFO_0.scala 49:16]
      end
    end
    if (reset) begin // @[FIFO_0.scala 25:25]
      rPointer <= 32'h0; // @[FIFO_0.scala 25:25]
    end else if (io_wr & io_rd) begin // @[FIFO_0.scala 33:46]
      if (!(count == 32'h0)) begin // @[FIFO_0.scala 34:25]
        if (rPointer == 32'h22) begin // @[FIFO_0.scala 30:10]
          rPointer <= 32'h0;
        end else begin
          rPointer <= _T_7;
        end
      end
    end else if (!(io_wr & ~io_rd)) begin // @[FIFO_0.scala 44:55]
      if (~io_wr & io_rd) begin // @[FIFO_0.scala 53:55]
        rPointer <= _GEN_22;
      end
    end
    if (reset) begin // @[FIFO_0.scala 26:24]
      dataout <= 32'h0; // @[FIFO_0.scala 26:24]
    end else if (io_wr & io_rd) begin // @[FIFO_0.scala 33:46]
      if (count == 32'h0) begin // @[FIFO_0.scala 34:25]
        dataout <= io_datain; // @[FIFO_0.scala 35:17]
      end else begin
        dataout <= mem_MPORT_data; // @[FIFO_0.scala 38:15]
      end
    end else if (io_wr & ~io_rd) begin // @[FIFO_0.scala 44:55]
      dataout <= 32'h0; // @[FIFO_0.scala 45:13]
    end else if (~io_wr & io_rd) begin // @[FIFO_0.scala 53:55]
      dataout <= _GEN_21;
    end else begin
      dataout <= 32'h0; // @[FIFO_0.scala 64:13]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {1{`RANDOM}};
  _RAND_2 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 35; initvar = initvar+1)
    mem[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  count = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  wPointer = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  rPointer = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  dataout = _RAND_6[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbitration_1(
  input         clock,
  input         reset,
  input  [31:0] io_node_id_0,
  input  [63:0] io_ray_id_0,
  input  [31:0] io_hit_0,
  input         io_valid_0,
  input  [31:0] io_node_id_1,
  input  [31:0] io_ray_id_1,
  input         io_valid_1,
  input  [31:0] io_ray_id_2,
  input         io_valid_2,
  output [31:0] io_node_id_out,
  output [31:0] io_ray_id_out,
  output [31:0] io_hit_out,
  output        io_valid_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  FIFO_A_1_0_node_clock; // @[Arbitration_1_1.scala 29:38]
  wire  FIFO_A_1_0_node_reset; // @[Arbitration_1_1.scala 29:38]
  wire [31:0] FIFO_A_1_0_node_io_datain; // @[Arbitration_1_1.scala 29:38]
  wire [31:0] FIFO_A_1_0_node_io_dataout; // @[Arbitration_1_1.scala 29:38]
  wire  FIFO_A_1_0_node_io_wr; // @[Arbitration_1_1.scala 29:38]
  wire  FIFO_A_1_0_node_io_rd; // @[Arbitration_1_1.scala 29:38]
  wire  FIFO_A_1_0_node_io_empty; // @[Arbitration_1_1.scala 29:38]
  wire  FIFO_A_1_0_ray_clock; // @[Arbitration_1_1.scala 30:41]
  wire  FIFO_A_1_0_ray_reset; // @[Arbitration_1_1.scala 30:41]
  wire [31:0] FIFO_A_1_0_ray_io_datain; // @[Arbitration_1_1.scala 30:41]
  wire [31:0] FIFO_A_1_0_ray_io_dataout; // @[Arbitration_1_1.scala 30:41]
  wire  FIFO_A_1_0_ray_io_wr; // @[Arbitration_1_1.scala 30:41]
  wire  FIFO_A_1_0_ray_io_rd; // @[Arbitration_1_1.scala 30:41]
  wire  FIFO_A_1_0_ray_io_empty; // @[Arbitration_1_1.scala 30:41]
  wire  FIFO_A_1_0_hit_clock; // @[Arbitration_1_1.scala 31:42]
  wire  FIFO_A_1_0_hit_reset; // @[Arbitration_1_1.scala 31:42]
  wire [31:0] FIFO_A_1_0_hit_io_datain; // @[Arbitration_1_1.scala 31:42]
  wire [31:0] FIFO_A_1_0_hit_io_dataout; // @[Arbitration_1_1.scala 31:42]
  wire  FIFO_A_1_0_hit_io_wr; // @[Arbitration_1_1.scala 31:42]
  wire  FIFO_A_1_0_hit_io_rd; // @[Arbitration_1_1.scala 31:42]
  wire  FIFO_A_1_0_hit_io_empty; // @[Arbitration_1_1.scala 31:42]
  wire  FIFO_A_1_1_node_clock; // @[Arbitration_1_1.scala 33:38]
  wire  FIFO_A_1_1_node_reset; // @[Arbitration_1_1.scala 33:38]
  wire [31:0] FIFO_A_1_1_node_io_datain; // @[Arbitration_1_1.scala 33:38]
  wire [31:0] FIFO_A_1_1_node_io_dataout; // @[Arbitration_1_1.scala 33:38]
  wire  FIFO_A_1_1_node_io_wr; // @[Arbitration_1_1.scala 33:38]
  wire  FIFO_A_1_1_node_io_rd; // @[Arbitration_1_1.scala 33:38]
  wire  FIFO_A_1_1_node_io_empty; // @[Arbitration_1_1.scala 33:38]
  wire  FIFO_A_1_1_ray_clock; // @[Arbitration_1_1.scala 34:41]
  wire  FIFO_A_1_1_ray_reset; // @[Arbitration_1_1.scala 34:41]
  wire [31:0] FIFO_A_1_1_ray_io_datain; // @[Arbitration_1_1.scala 34:41]
  wire [31:0] FIFO_A_1_1_ray_io_dataout; // @[Arbitration_1_1.scala 34:41]
  wire  FIFO_A_1_1_ray_io_wr; // @[Arbitration_1_1.scala 34:41]
  wire  FIFO_A_1_1_ray_io_rd; // @[Arbitration_1_1.scala 34:41]
  wire  FIFO_A_1_1_ray_io_empty; // @[Arbitration_1_1.scala 34:41]
  wire  FIFO_A_1_2_node_clock; // @[Arbitration_1_1.scala 36:38]
  wire  FIFO_A_1_2_node_reset; // @[Arbitration_1_1.scala 36:38]
  wire [31:0] FIFO_A_1_2_node_io_datain; // @[Arbitration_1_1.scala 36:38]
  wire [31:0] FIFO_A_1_2_node_io_dataout; // @[Arbitration_1_1.scala 36:38]
  wire  FIFO_A_1_2_node_io_wr; // @[Arbitration_1_1.scala 36:38]
  wire  FIFO_A_1_2_node_io_rd; // @[Arbitration_1_1.scala 36:38]
  wire  FIFO_A_1_2_node_io_empty; // @[Arbitration_1_1.scala 36:38]
  wire  FIFO_A_1_2_ray_clock; // @[Arbitration_1_1.scala 37:41]
  wire  FIFO_A_1_2_ray_reset; // @[Arbitration_1_1.scala 37:41]
  wire [31:0] FIFO_A_1_2_ray_io_datain; // @[Arbitration_1_1.scala 37:41]
  wire [31:0] FIFO_A_1_2_ray_io_dataout; // @[Arbitration_1_1.scala 37:41]
  wire  FIFO_A_1_2_ray_io_wr; // @[Arbitration_1_1.scala 37:41]
  wire  FIFO_A_1_2_ray_io_rd; // @[Arbitration_1_1.scala 37:41]
  wire  FIFO_A_1_2_ray_io_empty; // @[Arbitration_1_1.scala 37:41]
  reg  valid_out_temp; // @[Arbitration_1_1.scala 63:59]
  wire  _T_1 = FIFO_A_1_0_node_io_empty; // @[Arbitration_1_1.scala 78:45]
  wire  _T_3 = FIFO_A_1_0_node_io_empty & ~FIFO_A_1_1_node_io_empty; // @[Arbitration_1_1.scala 78:53]
  wire  _T_8 = _T_1 & FIFO_A_1_1_node_io_empty & ~FIFO_A_1_2_node_io_empty; // @[Arbitration_1_1.scala 91:88]
  wire  _GEN_4 = FIFO_A_1_0_node_io_empty & ~FIFO_A_1_1_node_io_empty ? 1'h0 : _T_8; // @[Arbitration_1_1.scala 78:89 Arbitration_1_1.scala 84:44]
  reg  FIFO_0_empty; // @[Arbitration_1_1.scala 116:58]
  reg  FIFO_1_empty; // @[Arbitration_1_1.scala 117:58]
  reg  FIFO_2_empty; // @[Arbitration_1_1.scala 118:58]
  wire [31:0] _GEN_8 = FIFO_0_empty & FIFO_1_empty & ~FIFO_2_empty ? $signed(FIFO_A_1_2_node_io_dataout) : $signed(32'sh0
    ); // @[Arbitration_1_1.scala 157:85 Arbitration_1_1.scala 158:45 Arbitration_1_1.scala 165:45]
  wire [31:0] _GEN_9 = FIFO_0_empty & FIFO_1_empty & ~FIFO_2_empty ? FIFO_A_1_2_ray_io_dataout : 32'h0; // @[Arbitration_1_1.scala 157:85 Arbitration_1_1.scala 159:48 Arbitration_1_1.scala 166:48]
  wire  _GEN_11 = FIFO_0_empty & FIFO_1_empty & ~FIFO_2_empty & valid_out_temp; // @[Arbitration_1_1.scala 157:85 Arbitration_1_1.scala 162:50 Arbitration_1_1.scala 168:50]
  wire [31:0] _GEN_12 = FIFO_0_empty & ~FIFO_1_empty ? $signed(FIFO_A_1_1_node_io_dataout) : $signed(_GEN_8); // @[Arbitration_1_1.scala 151:63 Arbitration_1_1.scala 152:46]
  wire [31:0] _GEN_13 = FIFO_0_empty & ~FIFO_1_empty ? FIFO_A_1_1_ray_io_dataout : _GEN_9; // @[Arbitration_1_1.scala 151:63 Arbitration_1_1.scala 153:49]
  wire  _GEN_15 = FIFO_0_empty & ~FIFO_1_empty ? valid_out_temp : _GEN_11; // @[Arbitration_1_1.scala 151:63 Arbitration_1_1.scala 155:50]
  FIFO FIFO_A_1_0_node ( // @[Arbitration_1_1.scala 29:38]
    .clock(FIFO_A_1_0_node_clock),
    .reset(FIFO_A_1_0_node_reset),
    .io_datain(FIFO_A_1_0_node_io_datain),
    .io_dataout(FIFO_A_1_0_node_io_dataout),
    .io_wr(FIFO_A_1_0_node_io_wr),
    .io_rd(FIFO_A_1_0_node_io_rd),
    .io_empty(FIFO_A_1_0_node_io_empty)
  );
  FIFO_0 FIFO_A_1_0_ray ( // @[Arbitration_1_1.scala 30:41]
    .clock(FIFO_A_1_0_ray_clock),
    .reset(FIFO_A_1_0_ray_reset),
    .io_datain(FIFO_A_1_0_ray_io_datain),
    .io_dataout(FIFO_A_1_0_ray_io_dataout),
    .io_wr(FIFO_A_1_0_ray_io_wr),
    .io_rd(FIFO_A_1_0_ray_io_rd),
    .io_empty(FIFO_A_1_0_ray_io_empty)
  );
  FIFO_0 FIFO_A_1_0_hit ( // @[Arbitration_1_1.scala 31:42]
    .clock(FIFO_A_1_0_hit_clock),
    .reset(FIFO_A_1_0_hit_reset),
    .io_datain(FIFO_A_1_0_hit_io_datain),
    .io_dataout(FIFO_A_1_0_hit_io_dataout),
    .io_wr(FIFO_A_1_0_hit_io_wr),
    .io_rd(FIFO_A_1_0_hit_io_rd),
    .io_empty(FIFO_A_1_0_hit_io_empty)
  );
  FIFO FIFO_A_1_1_node ( // @[Arbitration_1_1.scala 33:38]
    .clock(FIFO_A_1_1_node_clock),
    .reset(FIFO_A_1_1_node_reset),
    .io_datain(FIFO_A_1_1_node_io_datain),
    .io_dataout(FIFO_A_1_1_node_io_dataout),
    .io_wr(FIFO_A_1_1_node_io_wr),
    .io_rd(FIFO_A_1_1_node_io_rd),
    .io_empty(FIFO_A_1_1_node_io_empty)
  );
  FIFO_0 FIFO_A_1_1_ray ( // @[Arbitration_1_1.scala 34:41]
    .clock(FIFO_A_1_1_ray_clock),
    .reset(FIFO_A_1_1_ray_reset),
    .io_datain(FIFO_A_1_1_ray_io_datain),
    .io_dataout(FIFO_A_1_1_ray_io_dataout),
    .io_wr(FIFO_A_1_1_ray_io_wr),
    .io_rd(FIFO_A_1_1_ray_io_rd),
    .io_empty(FIFO_A_1_1_ray_io_empty)
  );
  FIFO FIFO_A_1_2_node ( // @[Arbitration_1_1.scala 36:38]
    .clock(FIFO_A_1_2_node_clock),
    .reset(FIFO_A_1_2_node_reset),
    .io_datain(FIFO_A_1_2_node_io_datain),
    .io_dataout(FIFO_A_1_2_node_io_dataout),
    .io_wr(FIFO_A_1_2_node_io_wr),
    .io_rd(FIFO_A_1_2_node_io_rd),
    .io_empty(FIFO_A_1_2_node_io_empty)
  );
  FIFO_0 FIFO_A_1_2_ray ( // @[Arbitration_1_1.scala 37:41]
    .clock(FIFO_A_1_2_ray_clock),
    .reset(FIFO_A_1_2_ray_reset),
    .io_datain(FIFO_A_1_2_ray_io_datain),
    .io_dataout(FIFO_A_1_2_ray_io_dataout),
    .io_wr(FIFO_A_1_2_ray_io_wr),
    .io_rd(FIFO_A_1_2_ray_io_rd),
    .io_empty(FIFO_A_1_2_ray_io_empty)
  );
  assign io_node_id_out = ~FIFO_0_empty ? $signed(FIFO_A_1_0_node_io_dataout) : $signed(_GEN_12); // @[Arbitration_1_1.scala 143:35 Arbitration_1_1.scala 144:45]
  assign io_ray_id_out = ~FIFO_0_empty ? FIFO_A_1_0_ray_io_dataout : _GEN_13; // @[Arbitration_1_1.scala 143:35 Arbitration_1_1.scala 145:46]
  assign io_hit_out = ~FIFO_0_empty ? FIFO_A_1_0_hit_io_dataout : 32'h0; // @[Arbitration_1_1.scala 143:35 Arbitration_1_1.scala 147:52]
  assign io_valid_out = ~FIFO_0_empty ? valid_out_temp : _GEN_15; // @[Arbitration_1_1.scala 143:35 Arbitration_1_1.scala 150:50]
  assign FIFO_A_1_0_node_clock = clock;
  assign FIFO_A_1_0_node_reset = reset;
  assign FIFO_A_1_0_node_io_datain = io_node_id_0; // @[Arbitration_1_1.scala 42:40]
  assign FIFO_A_1_0_node_io_wr = io_valid_0; // @[Arbitration_1_1.scala 39:44]
  assign FIFO_A_1_0_node_io_rd = ~FIFO_A_1_0_node_io_empty; // @[Arbitration_1_1.scala 65:39]
  assign FIFO_A_1_0_ray_clock = clock;
  assign FIFO_A_1_0_ray_reset = reset;
  assign FIFO_A_1_0_ray_io_datain = io_ray_id_0[31:0]; // @[Arbitration_1_1.scala 43:43]
  assign FIFO_A_1_0_ray_io_wr = io_valid_0; // @[Arbitration_1_1.scala 40:47]
  assign FIFO_A_1_0_ray_io_rd = ~FIFO_A_1_0_node_io_empty; // @[Arbitration_1_1.scala 65:39]
  assign FIFO_A_1_0_hit_clock = clock;
  assign FIFO_A_1_0_hit_reset = reset;
  assign FIFO_A_1_0_hit_io_datain = io_hit_0; // @[Arbitration_1_1.scala 44:44]
  assign FIFO_A_1_0_hit_io_wr = io_valid_0; // @[Arbitration_1_1.scala 41:48]
  assign FIFO_A_1_0_hit_io_rd = ~FIFO_A_1_0_node_io_empty; // @[Arbitration_1_1.scala 65:39]
  assign FIFO_A_1_1_node_clock = clock;
  assign FIFO_A_1_1_node_reset = reset;
  assign FIFO_A_1_1_node_io_datain = io_node_id_1; // @[Arbitration_1_1.scala 48:40]
  assign FIFO_A_1_1_node_io_wr = io_valid_1; // @[Arbitration_1_1.scala 46:44]
  assign FIFO_A_1_1_node_io_rd = ~FIFO_A_1_0_node_io_empty ? 1'h0 : _T_3; // @[Arbitration_1_1.scala 65:47 Arbitration_1_1.scala 69:44]
  assign FIFO_A_1_1_ray_clock = clock;
  assign FIFO_A_1_1_ray_reset = reset;
  assign FIFO_A_1_1_ray_io_datain = io_ray_id_1; // @[Arbitration_1_1.scala 49:43]
  assign FIFO_A_1_1_ray_io_wr = io_valid_1; // @[Arbitration_1_1.scala 47:47]
  assign FIFO_A_1_1_ray_io_rd = ~FIFO_A_1_0_node_io_empty ? 1'h0 : _T_3; // @[Arbitration_1_1.scala 65:47 Arbitration_1_1.scala 69:44]
  assign FIFO_A_1_2_node_clock = clock;
  assign FIFO_A_1_2_node_reset = reset;
  assign FIFO_A_1_2_node_io_datain = 32'sh0; // @[Arbitration_1_1.scala 53:40]
  assign FIFO_A_1_2_node_io_wr = io_valid_2; // @[Arbitration_1_1.scala 51:44]
  assign FIFO_A_1_2_node_io_rd = ~FIFO_A_1_0_node_io_empty ? 1'h0 : _GEN_4; // @[Arbitration_1_1.scala 65:47 Arbitration_1_1.scala 71:44]
  assign FIFO_A_1_2_ray_clock = clock;
  assign FIFO_A_1_2_ray_reset = reset;
  assign FIFO_A_1_2_ray_io_datain = io_ray_id_2; // @[Arbitration_1_1.scala 54:43]
  assign FIFO_A_1_2_ray_io_wr = io_valid_2; // @[Arbitration_1_1.scala 52:47]
  assign FIFO_A_1_2_ray_io_rd = ~FIFO_A_1_0_node_io_empty ? 1'h0 : _GEN_4; // @[Arbitration_1_1.scala 65:47 Arbitration_1_1.scala 71:44]
  always @(posedge clock) begin
    if (reset) begin // @[Arbitration_1_1.scala 63:59]
      valid_out_temp <= 1'h0; // @[Arbitration_1_1.scala 63:59]
    end else begin
      valid_out_temp <= FIFO_A_1_0_node_io_rd | FIFO_A_1_1_node_io_rd | FIFO_A_1_2_node_io_rd; // @[Arbitration_1_1.scala 139:51]
    end
    if (reset) begin // @[Arbitration_1_1.scala 116:58]
      FIFO_0_empty <= 1'h0; // @[Arbitration_1_1.scala 116:58]
    end else begin
      FIFO_0_empty <= FIFO_A_1_0_node_io_empty; // @[Arbitration_1_1.scala 120:52]
    end
    if (reset) begin // @[Arbitration_1_1.scala 117:58]
      FIFO_1_empty <= 1'h0; // @[Arbitration_1_1.scala 117:58]
    end else begin
      FIFO_1_empty <= FIFO_A_1_1_node_io_empty; // @[Arbitration_1_1.scala 121:52]
    end
    if (reset) begin // @[Arbitration_1_1.scala 118:58]
      FIFO_2_empty <= 1'h0; // @[Arbitration_1_1.scala 118:58]
    end else begin
      FIFO_2_empty <= FIFO_A_1_2_node_io_empty; // @[Arbitration_1_1.scala 122:52]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid_out_temp = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  FIFO_0_empty = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  FIFO_1_empty = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  FIFO_2_empty = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbitration_2_1(
  input         clock,
  input         reset,
  input  [31:0] io_ray_id_2_0,
  input  [31:0] io_hit_2_0,
  input         io_valid_2_0,
  input  [31:0] io_ray_id_2_1,
  input  [31:0] io_hit_2_1,
  input         io_valid_2_1,
  input  [31:0] io_ray_id_2_2,
  input  [31:0] io_hit_2_2,
  input         io_valid_2_2,
  input  [31:0] io_ray_id_2_3,
  input  [31:0] io_hit_2_3,
  input         io_valid_2_3,
  output [31:0] io_ray_id_out,
  output [31:0] io_hit_out,
  output        io_valid_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  FIFO_A_2_0_ray_clock; // @[Arbitration_2_1.scala 38:41]
  wire  FIFO_A_2_0_ray_reset; // @[Arbitration_2_1.scala 38:41]
  wire [31:0] FIFO_A_2_0_ray_io_datain; // @[Arbitration_2_1.scala 38:41]
  wire [31:0] FIFO_A_2_0_ray_io_dataout; // @[Arbitration_2_1.scala 38:41]
  wire  FIFO_A_2_0_ray_io_wr; // @[Arbitration_2_1.scala 38:41]
  wire  FIFO_A_2_0_ray_io_rd; // @[Arbitration_2_1.scala 38:41]
  wire  FIFO_A_2_0_ray_io_empty; // @[Arbitration_2_1.scala 38:41]
  wire  FIFO_A_2_0_hit_clock; // @[Arbitration_2_1.scala 39:42]
  wire  FIFO_A_2_0_hit_reset; // @[Arbitration_2_1.scala 39:42]
  wire [31:0] FIFO_A_2_0_hit_io_datain; // @[Arbitration_2_1.scala 39:42]
  wire [31:0] FIFO_A_2_0_hit_io_dataout; // @[Arbitration_2_1.scala 39:42]
  wire  FIFO_A_2_0_hit_io_wr; // @[Arbitration_2_1.scala 39:42]
  wire  FIFO_A_2_0_hit_io_rd; // @[Arbitration_2_1.scala 39:42]
  wire  FIFO_A_2_0_hit_io_empty; // @[Arbitration_2_1.scala 39:42]
  wire  FIFO_A_2_1_ray_clock; // @[Arbitration_2_1.scala 41:41]
  wire  FIFO_A_2_1_ray_reset; // @[Arbitration_2_1.scala 41:41]
  wire [31:0] FIFO_A_2_1_ray_io_datain; // @[Arbitration_2_1.scala 41:41]
  wire [31:0] FIFO_A_2_1_ray_io_dataout; // @[Arbitration_2_1.scala 41:41]
  wire  FIFO_A_2_1_ray_io_wr; // @[Arbitration_2_1.scala 41:41]
  wire  FIFO_A_2_1_ray_io_rd; // @[Arbitration_2_1.scala 41:41]
  wire  FIFO_A_2_1_ray_io_empty; // @[Arbitration_2_1.scala 41:41]
  wire  FIFO_A_2_1_hit_clock; // @[Arbitration_2_1.scala 42:42]
  wire  FIFO_A_2_1_hit_reset; // @[Arbitration_2_1.scala 42:42]
  wire [31:0] FIFO_A_2_1_hit_io_datain; // @[Arbitration_2_1.scala 42:42]
  wire [31:0] FIFO_A_2_1_hit_io_dataout; // @[Arbitration_2_1.scala 42:42]
  wire  FIFO_A_2_1_hit_io_wr; // @[Arbitration_2_1.scala 42:42]
  wire  FIFO_A_2_1_hit_io_rd; // @[Arbitration_2_1.scala 42:42]
  wire  FIFO_A_2_1_hit_io_empty; // @[Arbitration_2_1.scala 42:42]
  wire  FIFO_A_2_2_ray_clock; // @[Arbitration_2_1.scala 44:41]
  wire  FIFO_A_2_2_ray_reset; // @[Arbitration_2_1.scala 44:41]
  wire [31:0] FIFO_A_2_2_ray_io_datain; // @[Arbitration_2_1.scala 44:41]
  wire [31:0] FIFO_A_2_2_ray_io_dataout; // @[Arbitration_2_1.scala 44:41]
  wire  FIFO_A_2_2_ray_io_wr; // @[Arbitration_2_1.scala 44:41]
  wire  FIFO_A_2_2_ray_io_rd; // @[Arbitration_2_1.scala 44:41]
  wire  FIFO_A_2_2_ray_io_empty; // @[Arbitration_2_1.scala 44:41]
  wire  FIFO_A_2_2_hit_clock; // @[Arbitration_2_1.scala 45:42]
  wire  FIFO_A_2_2_hit_reset; // @[Arbitration_2_1.scala 45:42]
  wire [31:0] FIFO_A_2_2_hit_io_datain; // @[Arbitration_2_1.scala 45:42]
  wire [31:0] FIFO_A_2_2_hit_io_dataout; // @[Arbitration_2_1.scala 45:42]
  wire  FIFO_A_2_2_hit_io_wr; // @[Arbitration_2_1.scala 45:42]
  wire  FIFO_A_2_2_hit_io_rd; // @[Arbitration_2_1.scala 45:42]
  wire  FIFO_A_2_2_hit_io_empty; // @[Arbitration_2_1.scala 45:42]
  wire  FIFO_A_2_3_ray_clock; // @[Arbitration_2_1.scala 47:41]
  wire  FIFO_A_2_3_ray_reset; // @[Arbitration_2_1.scala 47:41]
  wire [31:0] FIFO_A_2_3_ray_io_datain; // @[Arbitration_2_1.scala 47:41]
  wire [31:0] FIFO_A_2_3_ray_io_dataout; // @[Arbitration_2_1.scala 47:41]
  wire  FIFO_A_2_3_ray_io_wr; // @[Arbitration_2_1.scala 47:41]
  wire  FIFO_A_2_3_ray_io_rd; // @[Arbitration_2_1.scala 47:41]
  wire  FIFO_A_2_3_ray_io_empty; // @[Arbitration_2_1.scala 47:41]
  wire  FIFO_A_2_3_hit_clock; // @[Arbitration_2_1.scala 48:42]
  wire  FIFO_A_2_3_hit_reset; // @[Arbitration_2_1.scala 48:42]
  wire [31:0] FIFO_A_2_3_hit_io_datain; // @[Arbitration_2_1.scala 48:42]
  wire [31:0] FIFO_A_2_3_hit_io_dataout; // @[Arbitration_2_1.scala 48:42]
  wire  FIFO_A_2_3_hit_io_wr; // @[Arbitration_2_1.scala 48:42]
  wire  FIFO_A_2_3_hit_io_rd; // @[Arbitration_2_1.scala 48:42]
  wire  FIFO_A_2_3_hit_io_empty; // @[Arbitration_2_1.scala 48:42]
  reg  valid_out_temp; // @[Arbitration_2_1.scala 73:59]
  wire  _T_1 = FIFO_A_2_0_ray_io_empty; // @[Arbitration_2_1.scala 84:44]
  wire  _T_3 = FIFO_A_2_0_ray_io_empty & ~FIFO_A_2_1_ray_io_empty; // @[Arbitration_2_1.scala 84:52]
  wire  _T_6 = _T_1 & FIFO_A_2_1_ray_io_empty; // @[Arbitration_2_1.scala 93:52]
  wire  _T_8 = _T_1 & FIFO_A_2_1_ray_io_empty & ~FIFO_A_2_2_ray_io_empty; // @[Arbitration_2_1.scala 93:86]
  wire  _T_15 = _T_6 & FIFO_A_2_2_ray_io_empty & ~FIFO_A_2_3_ray_io_empty; // @[Arbitration_2_1.scala 102:119]
  wire  _GEN_4 = _T_1 & FIFO_A_2_1_ray_io_empty & ~FIFO_A_2_2_ray_io_empty ? 1'h0 : _T_15; // @[Arbitration_2_1.scala 93:120 Arbitration_2_1.scala 100:47]
  wire  _GEN_7 = FIFO_A_2_0_ray_io_empty & ~FIFO_A_2_1_ray_io_empty ? 1'h0 : _T_8; // @[Arbitration_2_1.scala 84:87 Arbitration_2_1.scala 89:47]
  wire  _GEN_8 = FIFO_A_2_0_ray_io_empty & ~FIFO_A_2_1_ray_io_empty ? 1'h0 : _GEN_4; // @[Arbitration_2_1.scala 84:87 Arbitration_2_1.scala 91:47]
  reg  FIFO_0_empty; // @[Arbitration_2_1.scala 121:58]
  reg  FIFO_1_empty; // @[Arbitration_2_1.scala 122:58]
  reg  FIFO_2_empty; // @[Arbitration_2_1.scala 123:58]
  reg  FIFO_3_empty; // @[Arbitration_2_1.scala 124:58]
  wire  _T_26 = FIFO_0_empty & FIFO_1_empty; // @[Arbitration_2_1.scala 158:40]
  wire [31:0] _GEN_13 = _T_26 & FIFO_2_empty & ~FIFO_3_empty ? FIFO_A_2_3_ray_io_dataout : 32'h0; // @[Arbitration_2_1.scala 162:107 Arbitration_2_1.scala 166:56 Arbitration_2_1.scala 173:60]
  wire [31:0] _GEN_14 = _T_26 & FIFO_2_empty & ~FIFO_3_empty ? FIFO_A_2_3_hit_io_dataout : 32'h0; // @[Arbitration_2_1.scala 162:107 Arbitration_2_1.scala 167:61 Arbitration_2_1.scala 174:64]
  wire  _GEN_15 = _T_26 & FIFO_2_empty & ~FIFO_3_empty & valid_out_temp; // @[Arbitration_2_1.scala 162:107 Arbitration_2_1.scala 168:59 Arbitration_2_1.scala 175:62]
  wire [31:0] _GEN_16 = FIFO_0_empty & FIFO_1_empty & ~FIFO_2_empty ? FIFO_A_2_2_ray_io_dataout : _GEN_13; // @[Arbitration_2_1.scala 158:85 Arbitration_2_1.scala 159:56]
  wire [31:0] _GEN_17 = FIFO_0_empty & FIFO_1_empty & ~FIFO_2_empty ? FIFO_A_2_2_hit_io_dataout : _GEN_14; // @[Arbitration_2_1.scala 158:85 Arbitration_2_1.scala 160:61]
  wire  _GEN_18 = FIFO_0_empty & FIFO_1_empty & ~FIFO_2_empty ? valid_out_temp : _GEN_15; // @[Arbitration_2_1.scala 158:85 Arbitration_2_1.scala 161:59]
  wire [31:0] _GEN_19 = FIFO_0_empty & ~FIFO_1_empty ? FIFO_A_2_1_ray_io_dataout : _GEN_16; // @[Arbitration_2_1.scala 154:63 Arbitration_2_1.scala 155:56]
  wire [31:0] _GEN_20 = FIFO_0_empty & ~FIFO_1_empty ? FIFO_A_2_1_hit_io_dataout : _GEN_17; // @[Arbitration_2_1.scala 154:63 Arbitration_2_1.scala 156:61]
  wire  _GEN_21 = FIFO_0_empty & ~FIFO_1_empty ? valid_out_temp : _GEN_18; // @[Arbitration_2_1.scala 154:63 Arbitration_2_1.scala 157:59]
  FIFO_0 FIFO_A_2_0_ray ( // @[Arbitration_2_1.scala 38:41]
    .clock(FIFO_A_2_0_ray_clock),
    .reset(FIFO_A_2_0_ray_reset),
    .io_datain(FIFO_A_2_0_ray_io_datain),
    .io_dataout(FIFO_A_2_0_ray_io_dataout),
    .io_wr(FIFO_A_2_0_ray_io_wr),
    .io_rd(FIFO_A_2_0_ray_io_rd),
    .io_empty(FIFO_A_2_0_ray_io_empty)
  );
  FIFO_0 FIFO_A_2_0_hit ( // @[Arbitration_2_1.scala 39:42]
    .clock(FIFO_A_2_0_hit_clock),
    .reset(FIFO_A_2_0_hit_reset),
    .io_datain(FIFO_A_2_0_hit_io_datain),
    .io_dataout(FIFO_A_2_0_hit_io_dataout),
    .io_wr(FIFO_A_2_0_hit_io_wr),
    .io_rd(FIFO_A_2_0_hit_io_rd),
    .io_empty(FIFO_A_2_0_hit_io_empty)
  );
  FIFO_0 FIFO_A_2_1_ray ( // @[Arbitration_2_1.scala 41:41]
    .clock(FIFO_A_2_1_ray_clock),
    .reset(FIFO_A_2_1_ray_reset),
    .io_datain(FIFO_A_2_1_ray_io_datain),
    .io_dataout(FIFO_A_2_1_ray_io_dataout),
    .io_wr(FIFO_A_2_1_ray_io_wr),
    .io_rd(FIFO_A_2_1_ray_io_rd),
    .io_empty(FIFO_A_2_1_ray_io_empty)
  );
  FIFO_0 FIFO_A_2_1_hit ( // @[Arbitration_2_1.scala 42:42]
    .clock(FIFO_A_2_1_hit_clock),
    .reset(FIFO_A_2_1_hit_reset),
    .io_datain(FIFO_A_2_1_hit_io_datain),
    .io_dataout(FIFO_A_2_1_hit_io_dataout),
    .io_wr(FIFO_A_2_1_hit_io_wr),
    .io_rd(FIFO_A_2_1_hit_io_rd),
    .io_empty(FIFO_A_2_1_hit_io_empty)
  );
  FIFO_0 FIFO_A_2_2_ray ( // @[Arbitration_2_1.scala 44:41]
    .clock(FIFO_A_2_2_ray_clock),
    .reset(FIFO_A_2_2_ray_reset),
    .io_datain(FIFO_A_2_2_ray_io_datain),
    .io_dataout(FIFO_A_2_2_ray_io_dataout),
    .io_wr(FIFO_A_2_2_ray_io_wr),
    .io_rd(FIFO_A_2_2_ray_io_rd),
    .io_empty(FIFO_A_2_2_ray_io_empty)
  );
  FIFO_0 FIFO_A_2_2_hit ( // @[Arbitration_2_1.scala 45:42]
    .clock(FIFO_A_2_2_hit_clock),
    .reset(FIFO_A_2_2_hit_reset),
    .io_datain(FIFO_A_2_2_hit_io_datain),
    .io_dataout(FIFO_A_2_2_hit_io_dataout),
    .io_wr(FIFO_A_2_2_hit_io_wr),
    .io_rd(FIFO_A_2_2_hit_io_rd),
    .io_empty(FIFO_A_2_2_hit_io_empty)
  );
  FIFO_0 FIFO_A_2_3_ray ( // @[Arbitration_2_1.scala 47:41]
    .clock(FIFO_A_2_3_ray_clock),
    .reset(FIFO_A_2_3_ray_reset),
    .io_datain(FIFO_A_2_3_ray_io_datain),
    .io_dataout(FIFO_A_2_3_ray_io_dataout),
    .io_wr(FIFO_A_2_3_ray_io_wr),
    .io_rd(FIFO_A_2_3_ray_io_rd),
    .io_empty(FIFO_A_2_3_ray_io_empty)
  );
  FIFO_0 FIFO_A_2_3_hit ( // @[Arbitration_2_1.scala 48:42]
    .clock(FIFO_A_2_3_hit_clock),
    .reset(FIFO_A_2_3_hit_reset),
    .io_datain(FIFO_A_2_3_hit_io_datain),
    .io_dataout(FIFO_A_2_3_hit_io_dataout),
    .io_wr(FIFO_A_2_3_hit_io_wr),
    .io_rd(FIFO_A_2_3_hit_io_rd),
    .io_empty(FIFO_A_2_3_hit_io_empty)
  );
  assign io_ray_id_out = ~FIFO_0_empty ? FIFO_A_2_0_ray_io_dataout : _GEN_19; // @[Arbitration_2_1.scala 150:35 Arbitration_2_1.scala 151:55]
  assign io_hit_out = ~FIFO_0_empty ? FIFO_A_2_0_hit_io_dataout : _GEN_20; // @[Arbitration_2_1.scala 150:35 Arbitration_2_1.scala 152:59]
  assign io_valid_out = ~FIFO_0_empty ? valid_out_temp : _GEN_21; // @[Arbitration_2_1.scala 150:35 Arbitration_2_1.scala 153:57]
  assign FIFO_A_2_0_ray_clock = clock;
  assign FIFO_A_2_0_ray_reset = reset;
  assign FIFO_A_2_0_ray_io_datain = io_ray_id_2_0; // @[Arbitration_2_1.scala 52:43]
  assign FIFO_A_2_0_ray_io_wr = io_valid_2_0; // @[Arbitration_2_1.scala 50:47]
  assign FIFO_A_2_0_ray_io_rd = ~FIFO_A_2_0_ray_io_empty; // @[Arbitration_2_1.scala 75:38]
  assign FIFO_A_2_0_hit_clock = clock;
  assign FIFO_A_2_0_hit_reset = reset;
  assign FIFO_A_2_0_hit_io_datain = io_hit_2_0; // @[Arbitration_2_1.scala 53:44]
  assign FIFO_A_2_0_hit_io_wr = io_valid_2_0; // @[Arbitration_2_1.scala 51:48]
  assign FIFO_A_2_0_hit_io_rd = ~FIFO_A_2_0_ray_io_empty; // @[Arbitration_2_1.scala 75:38]
  assign FIFO_A_2_1_ray_clock = clock;
  assign FIFO_A_2_1_ray_reset = reset;
  assign FIFO_A_2_1_ray_io_datain = io_ray_id_2_1; // @[Arbitration_2_1.scala 57:43]
  assign FIFO_A_2_1_ray_io_wr = io_valid_2_1; // @[Arbitration_2_1.scala 55:47]
  assign FIFO_A_2_1_ray_io_rd = ~FIFO_A_2_0_ray_io_empty ? 1'h0 : _T_3; // @[Arbitration_2_1.scala 75:46 Arbitration_2_1.scala 78:47]
  assign FIFO_A_2_1_hit_clock = clock;
  assign FIFO_A_2_1_hit_reset = reset;
  assign FIFO_A_2_1_hit_io_datain = io_hit_2_1; // @[Arbitration_2_1.scala 58:44]
  assign FIFO_A_2_1_hit_io_wr = io_valid_2_1; // @[Arbitration_2_1.scala 56:48]
  assign FIFO_A_2_1_hit_io_rd = ~FIFO_A_2_0_ray_io_empty ? 1'h0 : _T_3; // @[Arbitration_2_1.scala 75:46 Arbitration_2_1.scala 78:47]
  assign FIFO_A_2_2_ray_clock = clock;
  assign FIFO_A_2_2_ray_reset = reset;
  assign FIFO_A_2_2_ray_io_datain = io_ray_id_2_2; // @[Arbitration_2_1.scala 62:43]
  assign FIFO_A_2_2_ray_io_wr = io_valid_2_2; // @[Arbitration_2_1.scala 60:47]
  assign FIFO_A_2_2_ray_io_rd = ~FIFO_A_2_0_ray_io_empty ? 1'h0 : _GEN_7; // @[Arbitration_2_1.scala 75:46 Arbitration_2_1.scala 80:47]
  assign FIFO_A_2_2_hit_clock = clock;
  assign FIFO_A_2_2_hit_reset = reset;
  assign FIFO_A_2_2_hit_io_datain = io_hit_2_2; // @[Arbitration_2_1.scala 63:44]
  assign FIFO_A_2_2_hit_io_wr = io_valid_2_2; // @[Arbitration_2_1.scala 61:48]
  assign FIFO_A_2_2_hit_io_rd = ~FIFO_A_2_0_ray_io_empty ? 1'h0 : _GEN_7; // @[Arbitration_2_1.scala 75:46 Arbitration_2_1.scala 80:47]
  assign FIFO_A_2_3_ray_clock = clock;
  assign FIFO_A_2_3_ray_reset = reset;
  assign FIFO_A_2_3_ray_io_datain = io_ray_id_2_3; // @[Arbitration_2_1.scala 67:43]
  assign FIFO_A_2_3_ray_io_wr = io_valid_2_3; // @[Arbitration_2_1.scala 65:47]
  assign FIFO_A_2_3_ray_io_rd = ~FIFO_A_2_0_ray_io_empty ? 1'h0 : _GEN_8; // @[Arbitration_2_1.scala 75:46 Arbitration_2_1.scala 82:47]
  assign FIFO_A_2_3_hit_clock = clock;
  assign FIFO_A_2_3_hit_reset = reset;
  assign FIFO_A_2_3_hit_io_datain = io_hit_2_3; // @[Arbitration_2_1.scala 68:44]
  assign FIFO_A_2_3_hit_io_wr = io_valid_2_3; // @[Arbitration_2_1.scala 66:48]
  assign FIFO_A_2_3_hit_io_rd = ~FIFO_A_2_0_ray_io_empty ? 1'h0 : _GEN_8; // @[Arbitration_2_1.scala 75:46 Arbitration_2_1.scala 82:47]
  always @(posedge clock) begin
    if (reset) begin // @[Arbitration_2_1.scala 73:59]
      valid_out_temp <= 1'h0; // @[Arbitration_2_1.scala 73:59]
    end else begin
      valid_out_temp <= FIFO_A_2_0_ray_io_rd | FIFO_A_2_1_ray_io_rd | FIFO_A_2_2_ray_io_rd | FIFO_A_2_3_ray_io_rd; // @[Arbitration_2_1.scala 149:51]
    end
    if (reset) begin // @[Arbitration_2_1.scala 121:58]
      FIFO_0_empty <= 1'h0; // @[Arbitration_2_1.scala 121:58]
    end else begin
      FIFO_0_empty <= FIFO_A_2_0_ray_io_empty; // @[Arbitration_2_1.scala 126:52]
    end
    if (reset) begin // @[Arbitration_2_1.scala 122:58]
      FIFO_1_empty <= 1'h0; // @[Arbitration_2_1.scala 122:58]
    end else begin
      FIFO_1_empty <= FIFO_A_2_1_ray_io_empty; // @[Arbitration_2_1.scala 127:52]
    end
    if (reset) begin // @[Arbitration_2_1.scala 123:58]
      FIFO_2_empty <= 1'h0; // @[Arbitration_2_1.scala 123:58]
    end else begin
      FIFO_2_empty <= FIFO_A_2_2_ray_io_empty; // @[Arbitration_2_1.scala 128:52]
    end
    if (reset) begin // @[Arbitration_2_1.scala 124:58]
      FIFO_3_empty <= 1'h0; // @[Arbitration_2_1.scala 124:58]
    end else begin
      FIFO_3_empty <= FIFO_A_2_3_ray_io_empty; // @[Arbitration_2_1.scala 129:52]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid_out_temp = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  FIFO_0_empty = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  FIFO_1_empty = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  FIFO_2_empty = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  FIFO_3_empty = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbitration_3(
  input         clock,
  input         reset,
  input  [31:0] io_node_id_3_0,
  input  [31:0] io_ray_id_3_0,
  input  [31:0] io_hit_3_0,
  input         io_valid_3_0,
  input  [31:0] io_node_id_3_1,
  input  [31:0] io_ray_id_3_1,
  input  [31:0] io_hit_3_1,
  input         io_valid_3_1,
  input  [31:0] io_node_id_3_2,
  input  [31:0] io_ray_id_3_2,
  input  [31:0] io_hit_3_2,
  input         io_valid_3_2,
  input  [31:0] io_node_id_3_3,
  input  [31:0] io_ray_id_3_3,
  input  [31:0] io_hit_3_3,
  input         io_valid_3_3,
  input  [31:0] io_node_id_3_4,
  input  [31:0] io_ray_id_3_4,
  input  [31:0] io_hit_3_4,
  input         io_valid_3_4,
  output [31:0] io_node_id_out,
  output [31:0] io_ray_id_out,
  output [31:0] io_hit_out,
  output        io_valid_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire  FIFO_A_3_0_node_clock; // @[Arbitration_3.scala 42:38]
  wire  FIFO_A_3_0_node_reset; // @[Arbitration_3.scala 42:38]
  wire [31:0] FIFO_A_3_0_node_io_datain; // @[Arbitration_3.scala 42:38]
  wire [31:0] FIFO_A_3_0_node_io_dataout; // @[Arbitration_3.scala 42:38]
  wire  FIFO_A_3_0_node_io_wr; // @[Arbitration_3.scala 42:38]
  wire  FIFO_A_3_0_node_io_rd; // @[Arbitration_3.scala 42:38]
  wire  FIFO_A_3_0_node_io_empty; // @[Arbitration_3.scala 42:38]
  wire  FIFO_A_3_0_ray_clock; // @[Arbitration_3.scala 43:41]
  wire  FIFO_A_3_0_ray_reset; // @[Arbitration_3.scala 43:41]
  wire [31:0] FIFO_A_3_0_ray_io_datain; // @[Arbitration_3.scala 43:41]
  wire [31:0] FIFO_A_3_0_ray_io_dataout; // @[Arbitration_3.scala 43:41]
  wire  FIFO_A_3_0_ray_io_wr; // @[Arbitration_3.scala 43:41]
  wire  FIFO_A_3_0_ray_io_rd; // @[Arbitration_3.scala 43:41]
  wire  FIFO_A_3_0_ray_io_empty; // @[Arbitration_3.scala 43:41]
  wire  FIFO_A_3_0_hit_clock; // @[Arbitration_3.scala 44:42]
  wire  FIFO_A_3_0_hit_reset; // @[Arbitration_3.scala 44:42]
  wire [31:0] FIFO_A_3_0_hit_io_datain; // @[Arbitration_3.scala 44:42]
  wire [31:0] FIFO_A_3_0_hit_io_dataout; // @[Arbitration_3.scala 44:42]
  wire  FIFO_A_3_0_hit_io_wr; // @[Arbitration_3.scala 44:42]
  wire  FIFO_A_3_0_hit_io_rd; // @[Arbitration_3.scala 44:42]
  wire  FIFO_A_3_0_hit_io_empty; // @[Arbitration_3.scala 44:42]
  wire  FIFO_A_3_1_node_clock; // @[Arbitration_3.scala 46:38]
  wire  FIFO_A_3_1_node_reset; // @[Arbitration_3.scala 46:38]
  wire [31:0] FIFO_A_3_1_node_io_datain; // @[Arbitration_3.scala 46:38]
  wire [31:0] FIFO_A_3_1_node_io_dataout; // @[Arbitration_3.scala 46:38]
  wire  FIFO_A_3_1_node_io_wr; // @[Arbitration_3.scala 46:38]
  wire  FIFO_A_3_1_node_io_rd; // @[Arbitration_3.scala 46:38]
  wire  FIFO_A_3_1_node_io_empty; // @[Arbitration_3.scala 46:38]
  wire  FIFO_A_3_1_ray_clock; // @[Arbitration_3.scala 47:41]
  wire  FIFO_A_3_1_ray_reset; // @[Arbitration_3.scala 47:41]
  wire [31:0] FIFO_A_3_1_ray_io_datain; // @[Arbitration_3.scala 47:41]
  wire [31:0] FIFO_A_3_1_ray_io_dataout; // @[Arbitration_3.scala 47:41]
  wire  FIFO_A_3_1_ray_io_wr; // @[Arbitration_3.scala 47:41]
  wire  FIFO_A_3_1_ray_io_rd; // @[Arbitration_3.scala 47:41]
  wire  FIFO_A_3_1_ray_io_empty; // @[Arbitration_3.scala 47:41]
  wire  FIFO_A_3_1_hit_clock; // @[Arbitration_3.scala 48:42]
  wire  FIFO_A_3_1_hit_reset; // @[Arbitration_3.scala 48:42]
  wire [31:0] FIFO_A_3_1_hit_io_datain; // @[Arbitration_3.scala 48:42]
  wire [31:0] FIFO_A_3_1_hit_io_dataout; // @[Arbitration_3.scala 48:42]
  wire  FIFO_A_3_1_hit_io_wr; // @[Arbitration_3.scala 48:42]
  wire  FIFO_A_3_1_hit_io_rd; // @[Arbitration_3.scala 48:42]
  wire  FIFO_A_3_1_hit_io_empty; // @[Arbitration_3.scala 48:42]
  wire  FIFO_A_3_2_node_clock; // @[Arbitration_3.scala 50:38]
  wire  FIFO_A_3_2_node_reset; // @[Arbitration_3.scala 50:38]
  wire [31:0] FIFO_A_3_2_node_io_datain; // @[Arbitration_3.scala 50:38]
  wire [31:0] FIFO_A_3_2_node_io_dataout; // @[Arbitration_3.scala 50:38]
  wire  FIFO_A_3_2_node_io_wr; // @[Arbitration_3.scala 50:38]
  wire  FIFO_A_3_2_node_io_rd; // @[Arbitration_3.scala 50:38]
  wire  FIFO_A_3_2_node_io_empty; // @[Arbitration_3.scala 50:38]
  wire  FIFO_A_3_2_ray_clock; // @[Arbitration_3.scala 51:41]
  wire  FIFO_A_3_2_ray_reset; // @[Arbitration_3.scala 51:41]
  wire [31:0] FIFO_A_3_2_ray_io_datain; // @[Arbitration_3.scala 51:41]
  wire [31:0] FIFO_A_3_2_ray_io_dataout; // @[Arbitration_3.scala 51:41]
  wire  FIFO_A_3_2_ray_io_wr; // @[Arbitration_3.scala 51:41]
  wire  FIFO_A_3_2_ray_io_rd; // @[Arbitration_3.scala 51:41]
  wire  FIFO_A_3_2_ray_io_empty; // @[Arbitration_3.scala 51:41]
  wire  FIFO_A_3_2_hit_clock; // @[Arbitration_3.scala 52:42]
  wire  FIFO_A_3_2_hit_reset; // @[Arbitration_3.scala 52:42]
  wire [31:0] FIFO_A_3_2_hit_io_datain; // @[Arbitration_3.scala 52:42]
  wire [31:0] FIFO_A_3_2_hit_io_dataout; // @[Arbitration_3.scala 52:42]
  wire  FIFO_A_3_2_hit_io_wr; // @[Arbitration_3.scala 52:42]
  wire  FIFO_A_3_2_hit_io_rd; // @[Arbitration_3.scala 52:42]
  wire  FIFO_A_3_2_hit_io_empty; // @[Arbitration_3.scala 52:42]
  wire  FIFO_A_3_3_node_clock; // @[Arbitration_3.scala 54:38]
  wire  FIFO_A_3_3_node_reset; // @[Arbitration_3.scala 54:38]
  wire [31:0] FIFO_A_3_3_node_io_datain; // @[Arbitration_3.scala 54:38]
  wire [31:0] FIFO_A_3_3_node_io_dataout; // @[Arbitration_3.scala 54:38]
  wire  FIFO_A_3_3_node_io_wr; // @[Arbitration_3.scala 54:38]
  wire  FIFO_A_3_3_node_io_rd; // @[Arbitration_3.scala 54:38]
  wire  FIFO_A_3_3_node_io_empty; // @[Arbitration_3.scala 54:38]
  wire  FIFO_A_3_3_ray_clock; // @[Arbitration_3.scala 55:41]
  wire  FIFO_A_3_3_ray_reset; // @[Arbitration_3.scala 55:41]
  wire [31:0] FIFO_A_3_3_ray_io_datain; // @[Arbitration_3.scala 55:41]
  wire [31:0] FIFO_A_3_3_ray_io_dataout; // @[Arbitration_3.scala 55:41]
  wire  FIFO_A_3_3_ray_io_wr; // @[Arbitration_3.scala 55:41]
  wire  FIFO_A_3_3_ray_io_rd; // @[Arbitration_3.scala 55:41]
  wire  FIFO_A_3_3_ray_io_empty; // @[Arbitration_3.scala 55:41]
  wire  FIFO_A_3_3_hit_clock; // @[Arbitration_3.scala 56:42]
  wire  FIFO_A_3_3_hit_reset; // @[Arbitration_3.scala 56:42]
  wire [31:0] FIFO_A_3_3_hit_io_datain; // @[Arbitration_3.scala 56:42]
  wire [31:0] FIFO_A_3_3_hit_io_dataout; // @[Arbitration_3.scala 56:42]
  wire  FIFO_A_3_3_hit_io_wr; // @[Arbitration_3.scala 56:42]
  wire  FIFO_A_3_3_hit_io_rd; // @[Arbitration_3.scala 56:42]
  wire  FIFO_A_3_3_hit_io_empty; // @[Arbitration_3.scala 56:42]
  wire  FIFO_A_3_4_node_clock; // @[Arbitration_3.scala 58:38]
  wire  FIFO_A_3_4_node_reset; // @[Arbitration_3.scala 58:38]
  wire [31:0] FIFO_A_3_4_node_io_datain; // @[Arbitration_3.scala 58:38]
  wire [31:0] FIFO_A_3_4_node_io_dataout; // @[Arbitration_3.scala 58:38]
  wire  FIFO_A_3_4_node_io_wr; // @[Arbitration_3.scala 58:38]
  wire  FIFO_A_3_4_node_io_rd; // @[Arbitration_3.scala 58:38]
  wire  FIFO_A_3_4_node_io_empty; // @[Arbitration_3.scala 58:38]
  wire  FIFO_A_3_4_ray_clock; // @[Arbitration_3.scala 59:41]
  wire  FIFO_A_3_4_ray_reset; // @[Arbitration_3.scala 59:41]
  wire [31:0] FIFO_A_3_4_ray_io_datain; // @[Arbitration_3.scala 59:41]
  wire [31:0] FIFO_A_3_4_ray_io_dataout; // @[Arbitration_3.scala 59:41]
  wire  FIFO_A_3_4_ray_io_wr; // @[Arbitration_3.scala 59:41]
  wire  FIFO_A_3_4_ray_io_rd; // @[Arbitration_3.scala 59:41]
  wire  FIFO_A_3_4_ray_io_empty; // @[Arbitration_3.scala 59:41]
  wire  FIFO_A_3_4_hit_clock; // @[Arbitration_3.scala 60:42]
  wire  FIFO_A_3_4_hit_reset; // @[Arbitration_3.scala 60:42]
  wire [31:0] FIFO_A_3_4_hit_io_datain; // @[Arbitration_3.scala 60:42]
  wire [31:0] FIFO_A_3_4_hit_io_dataout; // @[Arbitration_3.scala 60:42]
  wire  FIFO_A_3_4_hit_io_wr; // @[Arbitration_3.scala 60:42]
  wire  FIFO_A_3_4_hit_io_rd; // @[Arbitration_3.scala 60:42]
  wire  FIFO_A_3_4_hit_io_empty; // @[Arbitration_3.scala 60:42]
  reg  valid_out_temp; // @[Arbitration_3.scala 101:59]
  wire  _T_1 = FIFO_A_3_0_node_io_empty; // @[Arbitration_3.scala 119:45]
  wire  _T_3 = FIFO_A_3_0_node_io_empty & ~FIFO_A_3_1_node_io_empty; // @[Arbitration_3.scala 119:53]
  wire  _T_6 = _T_1 & FIFO_A_3_1_node_io_empty; // @[Arbitration_3.scala 135:53]
  wire  _T_8 = _T_1 & FIFO_A_3_1_node_io_empty & ~FIFO_A_3_2_node_io_empty; // @[Arbitration_3.scala 135:88]
  wire  _T_13 = _T_6 & FIFO_A_3_2_node_io_empty; // @[Arbitration_3.scala 151:88]
  wire  _T_15 = _T_6 & FIFO_A_3_2_node_io_empty & ~FIFO_A_3_3_node_io_empty; // @[Arbitration_3.scala 151:123]
  wire  _T_24 = _T_13 & FIFO_A_3_3_node_io_empty & ~FIFO_A_3_4_node_io_empty; // @[Arbitration_3.scala 167:157]
  wire  _GEN_4 = _T_6 & FIFO_A_3_2_node_io_empty & ~FIFO_A_3_3_node_io_empty ? 1'h0 : _T_24; // @[Arbitration_3.scala 151:158 Arbitration_3.scala 164:44]
  wire  _GEN_7 = _T_1 & FIFO_A_3_1_node_io_empty & ~FIFO_A_3_2_node_io_empty ? 1'h0 : _T_15; // @[Arbitration_3.scala 135:124 Arbitration_3.scala 145:44]
  wire  _GEN_8 = _T_1 & FIFO_A_3_1_node_io_empty & ~FIFO_A_3_2_node_io_empty ? 1'h0 : _GEN_4; // @[Arbitration_3.scala 135:124 Arbitration_3.scala 148:44]
  wire  _GEN_11 = FIFO_A_3_0_node_io_empty & ~FIFO_A_3_1_node_io_empty ? 1'h0 : _T_8; // @[Arbitration_3.scala 119:89 Arbitration_3.scala 126:44]
  wire  _GEN_12 = FIFO_A_3_0_node_io_empty & ~FIFO_A_3_1_node_io_empty ? 1'h0 : _GEN_7; // @[Arbitration_3.scala 119:89 Arbitration_3.scala 129:44]
  wire  _GEN_13 = FIFO_A_3_0_node_io_empty & ~FIFO_A_3_1_node_io_empty ? 1'h0 : _GEN_8; // @[Arbitration_3.scala 119:89 Arbitration_3.scala 132:44]
  reg  FIFO_0_empty; // @[Arbitration_3.scala 200:58]
  reg  FIFO_1_empty; // @[Arbitration_3.scala 201:58]
  reg  FIFO_2_empty; // @[Arbitration_3.scala 202:58]
  reg  FIFO_3_empty; // @[Arbitration_3.scala 203:58]
  reg  FIFO_4_empty; // @[Arbitration_3.scala 204:58]
  wire  _T_36 = FIFO_0_empty & FIFO_1_empty; // @[Arbitration_3.scala 237:40]
  wire  _T_43 = _T_36 & FIFO_2_empty; // @[Arbitration_3.scala 242:62]
  wire [31:0] _GEN_19 = _T_43 & FIFO_3_empty & ~FIFO_4_empty ? $signed(FIFO_A_3_4_node_io_dataout) : $signed(32'sh0); // @[Arbitration_3.scala 247:129 Arbitration_3.scala 248:46 Arbitration_3.scala 253:46]
  wire [31:0] _GEN_20 = _T_43 & FIFO_3_empty & ~FIFO_4_empty ? FIFO_A_3_4_ray_io_dataout : 32'h0; // @[Arbitration_3.scala 247:129 Arbitration_3.scala 249:48 Arbitration_3.scala 254:48]
  wire [31:0] _GEN_21 = _T_43 & FIFO_3_empty & ~FIFO_4_empty ? FIFO_A_3_4_hit_io_dataout : 32'h0; // @[Arbitration_3.scala 247:129 Arbitration_3.scala 250:52 Arbitration_3.scala 255:53]
  wire  _GEN_22 = _T_43 & FIFO_3_empty & ~FIFO_4_empty & valid_out_temp; // @[Arbitration_3.scala 247:129 Arbitration_3.scala 251:50 Arbitration_3.scala 256:50]
  wire [31:0] _GEN_23 = _T_36 & FIFO_2_empty & ~FIFO_3_empty ? $signed(FIFO_A_3_3_node_io_dataout) : $signed(_GEN_19); // @[Arbitration_3.scala 242:107 Arbitration_3.scala 243:46]
  wire [31:0] _GEN_24 = _T_36 & FIFO_2_empty & ~FIFO_3_empty ? FIFO_A_3_3_ray_io_dataout : _GEN_20; // @[Arbitration_3.scala 242:107 Arbitration_3.scala 244:47]
  wire [31:0] _GEN_25 = _T_36 & FIFO_2_empty & ~FIFO_3_empty ? FIFO_A_3_3_hit_io_dataout : _GEN_21; // @[Arbitration_3.scala 242:107 Arbitration_3.scala 245:53]
  wire  _GEN_26 = _T_36 & FIFO_2_empty & ~FIFO_3_empty ? valid_out_temp : _GEN_22; // @[Arbitration_3.scala 242:107 Arbitration_3.scala 246:50]
  wire [31:0] _GEN_27 = FIFO_0_empty & FIFO_1_empty & ~FIFO_2_empty ? $signed(FIFO_A_3_2_node_io_dataout) : $signed(
    _GEN_23); // @[Arbitration_3.scala 237:85 Arbitration_3.scala 238:46]
  wire [31:0] _GEN_28 = FIFO_0_empty & FIFO_1_empty & ~FIFO_2_empty ? FIFO_A_3_2_ray_io_dataout : _GEN_24; // @[Arbitration_3.scala 237:85 Arbitration_3.scala 239:48]
  wire [31:0] _GEN_29 = FIFO_0_empty & FIFO_1_empty & ~FIFO_2_empty ? FIFO_A_3_2_hit_io_dataout : _GEN_25; // @[Arbitration_3.scala 237:85 Arbitration_3.scala 240:53]
  wire  _GEN_30 = FIFO_0_empty & FIFO_1_empty & ~FIFO_2_empty ? valid_out_temp : _GEN_26; // @[Arbitration_3.scala 237:85 Arbitration_3.scala 241:50]
  wire [31:0] _GEN_31 = FIFO_0_empty & ~FIFO_1_empty ? $signed(FIFO_A_3_1_node_io_dataout) : $signed(_GEN_27); // @[Arbitration_3.scala 232:63 Arbitration_3.scala 233:45]
  wire [31:0] _GEN_32 = FIFO_0_empty & ~FIFO_1_empty ? FIFO_A_3_1_ray_io_dataout : _GEN_28; // @[Arbitration_3.scala 232:63 Arbitration_3.scala 234:48]
  wire [31:0] _GEN_33 = FIFO_0_empty & ~FIFO_1_empty ? FIFO_A_3_1_hit_io_dataout : _GEN_29; // @[Arbitration_3.scala 232:63 Arbitration_3.scala 235:53]
  wire  _GEN_34 = FIFO_0_empty & ~FIFO_1_empty ? valid_out_temp : _GEN_30; // @[Arbitration_3.scala 232:63 Arbitration_3.scala 236:50]
  FIFO FIFO_A_3_0_node ( // @[Arbitration_3.scala 42:38]
    .clock(FIFO_A_3_0_node_clock),
    .reset(FIFO_A_3_0_node_reset),
    .io_datain(FIFO_A_3_0_node_io_datain),
    .io_dataout(FIFO_A_3_0_node_io_dataout),
    .io_wr(FIFO_A_3_0_node_io_wr),
    .io_rd(FIFO_A_3_0_node_io_rd),
    .io_empty(FIFO_A_3_0_node_io_empty)
  );
  FIFO_0 FIFO_A_3_0_ray ( // @[Arbitration_3.scala 43:41]
    .clock(FIFO_A_3_0_ray_clock),
    .reset(FIFO_A_3_0_ray_reset),
    .io_datain(FIFO_A_3_0_ray_io_datain),
    .io_dataout(FIFO_A_3_0_ray_io_dataout),
    .io_wr(FIFO_A_3_0_ray_io_wr),
    .io_rd(FIFO_A_3_0_ray_io_rd),
    .io_empty(FIFO_A_3_0_ray_io_empty)
  );
  FIFO_0 FIFO_A_3_0_hit ( // @[Arbitration_3.scala 44:42]
    .clock(FIFO_A_3_0_hit_clock),
    .reset(FIFO_A_3_0_hit_reset),
    .io_datain(FIFO_A_3_0_hit_io_datain),
    .io_dataout(FIFO_A_3_0_hit_io_dataout),
    .io_wr(FIFO_A_3_0_hit_io_wr),
    .io_rd(FIFO_A_3_0_hit_io_rd),
    .io_empty(FIFO_A_3_0_hit_io_empty)
  );
  FIFO FIFO_A_3_1_node ( // @[Arbitration_3.scala 46:38]
    .clock(FIFO_A_3_1_node_clock),
    .reset(FIFO_A_3_1_node_reset),
    .io_datain(FIFO_A_3_1_node_io_datain),
    .io_dataout(FIFO_A_3_1_node_io_dataout),
    .io_wr(FIFO_A_3_1_node_io_wr),
    .io_rd(FIFO_A_3_1_node_io_rd),
    .io_empty(FIFO_A_3_1_node_io_empty)
  );
  FIFO_0 FIFO_A_3_1_ray ( // @[Arbitration_3.scala 47:41]
    .clock(FIFO_A_3_1_ray_clock),
    .reset(FIFO_A_3_1_ray_reset),
    .io_datain(FIFO_A_3_1_ray_io_datain),
    .io_dataout(FIFO_A_3_1_ray_io_dataout),
    .io_wr(FIFO_A_3_1_ray_io_wr),
    .io_rd(FIFO_A_3_1_ray_io_rd),
    .io_empty(FIFO_A_3_1_ray_io_empty)
  );
  FIFO_0 FIFO_A_3_1_hit ( // @[Arbitration_3.scala 48:42]
    .clock(FIFO_A_3_1_hit_clock),
    .reset(FIFO_A_3_1_hit_reset),
    .io_datain(FIFO_A_3_1_hit_io_datain),
    .io_dataout(FIFO_A_3_1_hit_io_dataout),
    .io_wr(FIFO_A_3_1_hit_io_wr),
    .io_rd(FIFO_A_3_1_hit_io_rd),
    .io_empty(FIFO_A_3_1_hit_io_empty)
  );
  FIFO FIFO_A_3_2_node ( // @[Arbitration_3.scala 50:38]
    .clock(FIFO_A_3_2_node_clock),
    .reset(FIFO_A_3_2_node_reset),
    .io_datain(FIFO_A_3_2_node_io_datain),
    .io_dataout(FIFO_A_3_2_node_io_dataout),
    .io_wr(FIFO_A_3_2_node_io_wr),
    .io_rd(FIFO_A_3_2_node_io_rd),
    .io_empty(FIFO_A_3_2_node_io_empty)
  );
  FIFO_0 FIFO_A_3_2_ray ( // @[Arbitration_3.scala 51:41]
    .clock(FIFO_A_3_2_ray_clock),
    .reset(FIFO_A_3_2_ray_reset),
    .io_datain(FIFO_A_3_2_ray_io_datain),
    .io_dataout(FIFO_A_3_2_ray_io_dataout),
    .io_wr(FIFO_A_3_2_ray_io_wr),
    .io_rd(FIFO_A_3_2_ray_io_rd),
    .io_empty(FIFO_A_3_2_ray_io_empty)
  );
  FIFO_0 FIFO_A_3_2_hit ( // @[Arbitration_3.scala 52:42]
    .clock(FIFO_A_3_2_hit_clock),
    .reset(FIFO_A_3_2_hit_reset),
    .io_datain(FIFO_A_3_2_hit_io_datain),
    .io_dataout(FIFO_A_3_2_hit_io_dataout),
    .io_wr(FIFO_A_3_2_hit_io_wr),
    .io_rd(FIFO_A_3_2_hit_io_rd),
    .io_empty(FIFO_A_3_2_hit_io_empty)
  );
  FIFO FIFO_A_3_3_node ( // @[Arbitration_3.scala 54:38]
    .clock(FIFO_A_3_3_node_clock),
    .reset(FIFO_A_3_3_node_reset),
    .io_datain(FIFO_A_3_3_node_io_datain),
    .io_dataout(FIFO_A_3_3_node_io_dataout),
    .io_wr(FIFO_A_3_3_node_io_wr),
    .io_rd(FIFO_A_3_3_node_io_rd),
    .io_empty(FIFO_A_3_3_node_io_empty)
  );
  FIFO_0 FIFO_A_3_3_ray ( // @[Arbitration_3.scala 55:41]
    .clock(FIFO_A_3_3_ray_clock),
    .reset(FIFO_A_3_3_ray_reset),
    .io_datain(FIFO_A_3_3_ray_io_datain),
    .io_dataout(FIFO_A_3_3_ray_io_dataout),
    .io_wr(FIFO_A_3_3_ray_io_wr),
    .io_rd(FIFO_A_3_3_ray_io_rd),
    .io_empty(FIFO_A_3_3_ray_io_empty)
  );
  FIFO_0 FIFO_A_3_3_hit ( // @[Arbitration_3.scala 56:42]
    .clock(FIFO_A_3_3_hit_clock),
    .reset(FIFO_A_3_3_hit_reset),
    .io_datain(FIFO_A_3_3_hit_io_datain),
    .io_dataout(FIFO_A_3_3_hit_io_dataout),
    .io_wr(FIFO_A_3_3_hit_io_wr),
    .io_rd(FIFO_A_3_3_hit_io_rd),
    .io_empty(FIFO_A_3_3_hit_io_empty)
  );
  FIFO FIFO_A_3_4_node ( // @[Arbitration_3.scala 58:38]
    .clock(FIFO_A_3_4_node_clock),
    .reset(FIFO_A_3_4_node_reset),
    .io_datain(FIFO_A_3_4_node_io_datain),
    .io_dataout(FIFO_A_3_4_node_io_dataout),
    .io_wr(FIFO_A_3_4_node_io_wr),
    .io_rd(FIFO_A_3_4_node_io_rd),
    .io_empty(FIFO_A_3_4_node_io_empty)
  );
  FIFO_0 FIFO_A_3_4_ray ( // @[Arbitration_3.scala 59:41]
    .clock(FIFO_A_3_4_ray_clock),
    .reset(FIFO_A_3_4_ray_reset),
    .io_datain(FIFO_A_3_4_ray_io_datain),
    .io_dataout(FIFO_A_3_4_ray_io_dataout),
    .io_wr(FIFO_A_3_4_ray_io_wr),
    .io_rd(FIFO_A_3_4_ray_io_rd),
    .io_empty(FIFO_A_3_4_ray_io_empty)
  );
  FIFO_0 FIFO_A_3_4_hit ( // @[Arbitration_3.scala 60:42]
    .clock(FIFO_A_3_4_hit_clock),
    .reset(FIFO_A_3_4_hit_reset),
    .io_datain(FIFO_A_3_4_hit_io_datain),
    .io_dataout(FIFO_A_3_4_hit_io_dataout),
    .io_wr(FIFO_A_3_4_hit_io_wr),
    .io_rd(FIFO_A_3_4_hit_io_rd),
    .io_empty(FIFO_A_3_4_hit_io_empty)
  );
  assign io_node_id_out = ~FIFO_0_empty ? $signed(FIFO_A_3_0_node_io_dataout) : $signed(_GEN_31); // @[Arbitration_3.scala 227:35 Arbitration_3.scala 228:46]
  assign io_ray_id_out = ~FIFO_0_empty ? FIFO_A_3_0_ray_io_dataout : _GEN_32; // @[Arbitration_3.scala 227:35 Arbitration_3.scala 229:48]
  assign io_hit_out = ~FIFO_0_empty ? FIFO_A_3_0_hit_io_dataout : _GEN_33; // @[Arbitration_3.scala 227:35 Arbitration_3.scala 230:53]
  assign io_valid_out = ~FIFO_0_empty ? valid_out_temp : _GEN_34; // @[Arbitration_3.scala 227:35 Arbitration_3.scala 231:50]
  assign FIFO_A_3_0_node_clock = clock;
  assign FIFO_A_3_0_node_reset = reset;
  assign FIFO_A_3_0_node_io_datain = io_node_id_3_0; // @[Arbitration_3.scala 66:40]
  assign FIFO_A_3_0_node_io_wr = io_valid_3_0; // @[Arbitration_3.scala 63:44]
  assign FIFO_A_3_0_node_io_rd = ~FIFO_A_3_0_node_io_empty; // @[Arbitration_3.scala 103:39]
  assign FIFO_A_3_0_ray_clock = clock;
  assign FIFO_A_3_0_ray_reset = reset;
  assign FIFO_A_3_0_ray_io_datain = io_ray_id_3_0; // @[Arbitration_3.scala 67:43]
  assign FIFO_A_3_0_ray_io_wr = io_valid_3_0; // @[Arbitration_3.scala 64:47]
  assign FIFO_A_3_0_ray_io_rd = ~FIFO_A_3_0_node_io_empty; // @[Arbitration_3.scala 103:39]
  assign FIFO_A_3_0_hit_clock = clock;
  assign FIFO_A_3_0_hit_reset = reset;
  assign FIFO_A_3_0_hit_io_datain = io_hit_3_0; // @[Arbitration_3.scala 68:44]
  assign FIFO_A_3_0_hit_io_wr = io_valid_3_0; // @[Arbitration_3.scala 65:48]
  assign FIFO_A_3_0_hit_io_rd = ~FIFO_A_3_0_node_io_empty; // @[Arbitration_3.scala 103:39]
  assign FIFO_A_3_1_node_clock = clock;
  assign FIFO_A_3_1_node_reset = reset;
  assign FIFO_A_3_1_node_io_datain = io_node_id_3_1; // @[Arbitration_3.scala 73:40]
  assign FIFO_A_3_1_node_io_wr = io_valid_3_1; // @[Arbitration_3.scala 70:44]
  assign FIFO_A_3_1_node_io_rd = ~FIFO_A_3_0_node_io_empty ? 1'h0 : _T_3; // @[Arbitration_3.scala 103:47 Arbitration_3.scala 107:44]
  assign FIFO_A_3_1_ray_clock = clock;
  assign FIFO_A_3_1_ray_reset = reset;
  assign FIFO_A_3_1_ray_io_datain = io_ray_id_3_1; // @[Arbitration_3.scala 74:43]
  assign FIFO_A_3_1_ray_io_wr = io_valid_3_1; // @[Arbitration_3.scala 71:47]
  assign FIFO_A_3_1_ray_io_rd = ~FIFO_A_3_0_node_io_empty ? 1'h0 : _T_3; // @[Arbitration_3.scala 103:47 Arbitration_3.scala 107:44]
  assign FIFO_A_3_1_hit_clock = clock;
  assign FIFO_A_3_1_hit_reset = reset;
  assign FIFO_A_3_1_hit_io_datain = io_hit_3_1; // @[Arbitration_3.scala 75:44]
  assign FIFO_A_3_1_hit_io_wr = io_valid_3_1; // @[Arbitration_3.scala 72:48]
  assign FIFO_A_3_1_hit_io_rd = ~FIFO_A_3_0_node_io_empty ? 1'h0 : _T_3; // @[Arbitration_3.scala 103:47 Arbitration_3.scala 107:44]
  assign FIFO_A_3_2_node_clock = clock;
  assign FIFO_A_3_2_node_reset = reset;
  assign FIFO_A_3_2_node_io_datain = io_node_id_3_2; // @[Arbitration_3.scala 80:40]
  assign FIFO_A_3_2_node_io_wr = io_valid_3_2; // @[Arbitration_3.scala 77:44]
  assign FIFO_A_3_2_node_io_rd = ~FIFO_A_3_0_node_io_empty ? 1'h0 : _GEN_11; // @[Arbitration_3.scala 103:47 Arbitration_3.scala 110:44]
  assign FIFO_A_3_2_ray_clock = clock;
  assign FIFO_A_3_2_ray_reset = reset;
  assign FIFO_A_3_2_ray_io_datain = io_ray_id_3_2; // @[Arbitration_3.scala 81:43]
  assign FIFO_A_3_2_ray_io_wr = io_valid_3_2; // @[Arbitration_3.scala 78:47]
  assign FIFO_A_3_2_ray_io_rd = ~FIFO_A_3_0_node_io_empty ? 1'h0 : _GEN_11; // @[Arbitration_3.scala 103:47 Arbitration_3.scala 110:44]
  assign FIFO_A_3_2_hit_clock = clock;
  assign FIFO_A_3_2_hit_reset = reset;
  assign FIFO_A_3_2_hit_io_datain = io_hit_3_2; // @[Arbitration_3.scala 82:44]
  assign FIFO_A_3_2_hit_io_wr = io_valid_3_2; // @[Arbitration_3.scala 79:48]
  assign FIFO_A_3_2_hit_io_rd = ~FIFO_A_3_0_node_io_empty ? 1'h0 : _GEN_11; // @[Arbitration_3.scala 103:47 Arbitration_3.scala 110:44]
  assign FIFO_A_3_3_node_clock = clock;
  assign FIFO_A_3_3_node_reset = reset;
  assign FIFO_A_3_3_node_io_datain = io_node_id_3_3; // @[Arbitration_3.scala 87:40]
  assign FIFO_A_3_3_node_io_wr = io_valid_3_3; // @[Arbitration_3.scala 84:44]
  assign FIFO_A_3_3_node_io_rd = ~FIFO_A_3_0_node_io_empty ? 1'h0 : _GEN_12; // @[Arbitration_3.scala 103:47 Arbitration_3.scala 113:44]
  assign FIFO_A_3_3_ray_clock = clock;
  assign FIFO_A_3_3_ray_reset = reset;
  assign FIFO_A_3_3_ray_io_datain = io_ray_id_3_3; // @[Arbitration_3.scala 88:43]
  assign FIFO_A_3_3_ray_io_wr = io_valid_3_3; // @[Arbitration_3.scala 85:47]
  assign FIFO_A_3_3_ray_io_rd = ~FIFO_A_3_0_node_io_empty ? 1'h0 : _GEN_12; // @[Arbitration_3.scala 103:47 Arbitration_3.scala 113:44]
  assign FIFO_A_3_3_hit_clock = clock;
  assign FIFO_A_3_3_hit_reset = reset;
  assign FIFO_A_3_3_hit_io_datain = io_hit_3_3; // @[Arbitration_3.scala 89:44]
  assign FIFO_A_3_3_hit_io_wr = io_valid_3_3; // @[Arbitration_3.scala 86:48]
  assign FIFO_A_3_3_hit_io_rd = ~FIFO_A_3_0_node_io_empty ? 1'h0 : _GEN_12; // @[Arbitration_3.scala 103:47 Arbitration_3.scala 113:44]
  assign FIFO_A_3_4_node_clock = clock;
  assign FIFO_A_3_4_node_reset = reset;
  assign FIFO_A_3_4_node_io_datain = io_node_id_3_4; // @[Arbitration_3.scala 94:40]
  assign FIFO_A_3_4_node_io_wr = io_valid_3_4; // @[Arbitration_3.scala 91:44]
  assign FIFO_A_3_4_node_io_rd = ~FIFO_A_3_0_node_io_empty ? 1'h0 : _GEN_13; // @[Arbitration_3.scala 103:47 Arbitration_3.scala 116:44]
  assign FIFO_A_3_4_ray_clock = clock;
  assign FIFO_A_3_4_ray_reset = reset;
  assign FIFO_A_3_4_ray_io_datain = io_ray_id_3_4; // @[Arbitration_3.scala 95:43]
  assign FIFO_A_3_4_ray_io_wr = io_valid_3_4; // @[Arbitration_3.scala 92:47]
  assign FIFO_A_3_4_ray_io_rd = ~FIFO_A_3_0_node_io_empty ? 1'h0 : _GEN_13; // @[Arbitration_3.scala 103:47 Arbitration_3.scala 116:44]
  assign FIFO_A_3_4_hit_clock = clock;
  assign FIFO_A_3_4_hit_reset = reset;
  assign FIFO_A_3_4_hit_io_datain = io_hit_3_4; // @[Arbitration_3.scala 96:44]
  assign FIFO_A_3_4_hit_io_wr = io_valid_3_4; // @[Arbitration_3.scala 93:48]
  assign FIFO_A_3_4_hit_io_rd = ~FIFO_A_3_0_node_io_empty ? 1'h0 : _GEN_13; // @[Arbitration_3.scala 103:47 Arbitration_3.scala 116:44]
  always @(posedge clock) begin
    if (reset) begin // @[Arbitration_3.scala 101:59]
      valid_out_temp <= 1'h0; // @[Arbitration_3.scala 101:59]
    end else begin
      valid_out_temp <= FIFO_A_3_0_node_io_rd | FIFO_A_3_1_node_io_rd | FIFO_A_3_2_node_io_rd | FIFO_A_3_3_node_io_rd |
        FIFO_A_3_4_node_io_rd; // @[Arbitration_3.scala 225:51]
    end
    if (reset) begin // @[Arbitration_3.scala 200:58]
      FIFO_0_empty <= 1'h0; // @[Arbitration_3.scala 200:58]
    end else begin
      FIFO_0_empty <= FIFO_A_3_0_node_io_empty; // @[Arbitration_3.scala 206:52]
    end
    if (reset) begin // @[Arbitration_3.scala 201:58]
      FIFO_1_empty <= 1'h0; // @[Arbitration_3.scala 201:58]
    end else begin
      FIFO_1_empty <= FIFO_A_3_1_node_io_empty; // @[Arbitration_3.scala 207:52]
    end
    if (reset) begin // @[Arbitration_3.scala 202:58]
      FIFO_2_empty <= 1'h0; // @[Arbitration_3.scala 202:58]
    end else begin
      FIFO_2_empty <= FIFO_A_3_2_node_io_empty; // @[Arbitration_3.scala 208:52]
    end
    if (reset) begin // @[Arbitration_3.scala 203:58]
      FIFO_3_empty <= 1'h0; // @[Arbitration_3.scala 203:58]
    end else begin
      FIFO_3_empty <= FIFO_A_3_3_node_io_empty; // @[Arbitration_3.scala 209:52]
    end
    if (reset) begin // @[Arbitration_3.scala 204:58]
      FIFO_4_empty <= 1'h0; // @[Arbitration_3.scala 204:58]
    end else begin
      FIFO_4_empty <= FIFO_A_3_4_node_io_empty; // @[Arbitration_3.scala 210:52]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid_out_temp = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  FIFO_0_empty = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  FIFO_1_empty = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  FIFO_2_empty = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  FIFO_3_empty = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  FIFO_4_empty = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FSM_1(
  input   clock,
  input   reset,
  input   io_request_0,
  input   io_request_1,
  output  io_grant_0,
  output  io_grant_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] grant; // @[FSM.scala 18:26]
  reg [1:0] stateReg; // @[FSM.scala 19:23]
  wire  _T = 2'h0 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_4 = ~io_request_1; // @[FSM.scala 29:44]
  wire [1:0] _GEN_2 = ~io_request_0 & io_request_1 ? 2'h2 : 2'h0; // @[FSM.scala 26:56 FSM.scala 27:27]
  wire [1:0] _GEN_4 = io_request_0 ? 2'h1 : _GEN_2; // @[FSM.scala 23:31 FSM.scala 24:27]
  wire  _T_6 = 2'h1 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_8 = _T_4 & io_request_0; // @[FSM.scala 41:39]
  wire  _T_12 = 2'h2 == stateReg; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_16 = io_request_0 ? 2'h1 : 2'h2; // @[FSM.scala 53:31 FSM.scala 54:27]
  assign io_grant_0 = grant == 2'h1; // @[FSM.scala 90:38]
  assign io_grant_1 = grant == 2'h2; // @[FSM.scala 91:38]
  always @(posedge clock) begin
    if (reset) begin // @[FSM.scala 18:26]
      grant <= 2'h0; // @[FSM.scala 18:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      grant <= _GEN_4;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      if (io_request_1) begin // @[FSM.scala 38:31]
        grant <= 2'h2; // @[FSM.scala 40:31]
      end else begin
        grant <= {{1'd0}, _T_8};
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      grant <= _GEN_4;
    end
    if (reset) begin // @[FSM.scala 19:23]
      stateReg <= 2'h0; // @[FSM.scala 19:23]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_request_0) begin // @[FSM.scala 23:31]
        stateReg <= 2'h1; // @[FSM.scala 24:27]
      end else if (~io_request_0 & io_request_1) begin // @[FSM.scala 26:56]
        stateReg <= 2'h2; // @[FSM.scala 27:27]
      end else begin
        stateReg <= 2'h0;
      end
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      if (io_request_1) begin // @[FSM.scala 38:31]
        stateReg <= 2'h2; // @[FSM.scala 39:27]
      end else begin
        stateReg <= 2'h1;
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      stateReg <= _GEN_16;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  grant = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  stateReg = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbitration_4(
  input         clock,
  input         reset,
  input  [31:0] io_node_id_4_0,
  input  [31:0] io_ray_id_4_0,
  input  [31:0] io_hit_4_0,
  input         io_valid_4_0,
  input  [31:0] io_node_id_4_1,
  input  [31:0] io_ray_id_4_1,
  input  [31:0] io_hit_4_1,
  input         io_valid_4_1,
  output [31:0] io_node_id_out,
  output [31:0] io_ray_id_out,
  output [31:0] io_hit_out,
  output        io_RAY_AABB_out,
  output        io_RAY_AABB_2_out,
  output        io_valid_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  FSM_clock; // @[Arbitration_4.scala 31:55]
  wire  FSM_reset; // @[Arbitration_4.scala 31:55]
  wire  FSM_io_request_0; // @[Arbitration_4.scala 31:55]
  wire  FSM_io_request_1; // @[Arbitration_4.scala 31:55]
  wire  FSM_io_grant_0; // @[Arbitration_4.scala 31:55]
  wire  FSM_io_grant_1; // @[Arbitration_4.scala 31:55]
  wire  FIFO_A_4_0_node_clock; // @[Arbitration_4.scala 33:38]
  wire  FIFO_A_4_0_node_reset; // @[Arbitration_4.scala 33:38]
  wire [31:0] FIFO_A_4_0_node_io_datain; // @[Arbitration_4.scala 33:38]
  wire [31:0] FIFO_A_4_0_node_io_dataout; // @[Arbitration_4.scala 33:38]
  wire  FIFO_A_4_0_node_io_wr; // @[Arbitration_4.scala 33:38]
  wire  FIFO_A_4_0_node_io_rd; // @[Arbitration_4.scala 33:38]
  wire  FIFO_A_4_0_node_io_empty; // @[Arbitration_4.scala 33:38]
  wire  FIFO_A_4_0_ray_clock; // @[Arbitration_4.scala 34:41]
  wire  FIFO_A_4_0_ray_reset; // @[Arbitration_4.scala 34:41]
  wire [31:0] FIFO_A_4_0_ray_io_datain; // @[Arbitration_4.scala 34:41]
  wire [31:0] FIFO_A_4_0_ray_io_dataout; // @[Arbitration_4.scala 34:41]
  wire  FIFO_A_4_0_ray_io_wr; // @[Arbitration_4.scala 34:41]
  wire  FIFO_A_4_0_ray_io_rd; // @[Arbitration_4.scala 34:41]
  wire  FIFO_A_4_0_ray_io_empty; // @[Arbitration_4.scala 34:41]
  wire  FIFO_A_4_0_hit_clock; // @[Arbitration_4.scala 35:42]
  wire  FIFO_A_4_0_hit_reset; // @[Arbitration_4.scala 35:42]
  wire [31:0] FIFO_A_4_0_hit_io_datain; // @[Arbitration_4.scala 35:42]
  wire [31:0] FIFO_A_4_0_hit_io_dataout; // @[Arbitration_4.scala 35:42]
  wire  FIFO_A_4_0_hit_io_wr; // @[Arbitration_4.scala 35:42]
  wire  FIFO_A_4_0_hit_io_rd; // @[Arbitration_4.scala 35:42]
  wire  FIFO_A_4_0_hit_io_empty; // @[Arbitration_4.scala 35:42]
  wire  FIFO_A_4_1_node_clock; // @[Arbitration_4.scala 37:38]
  wire  FIFO_A_4_1_node_reset; // @[Arbitration_4.scala 37:38]
  wire [31:0] FIFO_A_4_1_node_io_datain; // @[Arbitration_4.scala 37:38]
  wire [31:0] FIFO_A_4_1_node_io_dataout; // @[Arbitration_4.scala 37:38]
  wire  FIFO_A_4_1_node_io_wr; // @[Arbitration_4.scala 37:38]
  wire  FIFO_A_4_1_node_io_rd; // @[Arbitration_4.scala 37:38]
  wire  FIFO_A_4_1_node_io_empty; // @[Arbitration_4.scala 37:38]
  wire  FIFO_A_4_1_ray_clock; // @[Arbitration_4.scala 38:41]
  wire  FIFO_A_4_1_ray_reset; // @[Arbitration_4.scala 38:41]
  wire [31:0] FIFO_A_4_1_ray_io_datain; // @[Arbitration_4.scala 38:41]
  wire [31:0] FIFO_A_4_1_ray_io_dataout; // @[Arbitration_4.scala 38:41]
  wire  FIFO_A_4_1_ray_io_wr; // @[Arbitration_4.scala 38:41]
  wire  FIFO_A_4_1_ray_io_rd; // @[Arbitration_4.scala 38:41]
  wire  FIFO_A_4_1_ray_io_empty; // @[Arbitration_4.scala 38:41]
  wire  FIFO_A_4_1_hit_clock; // @[Arbitration_4.scala 39:42]
  wire  FIFO_A_4_1_hit_reset; // @[Arbitration_4.scala 39:42]
  wire [31:0] FIFO_A_4_1_hit_io_datain; // @[Arbitration_4.scala 39:42]
  wire [31:0] FIFO_A_4_1_hit_io_dataout; // @[Arbitration_4.scala 39:42]
  wire  FIFO_A_4_1_hit_io_wr; // @[Arbitration_4.scala 39:42]
  wire  FIFO_A_4_1_hit_io_rd; // @[Arbitration_4.scala 39:42]
  wire  FIFO_A_4_1_hit_io_empty; // @[Arbitration_4.scala 39:42]
  wire  _T = ~FIFO_A_4_0_ray_io_empty; // @[Arbitration_4.scala 59:76]
  wire  _T_1 = ~FIFO_A_4_1_ray_io_empty; // @[Arbitration_4.scala 60:76]
  reg  valid_0; // @[Arbitration_4.scala 61:66]
  reg  valid_1; // @[Arbitration_4.scala 62:66]
  wire  _T_3 = FSM_io_grant_0 & _T; // @[Arbitration_4.scala 63:28]
  wire  _T_5 = FSM_io_grant_1 & _T_1; // @[Arbitration_4.scala 72:35]
  wire [31:0] _GEN_4 = valid_1 ? $signed(FIFO_A_4_1_node_io_dataout) : $signed(32'sh0); // @[Arbitration_4.scala 134:34 Arbitration_4.scala 135:45 Arbitration_4.scala 151:46]
  wire [31:0] _GEN_5 = valid_1 ? FIFO_A_4_1_ray_io_dataout : 32'h0; // @[Arbitration_4.scala 134:34 Arbitration_4.scala 136:48 Arbitration_4.scala 152:48]
  wire [31:0] _GEN_6 = valid_1 ? FIFO_A_4_1_hit_io_dataout : 32'h0; // @[Arbitration_4.scala 134:34 Arbitration_4.scala 137:53 Arbitration_4.scala 153:53]
  FSM_1 FSM ( // @[Arbitration_4.scala 31:55]
    .clock(FSM_clock),
    .reset(FSM_reset),
    .io_request_0(FSM_io_request_0),
    .io_request_1(FSM_io_request_1),
    .io_grant_0(FSM_io_grant_0),
    .io_grant_1(FSM_io_grant_1)
  );
  FIFO FIFO_A_4_0_node ( // @[Arbitration_4.scala 33:38]
    .clock(FIFO_A_4_0_node_clock),
    .reset(FIFO_A_4_0_node_reset),
    .io_datain(FIFO_A_4_0_node_io_datain),
    .io_dataout(FIFO_A_4_0_node_io_dataout),
    .io_wr(FIFO_A_4_0_node_io_wr),
    .io_rd(FIFO_A_4_0_node_io_rd),
    .io_empty(FIFO_A_4_0_node_io_empty)
  );
  FIFO_0 FIFO_A_4_0_ray ( // @[Arbitration_4.scala 34:41]
    .clock(FIFO_A_4_0_ray_clock),
    .reset(FIFO_A_4_0_ray_reset),
    .io_datain(FIFO_A_4_0_ray_io_datain),
    .io_dataout(FIFO_A_4_0_ray_io_dataout),
    .io_wr(FIFO_A_4_0_ray_io_wr),
    .io_rd(FIFO_A_4_0_ray_io_rd),
    .io_empty(FIFO_A_4_0_ray_io_empty)
  );
  FIFO_0 FIFO_A_4_0_hit ( // @[Arbitration_4.scala 35:42]
    .clock(FIFO_A_4_0_hit_clock),
    .reset(FIFO_A_4_0_hit_reset),
    .io_datain(FIFO_A_4_0_hit_io_datain),
    .io_dataout(FIFO_A_4_0_hit_io_dataout),
    .io_wr(FIFO_A_4_0_hit_io_wr),
    .io_rd(FIFO_A_4_0_hit_io_rd),
    .io_empty(FIFO_A_4_0_hit_io_empty)
  );
  FIFO FIFO_A_4_1_node ( // @[Arbitration_4.scala 37:38]
    .clock(FIFO_A_4_1_node_clock),
    .reset(FIFO_A_4_1_node_reset),
    .io_datain(FIFO_A_4_1_node_io_datain),
    .io_dataout(FIFO_A_4_1_node_io_dataout),
    .io_wr(FIFO_A_4_1_node_io_wr),
    .io_rd(FIFO_A_4_1_node_io_rd),
    .io_empty(FIFO_A_4_1_node_io_empty)
  );
  FIFO_0 FIFO_A_4_1_ray ( // @[Arbitration_4.scala 38:41]
    .clock(FIFO_A_4_1_ray_clock),
    .reset(FIFO_A_4_1_ray_reset),
    .io_datain(FIFO_A_4_1_ray_io_datain),
    .io_dataout(FIFO_A_4_1_ray_io_dataout),
    .io_wr(FIFO_A_4_1_ray_io_wr),
    .io_rd(FIFO_A_4_1_ray_io_rd),
    .io_empty(FIFO_A_4_1_ray_io_empty)
  );
  FIFO_0 FIFO_A_4_1_hit ( // @[Arbitration_4.scala 39:42]
    .clock(FIFO_A_4_1_hit_clock),
    .reset(FIFO_A_4_1_hit_reset),
    .io_datain(FIFO_A_4_1_hit_io_datain),
    .io_dataout(FIFO_A_4_1_hit_io_dataout),
    .io_wr(FIFO_A_4_1_hit_io_wr),
    .io_rd(FIFO_A_4_1_hit_io_rd),
    .io_empty(FIFO_A_4_1_hit_io_empty)
  );
  assign io_node_id_out = valid_0 ? $signed(FIFO_A_4_0_node_io_dataout) : $signed(_GEN_4); // @[Arbitration_4.scala 126:29 Arbitration_4.scala 127:46]
  assign io_ray_id_out = valid_0 ? FIFO_A_4_0_ray_io_dataout : _GEN_5; // @[Arbitration_4.scala 126:29 Arbitration_4.scala 128:48]
  assign io_hit_out = valid_0 ? FIFO_A_4_0_hit_io_dataout : _GEN_6; // @[Arbitration_4.scala 126:29 Arbitration_4.scala 129:53]
  assign io_RAY_AABB_out = valid_0; // @[Arbitration_4.scala 126:29 Arbitration_4.scala 131:41]
  assign io_RAY_AABB_2_out = valid_0 ? 1'h0 : valid_1; // @[Arbitration_4.scala 126:29 Arbitration_4.scala 132:38]
  assign io_valid_out = valid_0 | valid_1; // @[Arbitration_4.scala 126:29 Arbitration_4.scala 130:50]
  assign FSM_clock = clock;
  assign FSM_reset = reset;
  assign FSM_io_request_0 = ~FIFO_A_4_0_ray_io_empty; // @[Arbitration_4.scala 59:76]
  assign FSM_io_request_1 = ~FIFO_A_4_1_ray_io_empty; // @[Arbitration_4.scala 60:76]
  assign FIFO_A_4_0_node_clock = clock;
  assign FIFO_A_4_0_node_reset = reset;
  assign FIFO_A_4_0_node_io_datain = io_node_id_4_0; // @[Arbitration_4.scala 44:40]
  assign FIFO_A_4_0_node_io_wr = io_valid_4_0; // @[Arbitration_4.scala 41:44]
  assign FIFO_A_4_0_node_io_rd = FSM_io_grant_0 & _T; // @[Arbitration_4.scala 63:28]
  assign FIFO_A_4_0_ray_clock = clock;
  assign FIFO_A_4_0_ray_reset = reset;
  assign FIFO_A_4_0_ray_io_datain = io_ray_id_4_0; // @[Arbitration_4.scala 45:43]
  assign FIFO_A_4_0_ray_io_wr = io_valid_4_0; // @[Arbitration_4.scala 42:47]
  assign FIFO_A_4_0_ray_io_rd = FSM_io_grant_0 & _T; // @[Arbitration_4.scala 63:28]
  assign FIFO_A_4_0_hit_clock = clock;
  assign FIFO_A_4_0_hit_reset = reset;
  assign FIFO_A_4_0_hit_io_datain = io_hit_4_0; // @[Arbitration_4.scala 46:44]
  assign FIFO_A_4_0_hit_io_wr = io_valid_4_0; // @[Arbitration_4.scala 43:48]
  assign FIFO_A_4_0_hit_io_rd = FSM_io_grant_0 & _T; // @[Arbitration_4.scala 63:28]
  assign FIFO_A_4_1_node_clock = clock;
  assign FIFO_A_4_1_node_reset = reset;
  assign FIFO_A_4_1_node_io_datain = io_node_id_4_1; // @[Arbitration_4.scala 51:40]
  assign FIFO_A_4_1_node_io_wr = io_valid_4_1; // @[Arbitration_4.scala 48:44]
  assign FIFO_A_4_1_node_io_rd = FSM_io_grant_0 & _T ? 1'h0 : _T_5; // @[Arbitration_4.scala 63:57 Arbitration_4.scala 67:44]
  assign FIFO_A_4_1_ray_clock = clock;
  assign FIFO_A_4_1_ray_reset = reset;
  assign FIFO_A_4_1_ray_io_datain = io_ray_id_4_1; // @[Arbitration_4.scala 52:43]
  assign FIFO_A_4_1_ray_io_wr = io_valid_4_1; // @[Arbitration_4.scala 49:47]
  assign FIFO_A_4_1_ray_io_rd = FSM_io_grant_0 & _T ? 1'h0 : _T_5; // @[Arbitration_4.scala 63:57 Arbitration_4.scala 67:44]
  assign FIFO_A_4_1_hit_clock = clock;
  assign FIFO_A_4_1_hit_reset = reset;
  assign FIFO_A_4_1_hit_io_datain = io_hit_4_1; // @[Arbitration_4.scala 53:44]
  assign FIFO_A_4_1_hit_io_wr = io_valid_4_1; // @[Arbitration_4.scala 50:48]
  assign FIFO_A_4_1_hit_io_rd = FSM_io_grant_0 & _T ? 1'h0 : _T_5; // @[Arbitration_4.scala 63:57 Arbitration_4.scala 67:44]
  always @(posedge clock) begin
    if (reset) begin // @[Arbitration_4.scala 61:66]
      valid_0 <= 1'h0; // @[Arbitration_4.scala 61:66]
    end else begin
      valid_0 <= _T_3;
    end
    if (reset) begin // @[Arbitration_4.scala 62:66]
      valid_1 <= 1'h0; // @[Arbitration_4.scala 62:66]
    end else if (FSM_io_grant_0 & _T) begin // @[Arbitration_4.scala 63:57]
      valid_1 <= 1'h0; // @[Arbitration_4.scala 67:44]
    end else begin
      valid_1 <= _T_5;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  valid_1 = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LUT(
  input         clock,
  input         reset,
  input         io_push,
  input         io_push_valid,
  input         io_pop,
  input         io_pop_valid,
  input         io_clear,
  input         io_empty_0,
  input         io_empty_1,
  input         io_empty_2,
  input         io_empty_3,
  input         io_empty_4,
  input         io_empty_5,
  input         io_empty_6,
  input         io_empty_7,
  input         io_empty_8,
  input         io_empty_9,
  input         io_empty_10,
  input         io_empty_11,
  input         io_empty_12,
  input         io_empty_13,
  input         io_empty_14,
  input         io_empty_15,
  input         io_empty_16,
  input         io_empty_17,
  input         io_empty_18,
  input         io_empty_19,
  input         io_empty_20,
  input         io_empty_21,
  input         io_empty_22,
  input         io_empty_23,
  input         io_empty_24,
  input         io_empty_25,
  input         io_empty_26,
  input         io_empty_27,
  input         io_empty_28,
  input         io_empty_29,
  input         io_empty_30,
  input         io_empty_31,
  input         io_empty_32,
  input         io_empty_33,
  input         io_empty_34,
  input         io_dispatch_0,
  input         io_dispatch_1,
  input         io_dispatch_2,
  input         io_dispatch_3,
  input         io_dispatch_4,
  input         io_dispatch_5,
  input         io_dispatch_6,
  input         io_dispatch_7,
  input         io_dispatch_8,
  input         io_dispatch_9,
  input         io_dispatch_10,
  input         io_dispatch_11,
  input         io_dispatch_12,
  input         io_dispatch_13,
  input         io_dispatch_14,
  input         io_dispatch_15,
  input         io_dispatch_16,
  input         io_dispatch_17,
  input         io_dispatch_18,
  input         io_dispatch_19,
  input         io_dispatch_20,
  input         io_dispatch_21,
  input         io_dispatch_22,
  input         io_dispatch_23,
  input         io_dispatch_24,
  input         io_dispatch_25,
  input         io_dispatch_26,
  input         io_dispatch_27,
  input         io_dispatch_28,
  input         io_dispatch_29,
  input         io_dispatch_30,
  input         io_dispatch_31,
  input         io_dispatch_32,
  input         io_dispatch_33,
  input         io_dispatch_34,
  input  [31:0] io_ray_id_push,
  input  [31:0] io_ray_id_pop,
  input  [31:0] io_node_id_push_in,
  input  [31:0] io_hitT_in,
  output [31:0] io_ray_id_pop_out,
  output [31:0] io_hitT_out,
  output        io_pop_0,
  output        io_pop_1,
  output        io_pop_2,
  output        io_pop_3,
  output        io_pop_4,
  output        io_pop_5,
  output        io_pop_6,
  output        io_pop_7,
  output        io_pop_8,
  output        io_pop_9,
  output        io_pop_10,
  output        io_pop_11,
  output        io_pop_12,
  output        io_pop_13,
  output        io_pop_14,
  output        io_pop_15,
  output        io_pop_16,
  output        io_pop_17,
  output        io_pop_18,
  output        io_pop_19,
  output        io_pop_20,
  output        io_pop_21,
  output        io_pop_22,
  output        io_pop_23,
  output        io_pop_24,
  output        io_pop_25,
  output        io_pop_26,
  output        io_pop_27,
  output        io_pop_28,
  output        io_pop_29,
  output        io_pop_30,
  output        io_pop_31,
  output        io_pop_32,
  output        io_pop_33,
  output        io_pop_34,
  output        io_pop_en,
  output        io_push_0,
  output        io_push_1,
  output        io_push_2,
  output        io_push_3,
  output        io_push_4,
  output        io_push_5,
  output        io_push_6,
  output        io_push_7,
  output        io_push_8,
  output        io_push_9,
  output        io_push_10,
  output        io_push_11,
  output        io_push_12,
  output        io_push_13,
  output        io_push_14,
  output        io_push_15,
  output        io_push_16,
  output        io_push_17,
  output        io_push_18,
  output        io_push_19,
  output        io_push_20,
  output        io_push_21,
  output        io_push_22,
  output        io_push_23,
  output        io_push_24,
  output        io_push_25,
  output        io_push_26,
  output        io_push_27,
  output        io_push_28,
  output        io_push_29,
  output        io_push_30,
  output        io_push_31,
  output        io_push_32,
  output        io_push_33,
  output        io_push_34,
  output        io_clear_0,
  output        io_clear_1,
  output        io_clear_2,
  output        io_clear_3,
  output        io_clear_4,
  output        io_clear_5,
  output        io_clear_6,
  output        io_clear_7,
  output        io_clear_8,
  output        io_clear_9,
  output        io_clear_10,
  output        io_clear_11,
  output        io_clear_12,
  output        io_clear_13,
  output        io_clear_14,
  output        io_clear_15,
  output        io_clear_16,
  output        io_clear_17,
  output        io_clear_18,
  output        io_clear_19,
  output        io_clear_20,
  output        io_clear_21,
  output        io_clear_22,
  output        io_clear_23,
  output        io_clear_24,
  output        io_clear_25,
  output        io_clear_26,
  output        io_clear_27,
  output        io_clear_28,
  output        io_clear_29,
  output        io_clear_30,
  output        io_clear_31,
  output        io_clear_32,
  output        io_clear_33,
  output        io_clear_34,
  output        io_push_en,
  output        io_no_match
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [63:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [63:0] _RAND_62;
  reg [63:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [63:0] _RAND_65;
  reg [63:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [63:0] _RAND_68;
  reg [63:0] _RAND_69;
  reg [63:0] _RAND_70;
  reg [63:0] _RAND_71;
  reg [63:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [63:0] _RAND_74;
  reg [63:0] _RAND_75;
  reg [63:0] _RAND_76;
  reg [63:0] _RAND_77;
  reg [63:0] _RAND_78;
  reg [63:0] _RAND_79;
  reg [63:0] _RAND_80;
  reg [63:0] _RAND_81;
  reg [63:0] _RAND_82;
  reg [63:0] _RAND_83;
  reg [63:0] _RAND_84;
  reg [63:0] _RAND_85;
  reg [63:0] _RAND_86;
  reg [63:0] _RAND_87;
  reg [63:0] _RAND_88;
  reg [63:0] _RAND_89;
  reg [63:0] _RAND_90;
  reg [63:0] _RAND_91;
  reg [63:0] _RAND_92;
  reg [63:0] _RAND_93;
  reg [63:0] _RAND_94;
  reg [63:0] _RAND_95;
  reg [63:0] _RAND_96;
  reg [63:0] _RAND_97;
  reg [63:0] _RAND_98;
  reg [63:0] _RAND_99;
  reg [63:0] _RAND_100;
  reg [63:0] _RAND_101;
  reg [63:0] _RAND_102;
  reg [63:0] _RAND_103;
  reg [63:0] _RAND_104;
  reg [63:0] _RAND_105;
  reg [63:0] _RAND_106;
  reg [63:0] _RAND_107;
  reg [63:0] _RAND_108;
  reg [63:0] _RAND_109;
  reg [63:0] _RAND_110;
  reg [63:0] _RAND_111;
  reg [63:0] _RAND_112;
  reg [63:0] _RAND_113;
  reg [63:0] _RAND_114;
  reg [63:0] _RAND_115;
  reg [63:0] _RAND_116;
  reg [63:0] _RAND_117;
  reg [63:0] _RAND_118;
  reg [63:0] _RAND_119;
  reg [63:0] _RAND_120;
  reg [63:0] _RAND_121;
  reg [63:0] _RAND_122;
  reg [63:0] _RAND_123;
  reg [63:0] _RAND_124;
  reg [63:0] _RAND_125;
  reg [63:0] _RAND_126;
  reg [63:0] _RAND_127;
  reg [63:0] _RAND_128;
  reg [63:0] _RAND_129;
  reg [63:0] _RAND_130;
  reg [63:0] _RAND_131;
  reg [63:0] _RAND_132;
  reg [63:0] _RAND_133;
  reg [63:0] _RAND_134;
  reg [63:0] _RAND_135;
  reg [63:0] _RAND_136;
  reg [63:0] _RAND_137;
  reg [63:0] _RAND_138;
  reg [63:0] _RAND_139;
  reg [63:0] _RAND_140;
  reg [63:0] _RAND_141;
  reg [63:0] _RAND_142;
  reg [63:0] _RAND_143;
  reg [63:0] _RAND_144;
  reg [63:0] _RAND_145;
  reg [63:0] _RAND_146;
  reg [63:0] _RAND_147;
  reg [63:0] _RAND_148;
  reg [63:0] _RAND_149;
  reg [63:0] _RAND_150;
  reg [63:0] _RAND_151;
  reg [63:0] _RAND_152;
  reg [63:0] _RAND_153;
  reg [63:0] _RAND_154;
  reg [63:0] _RAND_155;
  reg [63:0] _RAND_156;
  reg [63:0] _RAND_157;
  reg [63:0] _RAND_158;
  reg [63:0] _RAND_159;
  reg [63:0] _RAND_160;
  reg [63:0] _RAND_161;
  reg [63:0] _RAND_162;
  reg [63:0] _RAND_163;
  reg [63:0] _RAND_164;
  reg [63:0] _RAND_165;
  reg [63:0] _RAND_166;
  reg [63:0] _RAND_167;
  reg [63:0] _RAND_168;
  reg [63:0] _RAND_169;
  reg [63:0] _RAND_170;
  reg [63:0] _RAND_171;
  reg [63:0] _RAND_172;
  reg [63:0] _RAND_173;
  reg [63:0] _RAND_174;
  reg [63:0] _RAND_175;
  reg [63:0] _RAND_176;
  reg [63:0] _RAND_177;
  reg [63:0] _RAND_178;
  reg [63:0] _RAND_179;
  reg [63:0] _RAND_180;
  reg [63:0] _RAND_181;
  reg [63:0] _RAND_182;
  reg [63:0] _RAND_183;
  reg [63:0] _RAND_184;
  reg [63:0] _RAND_185;
  reg [63:0] _RAND_186;
  reg [63:0] _RAND_187;
  reg [63:0] _RAND_188;
  reg [63:0] _RAND_189;
  reg [63:0] _RAND_190;
  reg [63:0] _RAND_191;
  reg [63:0] _RAND_192;
  reg [63:0] _RAND_193;
  reg [63:0] _RAND_194;
  reg [63:0] _RAND_195;
  reg [63:0] _RAND_196;
  reg [63:0] _RAND_197;
  reg [63:0] _RAND_198;
  reg [63:0] _RAND_199;
  reg [63:0] _RAND_200;
  reg [63:0] _RAND_201;
  reg [63:0] _RAND_202;
  reg [63:0] _RAND_203;
  reg [63:0] _RAND_204;
  reg [63:0] _RAND_205;
  reg [63:0] _RAND_206;
  reg [63:0] _RAND_207;
  reg [63:0] _RAND_208;
  reg [63:0] _RAND_209;
  reg [63:0] _RAND_210;
  reg [63:0] _RAND_211;
  reg [63:0] _RAND_212;
  reg [63:0] _RAND_213;
  reg [63:0] _RAND_214;
  reg [63:0] _RAND_215;
  reg [63:0] _RAND_216;
  reg [63:0] _RAND_217;
  reg [63:0] _RAND_218;
  reg [63:0] _RAND_219;
  reg [63:0] _RAND_220;
  reg [63:0] _RAND_221;
  reg [63:0] _RAND_222;
  reg [63:0] _RAND_223;
  reg [63:0] _RAND_224;
  reg [63:0] _RAND_225;
  reg [63:0] _RAND_226;
  reg [63:0] _RAND_227;
  reg [63:0] _RAND_228;
  reg [63:0] _RAND_229;
  reg [63:0] _RAND_230;
  reg [63:0] _RAND_231;
  reg [63:0] _RAND_232;
  reg [63:0] _RAND_233;
  reg [63:0] _RAND_234;
  reg [63:0] _RAND_235;
  reg [63:0] _RAND_236;
  reg [63:0] _RAND_237;
  reg [63:0] _RAND_238;
  reg [63:0] _RAND_239;
  reg [63:0] _RAND_240;
  reg [63:0] _RAND_241;
  reg [63:0] _RAND_242;
  reg [63:0] _RAND_243;
  reg [63:0] _RAND_244;
  reg [63:0] _RAND_245;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
`endif // RANDOMIZE_REG_INIT
  reg [32:0] LUT_mem [0:34]; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_1_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_1_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_2_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_2_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_3_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_3_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_4_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_4_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_5_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_5_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_6_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_6_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_7_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_7_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_8_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_8_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_9_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_9_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_10_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_10_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_11_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_11_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_12_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_12_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_13_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_13_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_14_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_14_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_15_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_15_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_16_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_16_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_17_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_17_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_18_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_18_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_19_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_19_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_20_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_20_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_21_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_21_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_22_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_22_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_23_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_23_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_24_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_24_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_25_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_25_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_26_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_26_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_27_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_27_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_28_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_28_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_29_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_29_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_30_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_30_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_31_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_31_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_32_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_32_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_33_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_33_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_34_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_34_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_35_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_35_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_36_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_36_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_37_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_37_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_38_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_38_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_39_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_39_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_40_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_40_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_41_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_41_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_42_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_42_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_43_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_43_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_44_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_44_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_45_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_45_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_46_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_46_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_47_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_47_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_48_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_48_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_49_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_49_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_50_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_50_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_51_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_51_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_52_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_52_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_53_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_53_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_54_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_54_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_55_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_55_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_56_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_56_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_57_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_57_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_58_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_58_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_59_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_59_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_60_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_60_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_61_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_61_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_62_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_62_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_63_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_63_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_64_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_64_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_65_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_65_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_66_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_66_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_67_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_67_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_68_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_68_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_69_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_69_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_70_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_70_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_71_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_71_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_72_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_72_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_73_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_73_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_74_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_74_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_75_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_75_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_76_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_76_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_77_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_77_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_78_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_78_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_79_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_79_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_80_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_80_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_81_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_81_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_82_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_82_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_83_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_83_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_84_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_84_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_85_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_85_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_86_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_86_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_87_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_87_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_88_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_88_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_89_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_89_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_90_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_90_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_91_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_91_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_92_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_92_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_93_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_93_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_94_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_94_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_95_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_95_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_96_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_96_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_97_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_97_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_98_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_98_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_99_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_99_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_100_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_100_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_101_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_101_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_102_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_102_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_103_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_103_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_104_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_104_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_105_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_105_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_106_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_106_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_107_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_107_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_108_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_108_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_109_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_109_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_110_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_110_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_111_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_111_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_112_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_112_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_113_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_113_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_114_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_114_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_115_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_115_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_116_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_116_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_117_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_117_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_118_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_118_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_119_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_119_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_120_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_120_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_121_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_121_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_122_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_122_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_123_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_123_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_124_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_124_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_125_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_125_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_126_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_126_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_127_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_127_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_128_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_128_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_129_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_129_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_130_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_130_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_131_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_131_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_132_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_132_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_133_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_133_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_134_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_134_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_135_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_135_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_136_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_136_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_137_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_137_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_138_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_138_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_139_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_139_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_140_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_140_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_141_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_141_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_142_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_142_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_143_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_143_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_144_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_144_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_145_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_145_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_146_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_146_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_147_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_147_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_148_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_148_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_149_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_149_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_150_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_150_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_151_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_151_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_152_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_152_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_153_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_153_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_154_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_154_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_155_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_155_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_156_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_156_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_157_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_157_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_158_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_158_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_159_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_159_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_160_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_160_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_161_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_161_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_162_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_162_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_163_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_163_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_164_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_164_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_165_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_165_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_166_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_166_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_167_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_167_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_168_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_168_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_169_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_169_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_170_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_170_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_171_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_171_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_172_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_172_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_173_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_173_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_174_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_174_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_176_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_176_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_179_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_179_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_181_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_181_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_184_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_184_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_186_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_186_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_189_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_189_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_191_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_191_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_194_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_194_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_196_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_196_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_199_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_199_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_201_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_201_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_204_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_204_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_206_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_206_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_209_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_209_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_211_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_211_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_214_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_214_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_216_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_216_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_219_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_219_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_221_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_221_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_224_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_224_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_226_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_226_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_229_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_229_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_231_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_231_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_234_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_234_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_236_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_236_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_239_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_239_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_241_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_241_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_244_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_244_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_246_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_246_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_249_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_249_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_251_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_251_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_254_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_254_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_256_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_256_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_259_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_259_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_261_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_261_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_264_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_264_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_266_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_266_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_269_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_269_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_271_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_271_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_274_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_274_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_276_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_276_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_279_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_279_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_281_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_281_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_284_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_284_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_286_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_286_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_289_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_289_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_291_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_291_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_294_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_294_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_296_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_296_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_299_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_299_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_301_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_301_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_304_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_304_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_306_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_306_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_309_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_309_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_311_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_311_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_314_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_314_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_316_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_316_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_319_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_319_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_321_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_321_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_324_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_324_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_326_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_326_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_329_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_329_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_331_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_331_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_334_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_334_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_336_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_336_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_339_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_339_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_341_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_341_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_344_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_344_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_346_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_346_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_349_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_349_addr; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_175_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_175_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_175_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_175_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_177_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_177_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_177_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_177_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_178_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_178_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_178_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_178_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_180_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_180_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_180_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_180_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_182_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_182_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_182_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_182_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_183_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_183_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_183_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_183_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_185_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_185_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_185_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_185_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_187_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_187_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_187_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_187_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_188_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_188_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_188_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_188_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_190_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_190_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_190_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_190_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_192_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_192_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_192_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_192_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_193_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_193_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_193_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_193_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_195_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_195_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_195_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_195_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_197_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_197_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_197_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_197_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_198_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_198_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_198_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_198_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_200_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_200_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_200_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_200_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_202_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_202_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_202_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_202_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_203_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_203_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_203_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_203_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_205_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_205_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_205_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_205_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_207_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_207_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_207_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_207_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_208_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_208_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_208_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_208_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_210_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_210_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_210_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_210_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_212_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_212_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_212_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_212_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_213_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_213_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_213_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_213_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_215_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_215_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_215_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_215_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_217_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_217_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_217_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_217_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_218_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_218_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_218_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_218_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_220_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_220_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_220_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_220_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_222_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_222_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_222_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_222_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_223_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_223_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_223_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_223_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_225_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_225_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_225_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_225_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_227_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_227_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_227_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_227_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_228_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_228_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_228_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_228_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_230_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_230_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_230_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_230_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_232_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_232_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_232_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_232_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_233_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_233_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_233_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_233_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_235_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_235_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_235_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_235_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_237_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_237_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_237_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_237_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_238_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_238_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_238_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_238_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_240_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_240_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_240_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_240_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_242_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_242_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_242_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_242_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_243_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_243_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_243_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_243_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_245_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_245_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_245_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_245_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_247_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_247_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_247_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_247_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_248_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_248_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_248_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_248_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_250_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_250_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_250_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_250_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_252_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_252_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_252_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_252_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_253_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_253_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_253_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_253_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_255_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_255_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_255_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_255_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_257_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_257_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_257_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_257_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_258_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_258_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_258_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_258_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_260_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_260_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_260_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_260_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_262_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_262_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_262_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_262_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_263_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_263_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_263_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_263_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_265_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_265_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_265_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_265_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_267_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_267_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_267_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_267_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_268_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_268_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_268_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_268_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_270_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_270_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_270_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_270_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_272_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_272_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_272_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_272_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_273_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_273_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_273_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_273_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_275_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_275_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_275_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_275_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_277_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_277_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_277_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_277_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_278_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_278_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_278_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_278_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_280_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_280_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_280_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_280_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_282_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_282_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_282_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_282_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_283_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_283_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_283_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_283_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_285_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_285_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_285_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_285_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_287_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_287_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_287_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_287_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_288_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_288_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_288_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_288_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_290_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_290_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_290_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_290_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_292_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_292_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_292_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_292_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_293_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_293_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_293_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_293_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_295_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_295_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_295_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_295_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_297_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_297_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_297_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_297_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_298_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_298_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_298_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_298_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_300_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_300_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_300_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_300_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_302_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_302_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_302_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_302_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_303_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_303_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_303_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_303_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_305_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_305_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_305_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_305_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_307_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_307_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_307_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_307_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_308_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_308_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_308_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_308_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_310_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_310_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_310_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_310_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_312_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_312_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_312_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_312_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_313_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_313_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_313_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_313_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_315_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_315_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_315_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_315_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_317_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_317_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_317_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_317_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_318_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_318_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_318_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_318_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_320_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_320_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_320_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_320_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_322_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_322_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_322_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_322_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_323_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_323_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_323_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_323_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_325_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_325_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_325_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_325_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_327_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_327_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_327_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_327_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_328_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_328_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_328_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_328_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_330_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_330_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_330_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_330_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_332_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_332_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_332_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_332_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_333_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_333_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_333_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_333_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_335_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_335_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_335_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_335_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_337_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_337_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_337_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_337_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_338_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_338_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_338_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_338_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_340_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_340_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_340_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_340_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_342_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_342_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_342_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_342_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_343_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_343_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_343_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_343_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_345_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_345_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_345_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_345_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_347_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_347_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_347_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_347_en; // @[lut_35.scala 216:26]
  wire [32:0] LUT_mem_MPORT_348_data; // @[lut_35.scala 216:26]
  wire [5:0] LUT_mem_MPORT_348_addr; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_348_mask; // @[lut_35.scala 216:26]
  wire  LUT_mem_MPORT_348_en; // @[lut_35.scala 216:26]
  reg [31:0] read_stack0; // @[lut_35.scala 217:30]
  reg [31:0] read_stack1; // @[lut_35.scala 218:30]
  reg [31:0] read_stack2; // @[lut_35.scala 219:30]
  reg [31:0] read_stack3; // @[lut_35.scala 220:30]
  reg [31:0] read_stack4; // @[lut_35.scala 221:30]
  reg [31:0] read_stack5; // @[lut_35.scala 222:30]
  reg [31:0] read_stack6; // @[lut_35.scala 223:30]
  reg [31:0] read_stack7; // @[lut_35.scala 224:30]
  reg [31:0] read_stack8; // @[lut_35.scala 225:30]
  reg [31:0] read_stack9; // @[lut_35.scala 226:30]
  reg [31:0] read_stack10; // @[lut_35.scala 227:31]
  reg [31:0] read_stack11; // @[lut_35.scala 228:31]
  reg [31:0] read_stack12; // @[lut_35.scala 229:31]
  reg [31:0] read_stack13; // @[lut_35.scala 230:31]
  reg [31:0] read_stack14; // @[lut_35.scala 231:31]
  reg [31:0] read_stack15; // @[lut_35.scala 232:31]
  reg [31:0] read_stack16; // @[lut_35.scala 233:31]
  reg [31:0] read_stack17; // @[lut_35.scala 234:31]
  reg [31:0] read_stack18; // @[lut_35.scala 235:31]
  reg [31:0] read_stack19; // @[lut_35.scala 236:31]
  reg [31:0] read_stack20; // @[lut_35.scala 237:31]
  reg [31:0] read_stack21; // @[lut_35.scala 238:31]
  reg [31:0] read_stack22; // @[lut_35.scala 239:31]
  reg [31:0] read_stack23; // @[lut_35.scala 240:31]
  reg [31:0] read_stack24; // @[lut_35.scala 241:31]
  reg [31:0] read_stack25; // @[lut_35.scala 242:31]
  reg [31:0] read_stack26; // @[lut_35.scala 243:31]
  reg [31:0] read_stack27; // @[lut_35.scala 244:31]
  reg [31:0] read_stack28; // @[lut_35.scala 245:31]
  reg [31:0] read_stack29; // @[lut_35.scala 246:31]
  reg [31:0] read_stack30; // @[lut_35.scala 247:31]
  reg [31:0] read_stack31; // @[lut_35.scala 248:31]
  reg [31:0] read_stack32; // @[lut_35.scala 249:31]
  reg [31:0] read_stack33; // @[lut_35.scala 250:31]
  reg [31:0] read_stack34; // @[lut_35.scala 251:31]
  reg  push_0_1; // @[lut_35.scala 253:31]
  reg  push_1_1; // @[lut_35.scala 254:31]
  reg  push_2_1; // @[lut_35.scala 255:31]
  reg  push_3_1; // @[lut_35.scala 256:31]
  reg  push_4_1; // @[lut_35.scala 257:31]
  reg  push_5_1; // @[lut_35.scala 258:31]
  reg  push_6_1; // @[lut_35.scala 259:31]
  reg  push_7_1; // @[lut_35.scala 260:31]
  reg  push_8_1; // @[lut_35.scala 261:31]
  reg  push_9_1; // @[lut_35.scala 262:31]
  reg  push_10_1; // @[lut_35.scala 263:32]
  reg  push_11_1; // @[lut_35.scala 264:32]
  reg  push_12_1; // @[lut_35.scala 265:32]
  reg  push_13_1; // @[lut_35.scala 266:32]
  reg  push_14_1; // @[lut_35.scala 267:32]
  reg  push_15_1; // @[lut_35.scala 268:32]
  reg  push_16_1; // @[lut_35.scala 269:32]
  reg  push_17_1; // @[lut_35.scala 270:32]
  reg  push_18_1; // @[lut_35.scala 271:32]
  reg  push_19_1; // @[lut_35.scala 272:32]
  reg  push_20_1; // @[lut_35.scala 273:32]
  reg  push_21_1; // @[lut_35.scala 274:32]
  reg  push_22_1; // @[lut_35.scala 275:32]
  reg  push_23_1; // @[lut_35.scala 276:32]
  reg  push_24_1; // @[lut_35.scala 277:32]
  reg  push_25_1; // @[lut_35.scala 278:32]
  reg  push_26_1; // @[lut_35.scala 279:32]
  reg  push_27_1; // @[lut_35.scala 280:32]
  reg  push_28_1; // @[lut_35.scala 281:32]
  reg  push_29_1; // @[lut_35.scala 282:32]
  reg  push_30_1; // @[lut_35.scala 283:32]
  reg  push_31_1; // @[lut_35.scala 284:32]
  reg  push_32_1; // @[lut_35.scala 285:32]
  reg  push_33_1; // @[lut_35.scala 286:32]
  reg  push_34_1; // @[lut_35.scala 287:32]
  reg  push_1; // @[lut_35.scala 291:40]
  reg  push_valid; // @[lut_35.scala 292:41]
  reg [31:0] push_ray_id; // @[lut_35.scala 294:41]
  reg  push_valid_2; // @[lut_35.scala 334:41]
  reg  dispatch_reg_0; // @[lut_35.scala 340:33]
  reg  dispatch_reg_1; // @[lut_35.scala 341:33]
  reg  dispatch_reg_2; // @[lut_35.scala 342:33]
  reg  dispatch_reg_3; // @[lut_35.scala 343:33]
  reg  dispatch_reg_4; // @[lut_35.scala 344:33]
  reg  dispatch_reg_5; // @[lut_35.scala 345:33]
  reg  dispatch_reg_6; // @[lut_35.scala 346:33]
  reg  dispatch_reg_7; // @[lut_35.scala 347:33]
  reg  dispatch_reg_8; // @[lut_35.scala 348:33]
  reg  dispatch_reg_9; // @[lut_35.scala 349:33]
  reg  dispatch_reg_10; // @[lut_35.scala 350:34]
  reg  dispatch_reg_11; // @[lut_35.scala 351:34]
  reg  dispatch_reg_12; // @[lut_35.scala 352:34]
  reg  dispatch_reg_13; // @[lut_35.scala 353:34]
  reg  dispatch_reg_14; // @[lut_35.scala 354:34]
  reg  dispatch_reg_15; // @[lut_35.scala 355:34]
  reg  dispatch_reg_16; // @[lut_35.scala 356:34]
  reg  dispatch_reg_17; // @[lut_35.scala 357:34]
  reg  dispatch_reg_18; // @[lut_35.scala 358:34]
  reg  dispatch_reg_19; // @[lut_35.scala 359:34]
  reg  dispatch_reg_20; // @[lut_35.scala 360:34]
  reg  dispatch_reg_21; // @[lut_35.scala 361:34]
  reg  dispatch_reg_22; // @[lut_35.scala 362:34]
  reg  dispatch_reg_23; // @[lut_35.scala 363:34]
  reg  dispatch_reg_24; // @[lut_35.scala 364:34]
  reg  dispatch_reg_25; // @[lut_35.scala 365:34]
  reg  dispatch_reg_26; // @[lut_35.scala 366:34]
  reg  dispatch_reg_27; // @[lut_35.scala 367:34]
  reg  dispatch_reg_28; // @[lut_35.scala 368:34]
  reg  dispatch_reg_29; // @[lut_35.scala 369:34]
  reg  dispatch_reg_30; // @[lut_35.scala 370:34]
  reg  dispatch_reg_31; // @[lut_35.scala 371:34]
  reg  dispatch_reg_32; // @[lut_35.scala 372:34]
  reg  dispatch_reg_33; // @[lut_35.scala 373:34]
  reg  dispatch_reg_34; // @[lut_35.scala 374:34]
  wire  _T_36 = io_push & io_push_valid; // @[lut_35.scala 501:29]
  wire  _GEN_3 = io_push & io_push_valid & io_push_valid; // @[lut_35.scala 501:46 lut_35.scala 506:28 lut_35.scala 508:28]
  reg [5:0] push_mem_temp; // @[lut_35.scala 521:39]
  reg [31:0] push_id_temp; // @[lut_35.scala 522:39]
  wire  _T_39 = push_1 & push_valid; // @[lut_35.scala 524:24]
  wire  _T_196 = read_stack0 != push_ray_id & read_stack1 != push_ray_id & read_stack2 != push_ray_id & read_stack3 !=
    push_ray_id & read_stack4 != push_ray_id & read_stack5 != push_ray_id & read_stack6 != push_ray_id & read_stack7 !=
    push_ray_id & read_stack8 != push_ray_id; // @[lut_35.scala 1855:264]
  wire  _T_210 = _T_196 & read_stack9 != push_ray_id & read_stack10 != push_ray_id & read_stack11 != push_ray_id &
    read_stack12 != push_ray_id & read_stack13 != push_ray_id & read_stack14 != push_ray_id & read_stack15 !=
    push_ray_id; // @[lut_35.scala 1856:194]
  wire  _T_222 = _T_210 & read_stack16 != push_ray_id & read_stack17 != push_ray_id & read_stack18 != push_ray_id &
    read_stack19 != push_ray_id & read_stack20 != push_ray_id & read_stack21 != push_ray_id; // @[lut_35.scala 1857:164]
  wire  _T_234 = _T_222 & read_stack22 != push_ray_id & read_stack23 != push_ray_id & read_stack24 != push_ray_id &
    read_stack25 != push_ray_id & read_stack26 != push_ray_id & read_stack27 != push_ray_id; // @[lut_35.scala 1858:165]
  wire  _T_242 = _T_234 & read_stack28 != push_ray_id & read_stack29 != push_ray_id & read_stack30 != push_ray_id &
    read_stack31 != push_ray_id; // @[lut_35.scala 1859:102]
  wire  _T_250 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid; // @[lut_35.scala 1860:102]
  wire  _T_258 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32]; // @[lut_35.scala 1861:78]
  wire  _T_266 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32]; // @[lut_35.scala 1903:78]
  wire  _T_274 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32]; // @[lut_35.scala 1945:78]
  wire  _T_282 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32]; // @[lut_35.scala 1987:78]
  wire  _T_290 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32]; // @[lut_35.scala 2029:78]
  wire  _T_298 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32]; // @[lut_35.scala 2071:78]
  wire  _T_306 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32]; // @[lut_35.scala 2113:78]
  wire  _T_314 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32]; // @[lut_35.scala 2155:78]
  wire  _T_322 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32]; // @[lut_35.scala 2197:78]
  wire  _T_330 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32]; // @[lut_35.scala 2239:78]
  wire  _T_338 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32]; // @[lut_35.scala 2281:80]
  wire  _T_346 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32]; // @[lut_35.scala 2323:80]
  wire  _T_354 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32]; // @[lut_35.scala 2365:80]
  wire  _T_362 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32]; // @[lut_35.scala 2407:80]
  wire  _T_370 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32]; // @[lut_35.scala 2449:80]
  wire  _T_378 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_85_data[32]; // @[lut_35.scala 2491:80]
  wire  _T_386 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_86_data[32]; // @[lut_35.scala 2533:80]
  wire  _T_394 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_87_data[32]; // @[lut_35.scala 2575:80]
  wire  _T_402 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_88_data[32]; // @[lut_35.scala 2617:80]
  wire  _T_410 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_89_data[32]; // @[lut_35.scala 2659:80]
  wire  _T_418 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_90_data[32]; // @[lut_35.scala 2701:80]
  wire  _T_426 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_91_data[32]; // @[lut_35.scala 2743:80]
  wire  _T_434 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_92_data[32]; // @[lut_35.scala 2785:80]
  wire  _T_442 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_93_data[32]; // @[lut_35.scala 2827:80]
  wire  _T_450 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_94_data[32]; // @[lut_35.scala 2870:80]
  wire  _T_458 = io_empty_25 & push_valid & ~push_25_1 & ~LUT_mem_MPORT_95_data[32]; // @[lut_35.scala 2912:82]
  wire  _T_466 = io_empty_26 & push_valid & ~push_26_1 & ~LUT_mem_MPORT_96_data[32]; // @[lut_35.scala 2954:82]
  wire  _T_474 = io_empty_27 & push_valid & ~push_27_1 & ~LUT_mem_MPORT_97_data[32]; // @[lut_35.scala 2996:81]
  wire  _T_482 = io_empty_28 & push_valid & ~push_28_1 & ~LUT_mem_MPORT_98_data[32]; // @[lut_35.scala 3038:81]
  wire  _T_490 = io_empty_29 & push_valid & ~push_29_1 & ~LUT_mem_MPORT_99_data[32]; // @[lut_35.scala 3080:81]
  wire  _T_498 = io_empty_30 & push_valid & ~push_30_1 & ~LUT_mem_MPORT_100_data[32]; // @[lut_35.scala 3122:81]
  wire  _T_506 = io_empty_31 & push_valid & ~push_31_1 & ~LUT_mem_MPORT_101_data[32]; // @[lut_35.scala 3164:81]
  wire  _T_514 = io_empty_32 & push_valid & ~push_32_1 & ~LUT_mem_MPORT_102_data[32]; // @[lut_35.scala 3206:81]
  wire  _T_522 = io_empty_33 & push_valid & ~push_33_1 & ~LUT_mem_MPORT_103_data[32]; // @[lut_35.scala 3248:80]
  wire  _T_530 = io_empty_34 & push_valid & ~push_34_1 & ~LUT_mem_MPORT_104_data[32]; // @[lut_35.scala 3290:80]
  wire [5:0] _GEN_4 = io_empty_34 & push_valid & ~push_34_1 & ~LUT_mem_MPORT_104_data[32] ? 6'h22 : 6'h23; // @[lut_35.scala 3290:105 lut_35.scala 3291:42 lut_35.scala 3333:42]
  wire [31:0] _GEN_5 = io_empty_34 & push_valid & ~push_34_1 & ~LUT_mem_MPORT_104_data[32] ? push_ray_id : 32'h0; // @[lut_35.scala 3290:105 lut_35.scala 3292:42 lut_35.scala 3334:42]
  wire [5:0] _GEN_9 = io_empty_33 & push_valid & ~push_33_1 & ~LUT_mem_MPORT_103_data[32] ? 6'h21 : _GEN_4; // @[lut_35.scala 3248:105 lut_35.scala 3249:42]
  wire [31:0] _GEN_10 = io_empty_33 & push_valid & ~push_33_1 & ~LUT_mem_MPORT_103_data[32] ? push_ray_id : _GEN_5; // @[lut_35.scala 3248:105 lut_35.scala 3250:42]
  wire  _GEN_13 = io_empty_33 & push_valid & ~push_33_1 & ~LUT_mem_MPORT_103_data[32] ? 1'h0 : _T_530; // @[lut_35.scala 3248:105 lut_35.scala 3287:43]
  wire  _GEN_14 = io_empty_33 & push_valid & ~push_33_1 & ~LUT_mem_MPORT_103_data[32] | _T_530; // @[lut_35.scala 3248:105 lut_35.scala 3288:38]
  wire  _GEN_18 = io_empty_33 & push_valid & ~push_33_1 & ~LUT_mem_MPORT_103_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 3248:105 lut_35.scala 216:26 lut_35.scala 3290:89]
  wire [5:0] _GEN_19 = io_empty_32 & push_valid & ~push_32_1 & ~LUT_mem_MPORT_102_data[32] ? 6'h20 : _GEN_9; // @[lut_35.scala 3206:106 lut_35.scala 3207:42]
  wire [31:0] _GEN_20 = io_empty_32 & push_valid & ~push_32_1 & ~LUT_mem_MPORT_102_data[32] ? push_ray_id : _GEN_10; // @[lut_35.scala 3206:106 lut_35.scala 3208:42]
  wire  _GEN_23 = io_empty_32 & push_valid & ~push_32_1 & ~LUT_mem_MPORT_102_data[32] ? 1'h0 : _T_522; // @[lut_35.scala 3206:106 lut_35.scala 3244:43]
  wire  _GEN_24 = io_empty_32 & push_valid & ~push_32_1 & ~LUT_mem_MPORT_102_data[32] ? 1'h0 : _GEN_13; // @[lut_35.scala 3206:106 lut_35.scala 3245:43]
  wire  _GEN_25 = io_empty_32 & push_valid & ~push_32_1 & ~LUT_mem_MPORT_102_data[32] | _GEN_14; // @[lut_35.scala 3206:106 lut_35.scala 3246:38]
  wire  _GEN_29 = io_empty_32 & push_valid & ~push_32_1 & ~LUT_mem_MPORT_102_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 3206:106 lut_35.scala 216:26 lut_35.scala 3248:89]
  wire  _GEN_32 = io_empty_32 & push_valid & ~push_32_1 & ~LUT_mem_MPORT_102_data[32] ? 1'h0 : _GEN_18; // @[lut_35.scala 3206:106 lut_35.scala 216:26]
  wire [5:0] _GEN_33 = io_empty_31 & push_valid & ~push_31_1 & ~LUT_mem_MPORT_101_data[32] ? 6'h1f : _GEN_19; // @[lut_35.scala 3164:106 lut_35.scala 3165:42]
  wire [31:0] _GEN_34 = io_empty_31 & push_valid & ~push_31_1 & ~LUT_mem_MPORT_101_data[32] ? push_ray_id : _GEN_20; // @[lut_35.scala 3164:106 lut_35.scala 3166:42]
  wire  _GEN_37 = io_empty_31 & push_valid & ~push_31_1 & ~LUT_mem_MPORT_101_data[32] ? 1'h0 : _T_514; // @[lut_35.scala 3164:106 lut_35.scala 3201:43]
  wire  _GEN_38 = io_empty_31 & push_valid & ~push_31_1 & ~LUT_mem_MPORT_101_data[32] ? 1'h0 : _GEN_23; // @[lut_35.scala 3164:106 lut_35.scala 3202:43]
  wire  _GEN_39 = io_empty_31 & push_valid & ~push_31_1 & ~LUT_mem_MPORT_101_data[32] ? 1'h0 : _GEN_24; // @[lut_35.scala 3164:106 lut_35.scala 3203:43]
  wire  _GEN_40 = io_empty_31 & push_valid & ~push_31_1 & ~LUT_mem_MPORT_101_data[32] | _GEN_25; // @[lut_35.scala 3164:106 lut_35.scala 3204:38]
  wire  _GEN_44 = io_empty_31 & push_valid & ~push_31_1 & ~LUT_mem_MPORT_101_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 3164:106 lut_35.scala 216:26 lut_35.scala 3206:90]
  wire  _GEN_47 = io_empty_31 & push_valid & ~push_31_1 & ~LUT_mem_MPORT_101_data[32] ? 1'h0 : _GEN_29; // @[lut_35.scala 3164:106 lut_35.scala 216:26]
  wire  _GEN_50 = io_empty_31 & push_valid & ~push_31_1 & ~LUT_mem_MPORT_101_data[32] ? 1'h0 : _GEN_32; // @[lut_35.scala 3164:106 lut_35.scala 216:26]
  wire [5:0] _GEN_51 = io_empty_30 & push_valid & ~push_30_1 & ~LUT_mem_MPORT_100_data[32] ? 6'h1e : _GEN_33; // @[lut_35.scala 3122:106 lut_35.scala 3123:42]
  wire [31:0] _GEN_52 = io_empty_30 & push_valid & ~push_30_1 & ~LUT_mem_MPORT_100_data[32] ? push_ray_id : _GEN_34; // @[lut_35.scala 3122:106 lut_35.scala 3124:42]
  wire  _GEN_55 = io_empty_30 & push_valid & ~push_30_1 & ~LUT_mem_MPORT_100_data[32] ? 1'h0 : _T_506; // @[lut_35.scala 3122:106 lut_35.scala 3158:43]
  wire  _GEN_56 = io_empty_30 & push_valid & ~push_30_1 & ~LUT_mem_MPORT_100_data[32] ? 1'h0 : _GEN_37; // @[lut_35.scala 3122:106 lut_35.scala 3159:43]
  wire  _GEN_57 = io_empty_30 & push_valid & ~push_30_1 & ~LUT_mem_MPORT_100_data[32] ? 1'h0 : _GEN_38; // @[lut_35.scala 3122:106 lut_35.scala 3160:43]
  wire  _GEN_58 = io_empty_30 & push_valid & ~push_30_1 & ~LUT_mem_MPORT_100_data[32] ? 1'h0 : _GEN_39; // @[lut_35.scala 3122:106 lut_35.scala 3161:43]
  wire  _GEN_59 = io_empty_30 & push_valid & ~push_30_1 & ~LUT_mem_MPORT_100_data[32] | _GEN_40; // @[lut_35.scala 3122:106 lut_35.scala 3162:38]
  wire  _GEN_63 = io_empty_30 & push_valid & ~push_30_1 & ~LUT_mem_MPORT_100_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 3122:106 lut_35.scala 216:26 lut_35.scala 3164:90]
  wire  _GEN_66 = io_empty_30 & push_valid & ~push_30_1 & ~LUT_mem_MPORT_100_data[32] ? 1'h0 : _GEN_44; // @[lut_35.scala 3122:106 lut_35.scala 216:26]
  wire  _GEN_69 = io_empty_30 & push_valid & ~push_30_1 & ~LUT_mem_MPORT_100_data[32] ? 1'h0 : _GEN_47; // @[lut_35.scala 3122:106 lut_35.scala 216:26]
  wire  _GEN_72 = io_empty_30 & push_valid & ~push_30_1 & ~LUT_mem_MPORT_100_data[32] ? 1'h0 : _GEN_50; // @[lut_35.scala 3122:106 lut_35.scala 216:26]
  wire [5:0] _GEN_73 = io_empty_29 & push_valid & ~push_29_1 & ~LUT_mem_MPORT_99_data[32] ? 6'h1d : _GEN_51; // @[lut_35.scala 3080:106 lut_35.scala 3081:42]
  wire [31:0] _GEN_74 = io_empty_29 & push_valid & ~push_29_1 & ~LUT_mem_MPORT_99_data[32] ? push_ray_id : _GEN_52; // @[lut_35.scala 3080:106 lut_35.scala 3082:42]
  wire  _GEN_77 = io_empty_29 & push_valid & ~push_29_1 & ~LUT_mem_MPORT_99_data[32] ? 1'h0 : _T_498; // @[lut_35.scala 3080:106 lut_35.scala 3115:43]
  wire  _GEN_78 = io_empty_29 & push_valid & ~push_29_1 & ~LUT_mem_MPORT_99_data[32] ? 1'h0 : _GEN_55; // @[lut_35.scala 3080:106 lut_35.scala 3116:43]
  wire  _GEN_79 = io_empty_29 & push_valid & ~push_29_1 & ~LUT_mem_MPORT_99_data[32] ? 1'h0 : _GEN_56; // @[lut_35.scala 3080:106 lut_35.scala 3117:43]
  wire  _GEN_80 = io_empty_29 & push_valid & ~push_29_1 & ~LUT_mem_MPORT_99_data[32] ? 1'h0 : _GEN_57; // @[lut_35.scala 3080:106 lut_35.scala 3118:43]
  wire  _GEN_81 = io_empty_29 & push_valid & ~push_29_1 & ~LUT_mem_MPORT_99_data[32] ? 1'h0 : _GEN_58; // @[lut_35.scala 3080:106 lut_35.scala 3119:43]
  wire  _GEN_82 = io_empty_29 & push_valid & ~push_29_1 & ~LUT_mem_MPORT_99_data[32] | _GEN_59; // @[lut_35.scala 3080:106 lut_35.scala 3120:38]
  wire  _GEN_86 = io_empty_29 & push_valid & ~push_29_1 & ~LUT_mem_MPORT_99_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 3080:106 lut_35.scala 216:26 lut_35.scala 3122:90]
  wire  _GEN_89 = io_empty_29 & push_valid & ~push_29_1 & ~LUT_mem_MPORT_99_data[32] ? 1'h0 : _GEN_63; // @[lut_35.scala 3080:106 lut_35.scala 216:26]
  wire  _GEN_92 = io_empty_29 & push_valid & ~push_29_1 & ~LUT_mem_MPORT_99_data[32] ? 1'h0 : _GEN_66; // @[lut_35.scala 3080:106 lut_35.scala 216:26]
  wire  _GEN_95 = io_empty_29 & push_valid & ~push_29_1 & ~LUT_mem_MPORT_99_data[32] ? 1'h0 : _GEN_69; // @[lut_35.scala 3080:106 lut_35.scala 216:26]
  wire  _GEN_98 = io_empty_29 & push_valid & ~push_29_1 & ~LUT_mem_MPORT_99_data[32] ? 1'h0 : _GEN_72; // @[lut_35.scala 3080:106 lut_35.scala 216:26]
  wire [5:0] _GEN_99 = io_empty_28 & push_valid & ~push_28_1 & ~LUT_mem_MPORT_98_data[32] ? 6'h1c : _GEN_73; // @[lut_35.scala 3038:106 lut_35.scala 3039:42]
  wire [31:0] _GEN_100 = io_empty_28 & push_valid & ~push_28_1 & ~LUT_mem_MPORT_98_data[32] ? push_ray_id : _GEN_74; // @[lut_35.scala 3038:106 lut_35.scala 3040:42]
  wire  _GEN_103 = io_empty_28 & push_valid & ~push_28_1 & ~LUT_mem_MPORT_98_data[32] ? 1'h0 : _T_490; // @[lut_35.scala 3038:106 lut_35.scala 3072:43]
  wire  _GEN_104 = io_empty_28 & push_valid & ~push_28_1 & ~LUT_mem_MPORT_98_data[32] ? 1'h0 : _GEN_77; // @[lut_35.scala 3038:106 lut_35.scala 3073:43]
  wire  _GEN_105 = io_empty_28 & push_valid & ~push_28_1 & ~LUT_mem_MPORT_98_data[32] ? 1'h0 : _GEN_78; // @[lut_35.scala 3038:106 lut_35.scala 3074:43]
  wire  _GEN_106 = io_empty_28 & push_valid & ~push_28_1 & ~LUT_mem_MPORT_98_data[32] ? 1'h0 : _GEN_79; // @[lut_35.scala 3038:106 lut_35.scala 3075:43]
  wire  _GEN_107 = io_empty_28 & push_valid & ~push_28_1 & ~LUT_mem_MPORT_98_data[32] ? 1'h0 : _GEN_80; // @[lut_35.scala 3038:106 lut_35.scala 3076:43]
  wire  _GEN_108 = io_empty_28 & push_valid & ~push_28_1 & ~LUT_mem_MPORT_98_data[32] ? 1'h0 : _GEN_81; // @[lut_35.scala 3038:106 lut_35.scala 3077:43]
  wire  _GEN_109 = io_empty_28 & push_valid & ~push_28_1 & ~LUT_mem_MPORT_98_data[32] | _GEN_82; // @[lut_35.scala 3038:106 lut_35.scala 3078:38]
  wire  _GEN_113 = io_empty_28 & push_valid & ~push_28_1 & ~LUT_mem_MPORT_98_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 3038:106 lut_35.scala 216:26 lut_35.scala 3080:90]
  wire  _GEN_116 = io_empty_28 & push_valid & ~push_28_1 & ~LUT_mem_MPORT_98_data[32] ? 1'h0 : _GEN_86; // @[lut_35.scala 3038:106 lut_35.scala 216:26]
  wire  _GEN_119 = io_empty_28 & push_valid & ~push_28_1 & ~LUT_mem_MPORT_98_data[32] ? 1'h0 : _GEN_89; // @[lut_35.scala 3038:106 lut_35.scala 216:26]
  wire  _GEN_122 = io_empty_28 & push_valid & ~push_28_1 & ~LUT_mem_MPORT_98_data[32] ? 1'h0 : _GEN_92; // @[lut_35.scala 3038:106 lut_35.scala 216:26]
  wire  _GEN_125 = io_empty_28 & push_valid & ~push_28_1 & ~LUT_mem_MPORT_98_data[32] ? 1'h0 : _GEN_95; // @[lut_35.scala 3038:106 lut_35.scala 216:26]
  wire  _GEN_128 = io_empty_28 & push_valid & ~push_28_1 & ~LUT_mem_MPORT_98_data[32] ? 1'h0 : _GEN_98; // @[lut_35.scala 3038:106 lut_35.scala 216:26]
  wire [5:0] _GEN_129 = io_empty_27 & push_valid & ~push_27_1 & ~LUT_mem_MPORT_97_data[32] ? 6'h1b : _GEN_99; // @[lut_35.scala 2996:106 lut_35.scala 2997:42]
  wire [31:0] _GEN_130 = io_empty_27 & push_valid & ~push_27_1 & ~LUT_mem_MPORT_97_data[32] ? push_ray_id : _GEN_100; // @[lut_35.scala 2996:106 lut_35.scala 2998:42]
  wire  _GEN_133 = io_empty_27 & push_valid & ~push_27_1 & ~LUT_mem_MPORT_97_data[32] ? 1'h0 : _T_482; // @[lut_35.scala 2996:106 lut_35.scala 3029:43]
  wire  _GEN_134 = io_empty_27 & push_valid & ~push_27_1 & ~LUT_mem_MPORT_97_data[32] ? 1'h0 : _GEN_103; // @[lut_35.scala 2996:106 lut_35.scala 3030:43]
  wire  _GEN_135 = io_empty_27 & push_valid & ~push_27_1 & ~LUT_mem_MPORT_97_data[32] ? 1'h0 : _GEN_104; // @[lut_35.scala 2996:106 lut_35.scala 3031:43]
  wire  _GEN_136 = io_empty_27 & push_valid & ~push_27_1 & ~LUT_mem_MPORT_97_data[32] ? 1'h0 : _GEN_105; // @[lut_35.scala 2996:106 lut_35.scala 3032:43]
  wire  _GEN_137 = io_empty_27 & push_valid & ~push_27_1 & ~LUT_mem_MPORT_97_data[32] ? 1'h0 : _GEN_106; // @[lut_35.scala 2996:106 lut_35.scala 3033:43]
  wire  _GEN_138 = io_empty_27 & push_valid & ~push_27_1 & ~LUT_mem_MPORT_97_data[32] ? 1'h0 : _GEN_107; // @[lut_35.scala 2996:106 lut_35.scala 3034:43]
  wire  _GEN_139 = io_empty_27 & push_valid & ~push_27_1 & ~LUT_mem_MPORT_97_data[32] ? 1'h0 : _GEN_108; // @[lut_35.scala 2996:106 lut_35.scala 3035:43]
  wire  _GEN_140 = io_empty_27 & push_valid & ~push_27_1 & ~LUT_mem_MPORT_97_data[32] | _GEN_109; // @[lut_35.scala 2996:106 lut_35.scala 3036:38]
  wire  _GEN_144 = io_empty_27 & push_valid & ~push_27_1 & ~LUT_mem_MPORT_97_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2996:106 lut_35.scala 216:26 lut_35.scala 3038:90]
  wire  _GEN_147 = io_empty_27 & push_valid & ~push_27_1 & ~LUT_mem_MPORT_97_data[32] ? 1'h0 : _GEN_113; // @[lut_35.scala 2996:106 lut_35.scala 216:26]
  wire  _GEN_150 = io_empty_27 & push_valid & ~push_27_1 & ~LUT_mem_MPORT_97_data[32] ? 1'h0 : _GEN_116; // @[lut_35.scala 2996:106 lut_35.scala 216:26]
  wire  _GEN_153 = io_empty_27 & push_valid & ~push_27_1 & ~LUT_mem_MPORT_97_data[32] ? 1'h0 : _GEN_119; // @[lut_35.scala 2996:106 lut_35.scala 216:26]
  wire  _GEN_156 = io_empty_27 & push_valid & ~push_27_1 & ~LUT_mem_MPORT_97_data[32] ? 1'h0 : _GEN_122; // @[lut_35.scala 2996:106 lut_35.scala 216:26]
  wire  _GEN_159 = io_empty_27 & push_valid & ~push_27_1 & ~LUT_mem_MPORT_97_data[32] ? 1'h0 : _GEN_125; // @[lut_35.scala 2996:106 lut_35.scala 216:26]
  wire  _GEN_162 = io_empty_27 & push_valid & ~push_27_1 & ~LUT_mem_MPORT_97_data[32] ? 1'h0 : _GEN_128; // @[lut_35.scala 2996:106 lut_35.scala 216:26]
  wire [5:0] _GEN_163 = io_empty_26 & push_valid & ~push_26_1 & ~LUT_mem_MPORT_96_data[32] ? 6'h1a : _GEN_129; // @[lut_35.scala 2954:107 lut_35.scala 2955:42]
  wire [31:0] _GEN_164 = io_empty_26 & push_valid & ~push_26_1 & ~LUT_mem_MPORT_96_data[32] ? push_ray_id : _GEN_130; // @[lut_35.scala 2954:107 lut_35.scala 2956:42]
  wire  _GEN_167 = io_empty_26 & push_valid & ~push_26_1 & ~LUT_mem_MPORT_96_data[32] ? 1'h0 : _T_474; // @[lut_35.scala 2954:107 lut_35.scala 2986:43]
  wire  _GEN_168 = io_empty_26 & push_valid & ~push_26_1 & ~LUT_mem_MPORT_96_data[32] ? 1'h0 : _GEN_133; // @[lut_35.scala 2954:107 lut_35.scala 2987:43]
  wire  _GEN_169 = io_empty_26 & push_valid & ~push_26_1 & ~LUT_mem_MPORT_96_data[32] ? 1'h0 : _GEN_134; // @[lut_35.scala 2954:107 lut_35.scala 2988:43]
  wire  _GEN_170 = io_empty_26 & push_valid & ~push_26_1 & ~LUT_mem_MPORT_96_data[32] ? 1'h0 : _GEN_135; // @[lut_35.scala 2954:107 lut_35.scala 2989:43]
  wire  _GEN_171 = io_empty_26 & push_valid & ~push_26_1 & ~LUT_mem_MPORT_96_data[32] ? 1'h0 : _GEN_136; // @[lut_35.scala 2954:107 lut_35.scala 2990:43]
  wire  _GEN_172 = io_empty_26 & push_valid & ~push_26_1 & ~LUT_mem_MPORT_96_data[32] ? 1'h0 : _GEN_137; // @[lut_35.scala 2954:107 lut_35.scala 2991:43]
  wire  _GEN_173 = io_empty_26 & push_valid & ~push_26_1 & ~LUT_mem_MPORT_96_data[32] ? 1'h0 : _GEN_138; // @[lut_35.scala 2954:107 lut_35.scala 2992:43]
  wire  _GEN_174 = io_empty_26 & push_valid & ~push_26_1 & ~LUT_mem_MPORT_96_data[32] ? 1'h0 : _GEN_139; // @[lut_35.scala 2954:107 lut_35.scala 2993:43]
  wire  _GEN_175 = io_empty_26 & push_valid & ~push_26_1 & ~LUT_mem_MPORT_96_data[32] | _GEN_140; // @[lut_35.scala 2954:107 lut_35.scala 2994:38]
  wire  _GEN_179 = io_empty_26 & push_valid & ~push_26_1 & ~LUT_mem_MPORT_96_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2954:107 lut_35.scala 216:26 lut_35.scala 2996:90]
  wire  _GEN_182 = io_empty_26 & push_valid & ~push_26_1 & ~LUT_mem_MPORT_96_data[32] ? 1'h0 : _GEN_144; // @[lut_35.scala 2954:107 lut_35.scala 216:26]
  wire  _GEN_185 = io_empty_26 & push_valid & ~push_26_1 & ~LUT_mem_MPORT_96_data[32] ? 1'h0 : _GEN_147; // @[lut_35.scala 2954:107 lut_35.scala 216:26]
  wire  _GEN_188 = io_empty_26 & push_valid & ~push_26_1 & ~LUT_mem_MPORT_96_data[32] ? 1'h0 : _GEN_150; // @[lut_35.scala 2954:107 lut_35.scala 216:26]
  wire  _GEN_191 = io_empty_26 & push_valid & ~push_26_1 & ~LUT_mem_MPORT_96_data[32] ? 1'h0 : _GEN_153; // @[lut_35.scala 2954:107 lut_35.scala 216:26]
  wire  _GEN_194 = io_empty_26 & push_valid & ~push_26_1 & ~LUT_mem_MPORT_96_data[32] ? 1'h0 : _GEN_156; // @[lut_35.scala 2954:107 lut_35.scala 216:26]
  wire  _GEN_197 = io_empty_26 & push_valid & ~push_26_1 & ~LUT_mem_MPORT_96_data[32] ? 1'h0 : _GEN_159; // @[lut_35.scala 2954:107 lut_35.scala 216:26]
  wire  _GEN_200 = io_empty_26 & push_valid & ~push_26_1 & ~LUT_mem_MPORT_96_data[32] ? 1'h0 : _GEN_162; // @[lut_35.scala 2954:107 lut_35.scala 216:26]
  wire [5:0] _GEN_201 = io_empty_25 & push_valid & ~push_25_1 & ~LUT_mem_MPORT_95_data[32] ? 6'h19 : _GEN_163; // @[lut_35.scala 2912:107 lut_35.scala 2913:42]
  wire [31:0] _GEN_202 = io_empty_25 & push_valid & ~push_25_1 & ~LUT_mem_MPORT_95_data[32] ? push_ray_id : _GEN_164; // @[lut_35.scala 2912:107 lut_35.scala 2914:42]
  wire  _GEN_205 = io_empty_25 & push_valid & ~push_25_1 & ~LUT_mem_MPORT_95_data[32] ? 1'h0 : _T_466; // @[lut_35.scala 2912:107 lut_35.scala 2943:43]
  wire  _GEN_206 = io_empty_25 & push_valid & ~push_25_1 & ~LUT_mem_MPORT_95_data[32] ? 1'h0 : _GEN_167; // @[lut_35.scala 2912:107 lut_35.scala 2944:43]
  wire  _GEN_207 = io_empty_25 & push_valid & ~push_25_1 & ~LUT_mem_MPORT_95_data[32] ? 1'h0 : _GEN_168; // @[lut_35.scala 2912:107 lut_35.scala 2945:43]
  wire  _GEN_208 = io_empty_25 & push_valid & ~push_25_1 & ~LUT_mem_MPORT_95_data[32] ? 1'h0 : _GEN_169; // @[lut_35.scala 2912:107 lut_35.scala 2946:43]
  wire  _GEN_209 = io_empty_25 & push_valid & ~push_25_1 & ~LUT_mem_MPORT_95_data[32] ? 1'h0 : _GEN_170; // @[lut_35.scala 2912:107 lut_35.scala 2947:43]
  wire  _GEN_210 = io_empty_25 & push_valid & ~push_25_1 & ~LUT_mem_MPORT_95_data[32] ? 1'h0 : _GEN_171; // @[lut_35.scala 2912:107 lut_35.scala 2948:43]
  wire  _GEN_211 = io_empty_25 & push_valid & ~push_25_1 & ~LUT_mem_MPORT_95_data[32] ? 1'h0 : _GEN_172; // @[lut_35.scala 2912:107 lut_35.scala 2949:43]
  wire  _GEN_212 = io_empty_25 & push_valid & ~push_25_1 & ~LUT_mem_MPORT_95_data[32] ? 1'h0 : _GEN_173; // @[lut_35.scala 2912:107 lut_35.scala 2950:43]
  wire  _GEN_213 = io_empty_25 & push_valid & ~push_25_1 & ~LUT_mem_MPORT_95_data[32] ? 1'h0 : _GEN_174; // @[lut_35.scala 2912:107 lut_35.scala 2951:43]
  wire  _GEN_214 = io_empty_25 & push_valid & ~push_25_1 & ~LUT_mem_MPORT_95_data[32] | _GEN_175; // @[lut_35.scala 2912:107 lut_35.scala 2952:38]
  wire  _GEN_218 = io_empty_25 & push_valid & ~push_25_1 & ~LUT_mem_MPORT_95_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2912:107 lut_35.scala 216:26 lut_35.scala 2954:91]
  wire  _GEN_221 = io_empty_25 & push_valid & ~push_25_1 & ~LUT_mem_MPORT_95_data[32] ? 1'h0 : _GEN_179; // @[lut_35.scala 2912:107 lut_35.scala 216:26]
  wire  _GEN_224 = io_empty_25 & push_valid & ~push_25_1 & ~LUT_mem_MPORT_95_data[32] ? 1'h0 : _GEN_182; // @[lut_35.scala 2912:107 lut_35.scala 216:26]
  wire  _GEN_227 = io_empty_25 & push_valid & ~push_25_1 & ~LUT_mem_MPORT_95_data[32] ? 1'h0 : _GEN_185; // @[lut_35.scala 2912:107 lut_35.scala 216:26]
  wire  _GEN_230 = io_empty_25 & push_valid & ~push_25_1 & ~LUT_mem_MPORT_95_data[32] ? 1'h0 : _GEN_188; // @[lut_35.scala 2912:107 lut_35.scala 216:26]
  wire  _GEN_233 = io_empty_25 & push_valid & ~push_25_1 & ~LUT_mem_MPORT_95_data[32] ? 1'h0 : _GEN_191; // @[lut_35.scala 2912:107 lut_35.scala 216:26]
  wire  _GEN_236 = io_empty_25 & push_valid & ~push_25_1 & ~LUT_mem_MPORT_95_data[32] ? 1'h0 : _GEN_194; // @[lut_35.scala 2912:107 lut_35.scala 216:26]
  wire  _GEN_239 = io_empty_25 & push_valid & ~push_25_1 & ~LUT_mem_MPORT_95_data[32] ? 1'h0 : _GEN_197; // @[lut_35.scala 2912:107 lut_35.scala 216:26]
  wire  _GEN_242 = io_empty_25 & push_valid & ~push_25_1 & ~LUT_mem_MPORT_95_data[32] ? 1'h0 : _GEN_200; // @[lut_35.scala 2912:107 lut_35.scala 216:26]
  wire [5:0] _GEN_243 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_94_data[32] ? 6'h18 : _GEN_201; // @[lut_35.scala 2870:105 lut_35.scala 2871:42]
  wire [31:0] _GEN_244 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_94_data[32] ? push_ray_id : _GEN_202; // @[lut_35.scala 2870:105 lut_35.scala 2872:42]
  wire  _GEN_247 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_94_data[32] ? 1'h0 : _T_458; // @[lut_35.scala 2870:105 lut_35.scala 2900:43]
  wire  _GEN_248 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_94_data[32] ? 1'h0 : _GEN_205; // @[lut_35.scala 2870:105 lut_35.scala 2901:43]
  wire  _GEN_249 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_94_data[32] ? 1'h0 : _GEN_206; // @[lut_35.scala 2870:105 lut_35.scala 2902:43]
  wire  _GEN_250 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_94_data[32] ? 1'h0 : _GEN_207; // @[lut_35.scala 2870:105 lut_35.scala 2903:43]
  wire  _GEN_251 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_94_data[32] ? 1'h0 : _GEN_208; // @[lut_35.scala 2870:105 lut_35.scala 2904:43]
  wire  _GEN_252 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_94_data[32] ? 1'h0 : _GEN_209; // @[lut_35.scala 2870:105 lut_35.scala 2905:43]
  wire  _GEN_253 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_94_data[32] ? 1'h0 : _GEN_210; // @[lut_35.scala 2870:105 lut_35.scala 2906:43]
  wire  _GEN_254 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_94_data[32] ? 1'h0 : _GEN_211; // @[lut_35.scala 2870:105 lut_35.scala 2907:43]
  wire  _GEN_255 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_94_data[32] ? 1'h0 : _GEN_212; // @[lut_35.scala 2870:105 lut_35.scala 2908:43]
  wire  _GEN_256 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_94_data[32] ? 1'h0 : _GEN_213; // @[lut_35.scala 2870:105 lut_35.scala 2909:43]
  wire  _GEN_257 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_94_data[32] | _GEN_214; // @[lut_35.scala 2870:105 lut_35.scala 2910:38]
  wire  _GEN_261 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_94_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2870:105 lut_35.scala 216:26 lut_35.scala 2912:91]
  wire  _GEN_264 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_94_data[32] ? 1'h0 : _GEN_218; // @[lut_35.scala 2870:105 lut_35.scala 216:26]
  wire  _GEN_267 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_94_data[32] ? 1'h0 : _GEN_221; // @[lut_35.scala 2870:105 lut_35.scala 216:26]
  wire  _GEN_270 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_94_data[32] ? 1'h0 : _GEN_224; // @[lut_35.scala 2870:105 lut_35.scala 216:26]
  wire  _GEN_273 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_94_data[32] ? 1'h0 : _GEN_227; // @[lut_35.scala 2870:105 lut_35.scala 216:26]
  wire  _GEN_276 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_94_data[32] ? 1'h0 : _GEN_230; // @[lut_35.scala 2870:105 lut_35.scala 216:26]
  wire  _GEN_279 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_94_data[32] ? 1'h0 : _GEN_233; // @[lut_35.scala 2870:105 lut_35.scala 216:26]
  wire  _GEN_282 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_94_data[32] ? 1'h0 : _GEN_236; // @[lut_35.scala 2870:105 lut_35.scala 216:26]
  wire  _GEN_285 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_94_data[32] ? 1'h0 : _GEN_239; // @[lut_35.scala 2870:105 lut_35.scala 216:26]
  wire  _GEN_288 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_94_data[32] ? 1'h0 : _GEN_242; // @[lut_35.scala 2870:105 lut_35.scala 216:26]
  wire [5:0] _GEN_289 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_93_data[32] ? 6'h17 : _GEN_243; // @[lut_35.scala 2827:105 lut_35.scala 2828:42]
  wire [31:0] _GEN_290 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_93_data[32] ? push_ray_id : _GEN_244; // @[lut_35.scala 2827:105 lut_35.scala 2829:42]
  wire  _GEN_293 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_93_data[32] ? 1'h0 : _T_450; // @[lut_35.scala 2827:105 lut_35.scala 2856:43]
  wire  _GEN_294 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_93_data[32] ? 1'h0 : _GEN_247; // @[lut_35.scala 2827:105 lut_35.scala 2857:43]
  wire  _GEN_295 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_93_data[32] ? 1'h0 : _GEN_248; // @[lut_35.scala 2827:105 lut_35.scala 2858:43]
  wire  _GEN_296 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_93_data[32] ? 1'h0 : _GEN_249; // @[lut_35.scala 2827:105 lut_35.scala 2859:43]
  wire  _GEN_297 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_93_data[32] ? 1'h0 : _GEN_250; // @[lut_35.scala 2827:105 lut_35.scala 2860:43]
  wire  _GEN_298 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_93_data[32] ? 1'h0 : _GEN_251; // @[lut_35.scala 2827:105 lut_35.scala 2861:43]
  wire  _GEN_299 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_93_data[32] ? 1'h0 : _GEN_252; // @[lut_35.scala 2827:105 lut_35.scala 2862:43]
  wire  _GEN_300 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_93_data[32] ? 1'h0 : _GEN_253; // @[lut_35.scala 2827:105 lut_35.scala 2863:43]
  wire  _GEN_301 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_93_data[32] ? 1'h0 : _GEN_254; // @[lut_35.scala 2827:105 lut_35.scala 2864:43]
  wire  _GEN_302 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_93_data[32] ? 1'h0 : _GEN_255; // @[lut_35.scala 2827:105 lut_35.scala 2865:43]
  wire  _GEN_303 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_93_data[32] ? 1'h0 : _GEN_256; // @[lut_35.scala 2827:105 lut_35.scala 2866:43]
  wire  _GEN_304 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_93_data[32] | _GEN_257; // @[lut_35.scala 2827:105 lut_35.scala 2867:38]
  wire  _GEN_308 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_93_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2827:105 lut_35.scala 216:26 lut_35.scala 2870:89]
  wire  _GEN_311 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_93_data[32] ? 1'h0 : _GEN_261; // @[lut_35.scala 2827:105 lut_35.scala 216:26]
  wire  _GEN_314 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_93_data[32] ? 1'h0 : _GEN_264; // @[lut_35.scala 2827:105 lut_35.scala 216:26]
  wire  _GEN_317 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_93_data[32] ? 1'h0 : _GEN_267; // @[lut_35.scala 2827:105 lut_35.scala 216:26]
  wire  _GEN_320 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_93_data[32] ? 1'h0 : _GEN_270; // @[lut_35.scala 2827:105 lut_35.scala 216:26]
  wire  _GEN_323 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_93_data[32] ? 1'h0 : _GEN_273; // @[lut_35.scala 2827:105 lut_35.scala 216:26]
  wire  _GEN_326 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_93_data[32] ? 1'h0 : _GEN_276; // @[lut_35.scala 2827:105 lut_35.scala 216:26]
  wire  _GEN_329 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_93_data[32] ? 1'h0 : _GEN_279; // @[lut_35.scala 2827:105 lut_35.scala 216:26]
  wire  _GEN_332 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_93_data[32] ? 1'h0 : _GEN_282; // @[lut_35.scala 2827:105 lut_35.scala 216:26]
  wire  _GEN_335 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_93_data[32] ? 1'h0 : _GEN_285; // @[lut_35.scala 2827:105 lut_35.scala 216:26]
  wire  _GEN_338 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_93_data[32] ? 1'h0 : _GEN_288; // @[lut_35.scala 2827:105 lut_35.scala 216:26]
  wire [5:0] _GEN_339 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_92_data[32] ? 6'h16 : _GEN_289; // @[lut_35.scala 2785:105 lut_35.scala 2786:42]
  wire [31:0] _GEN_340 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_92_data[32] ? push_ray_id : _GEN_290; // @[lut_35.scala 2785:105 lut_35.scala 2787:42]
  wire  _GEN_343 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_92_data[32] ? 1'h0 : _T_442; // @[lut_35.scala 2785:105 lut_35.scala 2813:43]
  wire  _GEN_344 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_92_data[32] ? 1'h0 : _GEN_293; // @[lut_35.scala 2785:105 lut_35.scala 2814:43]
  wire  _GEN_345 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_92_data[32] ? 1'h0 : _GEN_294; // @[lut_35.scala 2785:105 lut_35.scala 2815:43]
  wire  _GEN_346 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_92_data[32] ? 1'h0 : _GEN_295; // @[lut_35.scala 2785:105 lut_35.scala 2816:43]
  wire  _GEN_347 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_92_data[32] ? 1'h0 : _GEN_296; // @[lut_35.scala 2785:105 lut_35.scala 2817:43]
  wire  _GEN_348 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_92_data[32] ? 1'h0 : _GEN_297; // @[lut_35.scala 2785:105 lut_35.scala 2818:43]
  wire  _GEN_349 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_92_data[32] ? 1'h0 : _GEN_298; // @[lut_35.scala 2785:105 lut_35.scala 2819:43]
  wire  _GEN_350 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_92_data[32] ? 1'h0 : _GEN_299; // @[lut_35.scala 2785:105 lut_35.scala 2820:43]
  wire  _GEN_351 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_92_data[32] ? 1'h0 : _GEN_300; // @[lut_35.scala 2785:105 lut_35.scala 2821:43]
  wire  _GEN_352 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_92_data[32] ? 1'h0 : _GEN_301; // @[lut_35.scala 2785:105 lut_35.scala 2822:43]
  wire  _GEN_353 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_92_data[32] ? 1'h0 : _GEN_302; // @[lut_35.scala 2785:105 lut_35.scala 2823:43]
  wire  _GEN_354 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_92_data[32] ? 1'h0 : _GEN_303; // @[lut_35.scala 2785:105 lut_35.scala 2824:43]
  wire  _GEN_355 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_92_data[32] | _GEN_304; // @[lut_35.scala 2785:105 lut_35.scala 2825:38]
  wire  _GEN_359 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_92_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2785:105 lut_35.scala 216:26 lut_35.scala 2827:89]
  wire  _GEN_362 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_92_data[32] ? 1'h0 : _GEN_308; // @[lut_35.scala 2785:105 lut_35.scala 216:26]
  wire  _GEN_365 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_92_data[32] ? 1'h0 : _GEN_311; // @[lut_35.scala 2785:105 lut_35.scala 216:26]
  wire  _GEN_368 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_92_data[32] ? 1'h0 : _GEN_314; // @[lut_35.scala 2785:105 lut_35.scala 216:26]
  wire  _GEN_371 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_92_data[32] ? 1'h0 : _GEN_317; // @[lut_35.scala 2785:105 lut_35.scala 216:26]
  wire  _GEN_374 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_92_data[32] ? 1'h0 : _GEN_320; // @[lut_35.scala 2785:105 lut_35.scala 216:26]
  wire  _GEN_377 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_92_data[32] ? 1'h0 : _GEN_323; // @[lut_35.scala 2785:105 lut_35.scala 216:26]
  wire  _GEN_380 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_92_data[32] ? 1'h0 : _GEN_326; // @[lut_35.scala 2785:105 lut_35.scala 216:26]
  wire  _GEN_383 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_92_data[32] ? 1'h0 : _GEN_329; // @[lut_35.scala 2785:105 lut_35.scala 216:26]
  wire  _GEN_386 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_92_data[32] ? 1'h0 : _GEN_332; // @[lut_35.scala 2785:105 lut_35.scala 216:26]
  wire  _GEN_389 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_92_data[32] ? 1'h0 : _GEN_335; // @[lut_35.scala 2785:105 lut_35.scala 216:26]
  wire  _GEN_392 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_92_data[32] ? 1'h0 : _GEN_338; // @[lut_35.scala 2785:105 lut_35.scala 216:26]
  wire [5:0] _GEN_393 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_91_data[32] ? 6'h15 : _GEN_339; // @[lut_35.scala 2743:105 lut_35.scala 2744:42]
  wire [31:0] _GEN_394 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_91_data[32] ? push_ray_id : _GEN_340; // @[lut_35.scala 2743:105 lut_35.scala 2745:42]
  wire  _GEN_397 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_91_data[32] ? 1'h0 : _T_434; // @[lut_35.scala 2743:105 lut_35.scala 2770:43]
  wire  _GEN_398 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_91_data[32] ? 1'h0 : _GEN_343; // @[lut_35.scala 2743:105 lut_35.scala 2771:43]
  wire  _GEN_399 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_91_data[32] ? 1'h0 : _GEN_344; // @[lut_35.scala 2743:105 lut_35.scala 2772:43]
  wire  _GEN_400 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_91_data[32] ? 1'h0 : _GEN_345; // @[lut_35.scala 2743:105 lut_35.scala 2773:43]
  wire  _GEN_401 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_91_data[32] ? 1'h0 : _GEN_346; // @[lut_35.scala 2743:105 lut_35.scala 2774:43]
  wire  _GEN_402 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_91_data[32] ? 1'h0 : _GEN_347; // @[lut_35.scala 2743:105 lut_35.scala 2775:43]
  wire  _GEN_403 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_91_data[32] ? 1'h0 : _GEN_348; // @[lut_35.scala 2743:105 lut_35.scala 2776:43]
  wire  _GEN_404 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_91_data[32] ? 1'h0 : _GEN_349; // @[lut_35.scala 2743:105 lut_35.scala 2777:43]
  wire  _GEN_405 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_91_data[32] ? 1'h0 : _GEN_350; // @[lut_35.scala 2743:105 lut_35.scala 2778:43]
  wire  _GEN_406 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_91_data[32] ? 1'h0 : _GEN_351; // @[lut_35.scala 2743:105 lut_35.scala 2779:43]
  wire  _GEN_407 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_91_data[32] ? 1'h0 : _GEN_352; // @[lut_35.scala 2743:105 lut_35.scala 2780:43]
  wire  _GEN_408 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_91_data[32] ? 1'h0 : _GEN_353; // @[lut_35.scala 2743:105 lut_35.scala 2781:43]
  wire  _GEN_409 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_91_data[32] ? 1'h0 : _GEN_354; // @[lut_35.scala 2743:105 lut_35.scala 2782:43]
  wire  _GEN_410 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_91_data[32] | _GEN_355; // @[lut_35.scala 2743:105 lut_35.scala 2783:38]
  wire  _GEN_414 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_91_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2743:105 lut_35.scala 216:26 lut_35.scala 2785:89]
  wire  _GEN_417 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_91_data[32] ? 1'h0 : _GEN_359; // @[lut_35.scala 2743:105 lut_35.scala 216:26]
  wire  _GEN_420 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_91_data[32] ? 1'h0 : _GEN_362; // @[lut_35.scala 2743:105 lut_35.scala 216:26]
  wire  _GEN_423 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_91_data[32] ? 1'h0 : _GEN_365; // @[lut_35.scala 2743:105 lut_35.scala 216:26]
  wire  _GEN_426 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_91_data[32] ? 1'h0 : _GEN_368; // @[lut_35.scala 2743:105 lut_35.scala 216:26]
  wire  _GEN_429 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_91_data[32] ? 1'h0 : _GEN_371; // @[lut_35.scala 2743:105 lut_35.scala 216:26]
  wire  _GEN_432 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_91_data[32] ? 1'h0 : _GEN_374; // @[lut_35.scala 2743:105 lut_35.scala 216:26]
  wire  _GEN_435 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_91_data[32] ? 1'h0 : _GEN_377; // @[lut_35.scala 2743:105 lut_35.scala 216:26]
  wire  _GEN_438 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_91_data[32] ? 1'h0 : _GEN_380; // @[lut_35.scala 2743:105 lut_35.scala 216:26]
  wire  _GEN_441 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_91_data[32] ? 1'h0 : _GEN_383; // @[lut_35.scala 2743:105 lut_35.scala 216:26]
  wire  _GEN_444 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_91_data[32] ? 1'h0 : _GEN_386; // @[lut_35.scala 2743:105 lut_35.scala 216:26]
  wire  _GEN_447 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_91_data[32] ? 1'h0 : _GEN_389; // @[lut_35.scala 2743:105 lut_35.scala 216:26]
  wire  _GEN_450 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_91_data[32] ? 1'h0 : _GEN_392; // @[lut_35.scala 2743:105 lut_35.scala 216:26]
  wire [5:0] _GEN_451 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_90_data[32] ? 6'h14 : _GEN_393; // @[lut_35.scala 2701:105 lut_35.scala 2702:42]
  wire [31:0] _GEN_452 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_90_data[32] ? push_ray_id : _GEN_394; // @[lut_35.scala 2701:105 lut_35.scala 2703:42]
  wire  _GEN_455 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_90_data[32] ? 1'h0 : _T_426; // @[lut_35.scala 2701:105 lut_35.scala 2727:43]
  wire  _GEN_456 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_90_data[32] ? 1'h0 : _GEN_397; // @[lut_35.scala 2701:105 lut_35.scala 2728:43]
  wire  _GEN_457 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_90_data[32] ? 1'h0 : _GEN_398; // @[lut_35.scala 2701:105 lut_35.scala 2729:43]
  wire  _GEN_458 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_90_data[32] ? 1'h0 : _GEN_399; // @[lut_35.scala 2701:105 lut_35.scala 2730:43]
  wire  _GEN_459 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_90_data[32] ? 1'h0 : _GEN_400; // @[lut_35.scala 2701:105 lut_35.scala 2731:43]
  wire  _GEN_460 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_90_data[32] ? 1'h0 : _GEN_401; // @[lut_35.scala 2701:105 lut_35.scala 2732:43]
  wire  _GEN_461 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_90_data[32] ? 1'h0 : _GEN_402; // @[lut_35.scala 2701:105 lut_35.scala 2733:43]
  wire  _GEN_462 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_90_data[32] ? 1'h0 : _GEN_403; // @[lut_35.scala 2701:105 lut_35.scala 2734:43]
  wire  _GEN_463 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_90_data[32] ? 1'h0 : _GEN_404; // @[lut_35.scala 2701:105 lut_35.scala 2735:43]
  wire  _GEN_464 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_90_data[32] ? 1'h0 : _GEN_405; // @[lut_35.scala 2701:105 lut_35.scala 2736:43]
  wire  _GEN_465 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_90_data[32] ? 1'h0 : _GEN_406; // @[lut_35.scala 2701:105 lut_35.scala 2737:43]
  wire  _GEN_466 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_90_data[32] ? 1'h0 : _GEN_407; // @[lut_35.scala 2701:105 lut_35.scala 2738:43]
  wire  _GEN_467 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_90_data[32] ? 1'h0 : _GEN_408; // @[lut_35.scala 2701:105 lut_35.scala 2739:43]
  wire  _GEN_468 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_90_data[32] ? 1'h0 : _GEN_409; // @[lut_35.scala 2701:105 lut_35.scala 2740:43]
  wire  _GEN_469 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_90_data[32] | _GEN_410; // @[lut_35.scala 2701:105 lut_35.scala 2741:38]
  wire  _GEN_473 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_90_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2701:105 lut_35.scala 216:26 lut_35.scala 2743:89]
  wire  _GEN_476 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_90_data[32] ? 1'h0 : _GEN_414; // @[lut_35.scala 2701:105 lut_35.scala 216:26]
  wire  _GEN_479 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_90_data[32] ? 1'h0 : _GEN_417; // @[lut_35.scala 2701:105 lut_35.scala 216:26]
  wire  _GEN_482 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_90_data[32] ? 1'h0 : _GEN_420; // @[lut_35.scala 2701:105 lut_35.scala 216:26]
  wire  _GEN_485 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_90_data[32] ? 1'h0 : _GEN_423; // @[lut_35.scala 2701:105 lut_35.scala 216:26]
  wire  _GEN_488 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_90_data[32] ? 1'h0 : _GEN_426; // @[lut_35.scala 2701:105 lut_35.scala 216:26]
  wire  _GEN_491 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_90_data[32] ? 1'h0 : _GEN_429; // @[lut_35.scala 2701:105 lut_35.scala 216:26]
  wire  _GEN_494 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_90_data[32] ? 1'h0 : _GEN_432; // @[lut_35.scala 2701:105 lut_35.scala 216:26]
  wire  _GEN_497 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_90_data[32] ? 1'h0 : _GEN_435; // @[lut_35.scala 2701:105 lut_35.scala 216:26]
  wire  _GEN_500 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_90_data[32] ? 1'h0 : _GEN_438; // @[lut_35.scala 2701:105 lut_35.scala 216:26]
  wire  _GEN_503 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_90_data[32] ? 1'h0 : _GEN_441; // @[lut_35.scala 2701:105 lut_35.scala 216:26]
  wire  _GEN_506 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_90_data[32] ? 1'h0 : _GEN_444; // @[lut_35.scala 2701:105 lut_35.scala 216:26]
  wire  _GEN_509 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_90_data[32] ? 1'h0 : _GEN_447; // @[lut_35.scala 2701:105 lut_35.scala 216:26]
  wire  _GEN_512 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_90_data[32] ? 1'h0 : _GEN_450; // @[lut_35.scala 2701:105 lut_35.scala 216:26]
  wire [5:0] _GEN_513 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_89_data[32] ? 6'h13 : _GEN_451; // @[lut_35.scala 2659:105 lut_35.scala 2660:42]
  wire [31:0] _GEN_514 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_89_data[32] ? push_ray_id : _GEN_452; // @[lut_35.scala 2659:105 lut_35.scala 2661:42]
  wire  _GEN_517 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_89_data[32] ? 1'h0 : _T_418; // @[lut_35.scala 2659:105 lut_35.scala 2684:43]
  wire  _GEN_518 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_89_data[32] ? 1'h0 : _GEN_455; // @[lut_35.scala 2659:105 lut_35.scala 2685:43]
  wire  _GEN_519 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_89_data[32] ? 1'h0 : _GEN_456; // @[lut_35.scala 2659:105 lut_35.scala 2686:43]
  wire  _GEN_520 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_89_data[32] ? 1'h0 : _GEN_457; // @[lut_35.scala 2659:105 lut_35.scala 2687:43]
  wire  _GEN_521 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_89_data[32] ? 1'h0 : _GEN_458; // @[lut_35.scala 2659:105 lut_35.scala 2688:43]
  wire  _GEN_522 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_89_data[32] ? 1'h0 : _GEN_459; // @[lut_35.scala 2659:105 lut_35.scala 2689:43]
  wire  _GEN_523 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_89_data[32] ? 1'h0 : _GEN_460; // @[lut_35.scala 2659:105 lut_35.scala 2690:43]
  wire  _GEN_524 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_89_data[32] ? 1'h0 : _GEN_461; // @[lut_35.scala 2659:105 lut_35.scala 2691:43]
  wire  _GEN_525 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_89_data[32] ? 1'h0 : _GEN_462; // @[lut_35.scala 2659:105 lut_35.scala 2692:43]
  wire  _GEN_526 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_89_data[32] ? 1'h0 : _GEN_463; // @[lut_35.scala 2659:105 lut_35.scala 2693:43]
  wire  _GEN_527 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_89_data[32] ? 1'h0 : _GEN_464; // @[lut_35.scala 2659:105 lut_35.scala 2694:43]
  wire  _GEN_528 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_89_data[32] ? 1'h0 : _GEN_465; // @[lut_35.scala 2659:105 lut_35.scala 2695:43]
  wire  _GEN_529 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_89_data[32] ? 1'h0 : _GEN_466; // @[lut_35.scala 2659:105 lut_35.scala 2696:43]
  wire  _GEN_530 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_89_data[32] ? 1'h0 : _GEN_467; // @[lut_35.scala 2659:105 lut_35.scala 2697:43]
  wire  _GEN_531 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_89_data[32] ? 1'h0 : _GEN_468; // @[lut_35.scala 2659:105 lut_35.scala 2698:43]
  wire  _GEN_532 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_89_data[32] | _GEN_469; // @[lut_35.scala 2659:105 lut_35.scala 2699:38]
  wire  _GEN_536 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_89_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2659:105 lut_35.scala 216:26 lut_35.scala 2701:89]
  wire  _GEN_539 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_89_data[32] ? 1'h0 : _GEN_473; // @[lut_35.scala 2659:105 lut_35.scala 216:26]
  wire  _GEN_542 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_89_data[32] ? 1'h0 : _GEN_476; // @[lut_35.scala 2659:105 lut_35.scala 216:26]
  wire  _GEN_545 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_89_data[32] ? 1'h0 : _GEN_479; // @[lut_35.scala 2659:105 lut_35.scala 216:26]
  wire  _GEN_548 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_89_data[32] ? 1'h0 : _GEN_482; // @[lut_35.scala 2659:105 lut_35.scala 216:26]
  wire  _GEN_551 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_89_data[32] ? 1'h0 : _GEN_485; // @[lut_35.scala 2659:105 lut_35.scala 216:26]
  wire  _GEN_554 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_89_data[32] ? 1'h0 : _GEN_488; // @[lut_35.scala 2659:105 lut_35.scala 216:26]
  wire  _GEN_557 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_89_data[32] ? 1'h0 : _GEN_491; // @[lut_35.scala 2659:105 lut_35.scala 216:26]
  wire  _GEN_560 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_89_data[32] ? 1'h0 : _GEN_494; // @[lut_35.scala 2659:105 lut_35.scala 216:26]
  wire  _GEN_563 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_89_data[32] ? 1'h0 : _GEN_497; // @[lut_35.scala 2659:105 lut_35.scala 216:26]
  wire  _GEN_566 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_89_data[32] ? 1'h0 : _GEN_500; // @[lut_35.scala 2659:105 lut_35.scala 216:26]
  wire  _GEN_569 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_89_data[32] ? 1'h0 : _GEN_503; // @[lut_35.scala 2659:105 lut_35.scala 216:26]
  wire  _GEN_572 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_89_data[32] ? 1'h0 : _GEN_506; // @[lut_35.scala 2659:105 lut_35.scala 216:26]
  wire  _GEN_575 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_89_data[32] ? 1'h0 : _GEN_509; // @[lut_35.scala 2659:105 lut_35.scala 216:26]
  wire  _GEN_578 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_89_data[32] ? 1'h0 : _GEN_512; // @[lut_35.scala 2659:105 lut_35.scala 216:26]
  wire [5:0] _GEN_579 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_88_data[32] ? 6'h12 : _GEN_513; // @[lut_35.scala 2617:105 lut_35.scala 2618:42]
  wire [31:0] _GEN_580 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_88_data[32] ? push_ray_id : _GEN_514; // @[lut_35.scala 2617:105 lut_35.scala 2619:42]
  wire  _GEN_583 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_88_data[32] ? 1'h0 : _T_410; // @[lut_35.scala 2617:105 lut_35.scala 2641:43]
  wire  _GEN_584 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_88_data[32] ? 1'h0 : _GEN_517; // @[lut_35.scala 2617:105 lut_35.scala 2642:43]
  wire  _GEN_585 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_88_data[32] ? 1'h0 : _GEN_518; // @[lut_35.scala 2617:105 lut_35.scala 2643:43]
  wire  _GEN_586 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_88_data[32] ? 1'h0 : _GEN_519; // @[lut_35.scala 2617:105 lut_35.scala 2644:43]
  wire  _GEN_587 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_88_data[32] ? 1'h0 : _GEN_520; // @[lut_35.scala 2617:105 lut_35.scala 2645:43]
  wire  _GEN_588 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_88_data[32] ? 1'h0 : _GEN_521; // @[lut_35.scala 2617:105 lut_35.scala 2646:43]
  wire  _GEN_589 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_88_data[32] ? 1'h0 : _GEN_522; // @[lut_35.scala 2617:105 lut_35.scala 2647:43]
  wire  _GEN_590 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_88_data[32] ? 1'h0 : _GEN_523; // @[lut_35.scala 2617:105 lut_35.scala 2648:43]
  wire  _GEN_591 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_88_data[32] ? 1'h0 : _GEN_524; // @[lut_35.scala 2617:105 lut_35.scala 2649:43]
  wire  _GEN_592 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_88_data[32] ? 1'h0 : _GEN_525; // @[lut_35.scala 2617:105 lut_35.scala 2650:43]
  wire  _GEN_593 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_88_data[32] ? 1'h0 : _GEN_526; // @[lut_35.scala 2617:105 lut_35.scala 2651:43]
  wire  _GEN_594 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_88_data[32] ? 1'h0 : _GEN_527; // @[lut_35.scala 2617:105 lut_35.scala 2652:43]
  wire  _GEN_595 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_88_data[32] ? 1'h0 : _GEN_528; // @[lut_35.scala 2617:105 lut_35.scala 2653:43]
  wire  _GEN_596 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_88_data[32] ? 1'h0 : _GEN_529; // @[lut_35.scala 2617:105 lut_35.scala 2654:43]
  wire  _GEN_597 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_88_data[32] ? 1'h0 : _GEN_530; // @[lut_35.scala 2617:105 lut_35.scala 2655:43]
  wire  _GEN_598 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_88_data[32] ? 1'h0 : _GEN_531; // @[lut_35.scala 2617:105 lut_35.scala 2656:43]
  wire  _GEN_599 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_88_data[32] | _GEN_532; // @[lut_35.scala 2617:105 lut_35.scala 2657:38]
  wire  _GEN_603 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_88_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2617:105 lut_35.scala 216:26 lut_35.scala 2659:89]
  wire  _GEN_606 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_88_data[32] ? 1'h0 : _GEN_536; // @[lut_35.scala 2617:105 lut_35.scala 216:26]
  wire  _GEN_609 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_88_data[32] ? 1'h0 : _GEN_539; // @[lut_35.scala 2617:105 lut_35.scala 216:26]
  wire  _GEN_612 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_88_data[32] ? 1'h0 : _GEN_542; // @[lut_35.scala 2617:105 lut_35.scala 216:26]
  wire  _GEN_615 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_88_data[32] ? 1'h0 : _GEN_545; // @[lut_35.scala 2617:105 lut_35.scala 216:26]
  wire  _GEN_618 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_88_data[32] ? 1'h0 : _GEN_548; // @[lut_35.scala 2617:105 lut_35.scala 216:26]
  wire  _GEN_621 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_88_data[32] ? 1'h0 : _GEN_551; // @[lut_35.scala 2617:105 lut_35.scala 216:26]
  wire  _GEN_624 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_88_data[32] ? 1'h0 : _GEN_554; // @[lut_35.scala 2617:105 lut_35.scala 216:26]
  wire  _GEN_627 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_88_data[32] ? 1'h0 : _GEN_557; // @[lut_35.scala 2617:105 lut_35.scala 216:26]
  wire  _GEN_630 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_88_data[32] ? 1'h0 : _GEN_560; // @[lut_35.scala 2617:105 lut_35.scala 216:26]
  wire  _GEN_633 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_88_data[32] ? 1'h0 : _GEN_563; // @[lut_35.scala 2617:105 lut_35.scala 216:26]
  wire  _GEN_636 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_88_data[32] ? 1'h0 : _GEN_566; // @[lut_35.scala 2617:105 lut_35.scala 216:26]
  wire  _GEN_639 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_88_data[32] ? 1'h0 : _GEN_569; // @[lut_35.scala 2617:105 lut_35.scala 216:26]
  wire  _GEN_642 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_88_data[32] ? 1'h0 : _GEN_572; // @[lut_35.scala 2617:105 lut_35.scala 216:26]
  wire  _GEN_645 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_88_data[32] ? 1'h0 : _GEN_575; // @[lut_35.scala 2617:105 lut_35.scala 216:26]
  wire  _GEN_648 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_88_data[32] ? 1'h0 : _GEN_578; // @[lut_35.scala 2617:105 lut_35.scala 216:26]
  wire [5:0] _GEN_649 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_87_data[32] ? 6'h11 : _GEN_579; // @[lut_35.scala 2575:105 lut_35.scala 2576:42]
  wire [31:0] _GEN_650 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_87_data[32] ? push_ray_id : _GEN_580; // @[lut_35.scala 2575:105 lut_35.scala 2577:42]
  wire  _GEN_653 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_87_data[32] ? 1'h0 : _T_402; // @[lut_35.scala 2575:105 lut_35.scala 2598:43]
  wire  _GEN_654 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_87_data[32] ? 1'h0 : _GEN_583; // @[lut_35.scala 2575:105 lut_35.scala 2599:43]
  wire  _GEN_655 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_87_data[32] ? 1'h0 : _GEN_584; // @[lut_35.scala 2575:105 lut_35.scala 2600:43]
  wire  _GEN_656 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_87_data[32] ? 1'h0 : _GEN_585; // @[lut_35.scala 2575:105 lut_35.scala 2601:43]
  wire  _GEN_657 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_87_data[32] ? 1'h0 : _GEN_586; // @[lut_35.scala 2575:105 lut_35.scala 2602:43]
  wire  _GEN_658 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_87_data[32] ? 1'h0 : _GEN_587; // @[lut_35.scala 2575:105 lut_35.scala 2603:43]
  wire  _GEN_659 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_87_data[32] ? 1'h0 : _GEN_588; // @[lut_35.scala 2575:105 lut_35.scala 2604:43]
  wire  _GEN_660 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_87_data[32] ? 1'h0 : _GEN_589; // @[lut_35.scala 2575:105 lut_35.scala 2605:43]
  wire  _GEN_661 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_87_data[32] ? 1'h0 : _GEN_590; // @[lut_35.scala 2575:105 lut_35.scala 2606:43]
  wire  _GEN_662 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_87_data[32] ? 1'h0 : _GEN_591; // @[lut_35.scala 2575:105 lut_35.scala 2607:43]
  wire  _GEN_663 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_87_data[32] ? 1'h0 : _GEN_592; // @[lut_35.scala 2575:105 lut_35.scala 2608:43]
  wire  _GEN_664 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_87_data[32] ? 1'h0 : _GEN_593; // @[lut_35.scala 2575:105 lut_35.scala 2609:43]
  wire  _GEN_665 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_87_data[32] ? 1'h0 : _GEN_594; // @[lut_35.scala 2575:105 lut_35.scala 2610:43]
  wire  _GEN_666 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_87_data[32] ? 1'h0 : _GEN_595; // @[lut_35.scala 2575:105 lut_35.scala 2611:43]
  wire  _GEN_667 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_87_data[32] ? 1'h0 : _GEN_596; // @[lut_35.scala 2575:105 lut_35.scala 2612:43]
  wire  _GEN_668 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_87_data[32] ? 1'h0 : _GEN_597; // @[lut_35.scala 2575:105 lut_35.scala 2613:43]
  wire  _GEN_669 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_87_data[32] ? 1'h0 : _GEN_598; // @[lut_35.scala 2575:105 lut_35.scala 2614:43]
  wire  _GEN_670 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_87_data[32] | _GEN_599; // @[lut_35.scala 2575:105 lut_35.scala 2615:38]
  wire  _GEN_674 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_87_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2575:105 lut_35.scala 216:26 lut_35.scala 2617:89]
  wire  _GEN_677 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_87_data[32] ? 1'h0 : _GEN_603; // @[lut_35.scala 2575:105 lut_35.scala 216:26]
  wire  _GEN_680 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_87_data[32] ? 1'h0 : _GEN_606; // @[lut_35.scala 2575:105 lut_35.scala 216:26]
  wire  _GEN_683 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_87_data[32] ? 1'h0 : _GEN_609; // @[lut_35.scala 2575:105 lut_35.scala 216:26]
  wire  _GEN_686 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_87_data[32] ? 1'h0 : _GEN_612; // @[lut_35.scala 2575:105 lut_35.scala 216:26]
  wire  _GEN_689 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_87_data[32] ? 1'h0 : _GEN_615; // @[lut_35.scala 2575:105 lut_35.scala 216:26]
  wire  _GEN_692 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_87_data[32] ? 1'h0 : _GEN_618; // @[lut_35.scala 2575:105 lut_35.scala 216:26]
  wire  _GEN_695 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_87_data[32] ? 1'h0 : _GEN_621; // @[lut_35.scala 2575:105 lut_35.scala 216:26]
  wire  _GEN_698 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_87_data[32] ? 1'h0 : _GEN_624; // @[lut_35.scala 2575:105 lut_35.scala 216:26]
  wire  _GEN_701 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_87_data[32] ? 1'h0 : _GEN_627; // @[lut_35.scala 2575:105 lut_35.scala 216:26]
  wire  _GEN_704 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_87_data[32] ? 1'h0 : _GEN_630; // @[lut_35.scala 2575:105 lut_35.scala 216:26]
  wire  _GEN_707 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_87_data[32] ? 1'h0 : _GEN_633; // @[lut_35.scala 2575:105 lut_35.scala 216:26]
  wire  _GEN_710 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_87_data[32] ? 1'h0 : _GEN_636; // @[lut_35.scala 2575:105 lut_35.scala 216:26]
  wire  _GEN_713 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_87_data[32] ? 1'h0 : _GEN_639; // @[lut_35.scala 2575:105 lut_35.scala 216:26]
  wire  _GEN_716 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_87_data[32] ? 1'h0 : _GEN_642; // @[lut_35.scala 2575:105 lut_35.scala 216:26]
  wire  _GEN_719 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_87_data[32] ? 1'h0 : _GEN_645; // @[lut_35.scala 2575:105 lut_35.scala 216:26]
  wire  _GEN_722 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_87_data[32] ? 1'h0 : _GEN_648; // @[lut_35.scala 2575:105 lut_35.scala 216:26]
  wire [5:0] _GEN_723 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_86_data[32] ? 6'h10 : _GEN_649; // @[lut_35.scala 2533:105 lut_35.scala 2534:42]
  wire [31:0] _GEN_724 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_86_data[32] ? push_ray_id : _GEN_650; // @[lut_35.scala 2533:105 lut_35.scala 2535:42]
  wire  _GEN_727 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_86_data[32] ? 1'h0 : _T_394; // @[lut_35.scala 2533:105 lut_35.scala 2555:43]
  wire  _GEN_728 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_86_data[32] ? 1'h0 : _GEN_653; // @[lut_35.scala 2533:105 lut_35.scala 2556:43]
  wire  _GEN_729 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_86_data[32] ? 1'h0 : _GEN_654; // @[lut_35.scala 2533:105 lut_35.scala 2557:43]
  wire  _GEN_730 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_86_data[32] ? 1'h0 : _GEN_655; // @[lut_35.scala 2533:105 lut_35.scala 2558:43]
  wire  _GEN_731 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_86_data[32] ? 1'h0 : _GEN_656; // @[lut_35.scala 2533:105 lut_35.scala 2559:43]
  wire  _GEN_732 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_86_data[32] ? 1'h0 : _GEN_657; // @[lut_35.scala 2533:105 lut_35.scala 2560:43]
  wire  _GEN_733 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_86_data[32] ? 1'h0 : _GEN_658; // @[lut_35.scala 2533:105 lut_35.scala 2561:43]
  wire  _GEN_734 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_86_data[32] ? 1'h0 : _GEN_659; // @[lut_35.scala 2533:105 lut_35.scala 2562:43]
  wire  _GEN_735 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_86_data[32] ? 1'h0 : _GEN_660; // @[lut_35.scala 2533:105 lut_35.scala 2563:43]
  wire  _GEN_736 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_86_data[32] ? 1'h0 : _GEN_661; // @[lut_35.scala 2533:105 lut_35.scala 2564:43]
  wire  _GEN_737 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_86_data[32] ? 1'h0 : _GEN_662; // @[lut_35.scala 2533:105 lut_35.scala 2565:43]
  wire  _GEN_738 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_86_data[32] ? 1'h0 : _GEN_663; // @[lut_35.scala 2533:105 lut_35.scala 2566:43]
  wire  _GEN_739 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_86_data[32] ? 1'h0 : _GEN_664; // @[lut_35.scala 2533:105 lut_35.scala 2567:43]
  wire  _GEN_740 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_86_data[32] ? 1'h0 : _GEN_665; // @[lut_35.scala 2533:105 lut_35.scala 2568:43]
  wire  _GEN_741 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_86_data[32] ? 1'h0 : _GEN_666; // @[lut_35.scala 2533:105 lut_35.scala 2569:43]
  wire  _GEN_742 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_86_data[32] ? 1'h0 : _GEN_667; // @[lut_35.scala 2533:105 lut_35.scala 2570:43]
  wire  _GEN_743 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_86_data[32] ? 1'h0 : _GEN_668; // @[lut_35.scala 2533:105 lut_35.scala 2571:43]
  wire  _GEN_744 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_86_data[32] ? 1'h0 : _GEN_669; // @[lut_35.scala 2533:105 lut_35.scala 2572:43]
  wire  _GEN_745 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_86_data[32] | _GEN_670; // @[lut_35.scala 2533:105 lut_35.scala 2573:38]
  wire  _GEN_749 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_86_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2533:105 lut_35.scala 216:26 lut_35.scala 2575:89]
  wire  _GEN_752 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_86_data[32] ? 1'h0 : _GEN_674; // @[lut_35.scala 2533:105 lut_35.scala 216:26]
  wire  _GEN_755 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_86_data[32] ? 1'h0 : _GEN_677; // @[lut_35.scala 2533:105 lut_35.scala 216:26]
  wire  _GEN_758 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_86_data[32] ? 1'h0 : _GEN_680; // @[lut_35.scala 2533:105 lut_35.scala 216:26]
  wire  _GEN_761 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_86_data[32] ? 1'h0 : _GEN_683; // @[lut_35.scala 2533:105 lut_35.scala 216:26]
  wire  _GEN_764 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_86_data[32] ? 1'h0 : _GEN_686; // @[lut_35.scala 2533:105 lut_35.scala 216:26]
  wire  _GEN_767 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_86_data[32] ? 1'h0 : _GEN_689; // @[lut_35.scala 2533:105 lut_35.scala 216:26]
  wire  _GEN_770 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_86_data[32] ? 1'h0 : _GEN_692; // @[lut_35.scala 2533:105 lut_35.scala 216:26]
  wire  _GEN_773 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_86_data[32] ? 1'h0 : _GEN_695; // @[lut_35.scala 2533:105 lut_35.scala 216:26]
  wire  _GEN_776 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_86_data[32] ? 1'h0 : _GEN_698; // @[lut_35.scala 2533:105 lut_35.scala 216:26]
  wire  _GEN_779 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_86_data[32] ? 1'h0 : _GEN_701; // @[lut_35.scala 2533:105 lut_35.scala 216:26]
  wire  _GEN_782 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_86_data[32] ? 1'h0 : _GEN_704; // @[lut_35.scala 2533:105 lut_35.scala 216:26]
  wire  _GEN_785 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_86_data[32] ? 1'h0 : _GEN_707; // @[lut_35.scala 2533:105 lut_35.scala 216:26]
  wire  _GEN_788 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_86_data[32] ? 1'h0 : _GEN_710; // @[lut_35.scala 2533:105 lut_35.scala 216:26]
  wire  _GEN_791 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_86_data[32] ? 1'h0 : _GEN_713; // @[lut_35.scala 2533:105 lut_35.scala 216:26]
  wire  _GEN_794 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_86_data[32] ? 1'h0 : _GEN_716; // @[lut_35.scala 2533:105 lut_35.scala 216:26]
  wire  _GEN_797 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_86_data[32] ? 1'h0 : _GEN_719; // @[lut_35.scala 2533:105 lut_35.scala 216:26]
  wire  _GEN_800 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_86_data[32] ? 1'h0 : _GEN_722; // @[lut_35.scala 2533:105 lut_35.scala 216:26]
  wire [5:0] _GEN_801 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_85_data[32] ? 6'hf : _GEN_723; // @[lut_35.scala 2491:105 lut_35.scala 2492:42]
  wire [31:0] _GEN_802 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_85_data[32] ? push_ray_id : _GEN_724; // @[lut_35.scala 2491:105 lut_35.scala 2493:42]
  wire  _GEN_805 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_85_data[32] ? 1'h0 : _T_386; // @[lut_35.scala 2491:105 lut_35.scala 2512:43]
  wire  _GEN_806 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_85_data[32] ? 1'h0 : _GEN_727; // @[lut_35.scala 2491:105 lut_35.scala 2513:43]
  wire  _GEN_807 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_85_data[32] ? 1'h0 : _GEN_728; // @[lut_35.scala 2491:105 lut_35.scala 2514:43]
  wire  _GEN_808 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_85_data[32] ? 1'h0 : _GEN_729; // @[lut_35.scala 2491:105 lut_35.scala 2515:43]
  wire  _GEN_809 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_85_data[32] ? 1'h0 : _GEN_730; // @[lut_35.scala 2491:105 lut_35.scala 2516:43]
  wire  _GEN_810 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_85_data[32] ? 1'h0 : _GEN_731; // @[lut_35.scala 2491:105 lut_35.scala 2517:43]
  wire  _GEN_811 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_85_data[32] ? 1'h0 : _GEN_732; // @[lut_35.scala 2491:105 lut_35.scala 2518:43]
  wire  _GEN_812 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_85_data[32] ? 1'h0 : _GEN_733; // @[lut_35.scala 2491:105 lut_35.scala 2519:43]
  wire  _GEN_813 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_85_data[32] ? 1'h0 : _GEN_734; // @[lut_35.scala 2491:105 lut_35.scala 2520:43]
  wire  _GEN_814 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_85_data[32] ? 1'h0 : _GEN_735; // @[lut_35.scala 2491:105 lut_35.scala 2521:43]
  wire  _GEN_815 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_85_data[32] ? 1'h0 : _GEN_736; // @[lut_35.scala 2491:105 lut_35.scala 2522:43]
  wire  _GEN_816 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_85_data[32] ? 1'h0 : _GEN_737; // @[lut_35.scala 2491:105 lut_35.scala 2523:43]
  wire  _GEN_817 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_85_data[32] ? 1'h0 : _GEN_738; // @[lut_35.scala 2491:105 lut_35.scala 2524:43]
  wire  _GEN_818 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_85_data[32] ? 1'h0 : _GEN_739; // @[lut_35.scala 2491:105 lut_35.scala 2525:43]
  wire  _GEN_819 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_85_data[32] ? 1'h0 : _GEN_740; // @[lut_35.scala 2491:105 lut_35.scala 2526:43]
  wire  _GEN_820 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_85_data[32] ? 1'h0 : _GEN_741; // @[lut_35.scala 2491:105 lut_35.scala 2527:43]
  wire  _GEN_821 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_85_data[32] ? 1'h0 : _GEN_742; // @[lut_35.scala 2491:105 lut_35.scala 2528:43]
  wire  _GEN_822 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_85_data[32] ? 1'h0 : _GEN_743; // @[lut_35.scala 2491:105 lut_35.scala 2529:43]
  wire  _GEN_823 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_85_data[32] ? 1'h0 : _GEN_744; // @[lut_35.scala 2491:105 lut_35.scala 2530:43]
  wire  _GEN_824 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_85_data[32] | _GEN_745; // @[lut_35.scala 2491:105 lut_35.scala 2531:38]
  wire  _GEN_828 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_85_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2491:105 lut_35.scala 216:26 lut_35.scala 2533:89]
  wire  _GEN_831 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_85_data[32] ? 1'h0 : _GEN_749; // @[lut_35.scala 2491:105 lut_35.scala 216:26]
  wire  _GEN_834 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_85_data[32] ? 1'h0 : _GEN_752; // @[lut_35.scala 2491:105 lut_35.scala 216:26]
  wire  _GEN_837 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_85_data[32] ? 1'h0 : _GEN_755; // @[lut_35.scala 2491:105 lut_35.scala 216:26]
  wire  _GEN_840 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_85_data[32] ? 1'h0 : _GEN_758; // @[lut_35.scala 2491:105 lut_35.scala 216:26]
  wire  _GEN_843 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_85_data[32] ? 1'h0 : _GEN_761; // @[lut_35.scala 2491:105 lut_35.scala 216:26]
  wire  _GEN_846 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_85_data[32] ? 1'h0 : _GEN_764; // @[lut_35.scala 2491:105 lut_35.scala 216:26]
  wire  _GEN_849 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_85_data[32] ? 1'h0 : _GEN_767; // @[lut_35.scala 2491:105 lut_35.scala 216:26]
  wire  _GEN_852 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_85_data[32] ? 1'h0 : _GEN_770; // @[lut_35.scala 2491:105 lut_35.scala 216:26]
  wire  _GEN_855 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_85_data[32] ? 1'h0 : _GEN_773; // @[lut_35.scala 2491:105 lut_35.scala 216:26]
  wire  _GEN_858 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_85_data[32] ? 1'h0 : _GEN_776; // @[lut_35.scala 2491:105 lut_35.scala 216:26]
  wire  _GEN_861 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_85_data[32] ? 1'h0 : _GEN_779; // @[lut_35.scala 2491:105 lut_35.scala 216:26]
  wire  _GEN_864 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_85_data[32] ? 1'h0 : _GEN_782; // @[lut_35.scala 2491:105 lut_35.scala 216:26]
  wire  _GEN_867 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_85_data[32] ? 1'h0 : _GEN_785; // @[lut_35.scala 2491:105 lut_35.scala 216:26]
  wire  _GEN_870 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_85_data[32] ? 1'h0 : _GEN_788; // @[lut_35.scala 2491:105 lut_35.scala 216:26]
  wire  _GEN_873 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_85_data[32] ? 1'h0 : _GEN_791; // @[lut_35.scala 2491:105 lut_35.scala 216:26]
  wire  _GEN_876 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_85_data[32] ? 1'h0 : _GEN_794; // @[lut_35.scala 2491:105 lut_35.scala 216:26]
  wire  _GEN_879 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_85_data[32] ? 1'h0 : _GEN_797; // @[lut_35.scala 2491:105 lut_35.scala 216:26]
  wire  _GEN_882 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_85_data[32] ? 1'h0 : _GEN_800; // @[lut_35.scala 2491:105 lut_35.scala 216:26]
  wire [5:0] _GEN_883 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] ? 6'he : _GEN_801; // @[lut_35.scala 2449:105 lut_35.scala 2450:42]
  wire [31:0] _GEN_884 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] ? push_ray_id : _GEN_802; // @[lut_35.scala 2449:105 lut_35.scala 2451:42]
  wire  _GEN_887 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] ? 1'h0 : _T_378; // @[lut_35.scala 2449:105 lut_35.scala 2469:43]
  wire  _GEN_888 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] ? 1'h0 : _GEN_805; // @[lut_35.scala 2449:105 lut_35.scala 2470:43]
  wire  _GEN_889 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] ? 1'h0 : _GEN_806; // @[lut_35.scala 2449:105 lut_35.scala 2471:43]
  wire  _GEN_890 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] ? 1'h0 : _GEN_807; // @[lut_35.scala 2449:105 lut_35.scala 2472:43]
  wire  _GEN_891 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] ? 1'h0 : _GEN_808; // @[lut_35.scala 2449:105 lut_35.scala 2473:43]
  wire  _GEN_892 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] ? 1'h0 : _GEN_809; // @[lut_35.scala 2449:105 lut_35.scala 2474:43]
  wire  _GEN_893 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] ? 1'h0 : _GEN_810; // @[lut_35.scala 2449:105 lut_35.scala 2475:43]
  wire  _GEN_894 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] ? 1'h0 : _GEN_811; // @[lut_35.scala 2449:105 lut_35.scala 2476:43]
  wire  _GEN_895 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] ? 1'h0 : _GEN_812; // @[lut_35.scala 2449:105 lut_35.scala 2477:43]
  wire  _GEN_896 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] ? 1'h0 : _GEN_813; // @[lut_35.scala 2449:105 lut_35.scala 2478:43]
  wire  _GEN_897 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] ? 1'h0 : _GEN_814; // @[lut_35.scala 2449:105 lut_35.scala 2479:43]
  wire  _GEN_898 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] ? 1'h0 : _GEN_815; // @[lut_35.scala 2449:105 lut_35.scala 2480:43]
  wire  _GEN_899 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] ? 1'h0 : _GEN_816; // @[lut_35.scala 2449:105 lut_35.scala 2481:43]
  wire  _GEN_900 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] ? 1'h0 : _GEN_817; // @[lut_35.scala 2449:105 lut_35.scala 2482:43]
  wire  _GEN_901 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] ? 1'h0 : _GEN_818; // @[lut_35.scala 2449:105 lut_35.scala 2483:43]
  wire  _GEN_902 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] ? 1'h0 : _GEN_819; // @[lut_35.scala 2449:105 lut_35.scala 2484:43]
  wire  _GEN_903 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] ? 1'h0 : _GEN_820; // @[lut_35.scala 2449:105 lut_35.scala 2485:43]
  wire  _GEN_904 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] ? 1'h0 : _GEN_821; // @[lut_35.scala 2449:105 lut_35.scala 2486:43]
  wire  _GEN_905 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] ? 1'h0 : _GEN_822; // @[lut_35.scala 2449:105 lut_35.scala 2487:43]
  wire  _GEN_906 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] ? 1'h0 : _GEN_823; // @[lut_35.scala 2449:105 lut_35.scala 2488:43]
  wire  _GEN_907 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] | _GEN_824; // @[lut_35.scala 2449:105 lut_35.scala 2489:38]
  wire  _GEN_911 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2449:105 lut_35.scala 216:26 lut_35.scala 2491:89]
  wire  _GEN_914 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] ? 1'h0 : _GEN_828; // @[lut_35.scala 2449:105 lut_35.scala 216:26]
  wire  _GEN_917 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] ? 1'h0 : _GEN_831; // @[lut_35.scala 2449:105 lut_35.scala 216:26]
  wire  _GEN_920 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] ? 1'h0 : _GEN_834; // @[lut_35.scala 2449:105 lut_35.scala 216:26]
  wire  _GEN_923 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] ? 1'h0 : _GEN_837; // @[lut_35.scala 2449:105 lut_35.scala 216:26]
  wire  _GEN_926 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] ? 1'h0 : _GEN_840; // @[lut_35.scala 2449:105 lut_35.scala 216:26]
  wire  _GEN_929 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] ? 1'h0 : _GEN_843; // @[lut_35.scala 2449:105 lut_35.scala 216:26]
  wire  _GEN_932 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] ? 1'h0 : _GEN_846; // @[lut_35.scala 2449:105 lut_35.scala 216:26]
  wire  _GEN_935 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] ? 1'h0 : _GEN_849; // @[lut_35.scala 2449:105 lut_35.scala 216:26]
  wire  _GEN_938 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] ? 1'h0 : _GEN_852; // @[lut_35.scala 2449:105 lut_35.scala 216:26]
  wire  _GEN_941 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] ? 1'h0 : _GEN_855; // @[lut_35.scala 2449:105 lut_35.scala 216:26]
  wire  _GEN_944 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] ? 1'h0 : _GEN_858; // @[lut_35.scala 2449:105 lut_35.scala 216:26]
  wire  _GEN_947 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] ? 1'h0 : _GEN_861; // @[lut_35.scala 2449:105 lut_35.scala 216:26]
  wire  _GEN_950 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] ? 1'h0 : _GEN_864; // @[lut_35.scala 2449:105 lut_35.scala 216:26]
  wire  _GEN_953 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] ? 1'h0 : _GEN_867; // @[lut_35.scala 2449:105 lut_35.scala 216:26]
  wire  _GEN_956 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] ? 1'h0 : _GEN_870; // @[lut_35.scala 2449:105 lut_35.scala 216:26]
  wire  _GEN_959 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] ? 1'h0 : _GEN_873; // @[lut_35.scala 2449:105 lut_35.scala 216:26]
  wire  _GEN_962 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] ? 1'h0 : _GEN_876; // @[lut_35.scala 2449:105 lut_35.scala 216:26]
  wire  _GEN_965 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] ? 1'h0 : _GEN_879; // @[lut_35.scala 2449:105 lut_35.scala 216:26]
  wire  _GEN_968 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_84_data[32] ? 1'h0 : _GEN_882; // @[lut_35.scala 2449:105 lut_35.scala 216:26]
  wire [5:0] _GEN_969 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 6'hd : _GEN_883; // @[lut_35.scala 2407:105 lut_35.scala 2408:42]
  wire [31:0] _GEN_970 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? push_ray_id : _GEN_884; // @[lut_35.scala 2407:105 lut_35.scala 2409:42]
  wire  _GEN_973 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 1'h0 : _T_370; // @[lut_35.scala 2407:105 lut_35.scala 2426:43]
  wire  _GEN_974 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 1'h0 : _GEN_887; // @[lut_35.scala 2407:105 lut_35.scala 2427:43]
  wire  _GEN_975 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 1'h0 : _GEN_888; // @[lut_35.scala 2407:105 lut_35.scala 2428:43]
  wire  _GEN_976 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 1'h0 : _GEN_889; // @[lut_35.scala 2407:105 lut_35.scala 2429:43]
  wire  _GEN_977 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 1'h0 : _GEN_890; // @[lut_35.scala 2407:105 lut_35.scala 2430:43]
  wire  _GEN_978 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 1'h0 : _GEN_891; // @[lut_35.scala 2407:105 lut_35.scala 2431:43]
  wire  _GEN_979 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 1'h0 : _GEN_892; // @[lut_35.scala 2407:105 lut_35.scala 2432:43]
  wire  _GEN_980 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 1'h0 : _GEN_893; // @[lut_35.scala 2407:105 lut_35.scala 2433:43]
  wire  _GEN_981 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 1'h0 : _GEN_894; // @[lut_35.scala 2407:105 lut_35.scala 2434:43]
  wire  _GEN_982 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 1'h0 : _GEN_895; // @[lut_35.scala 2407:105 lut_35.scala 2435:43]
  wire  _GEN_983 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 1'h0 : _GEN_896; // @[lut_35.scala 2407:105 lut_35.scala 2436:43]
  wire  _GEN_984 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 1'h0 : _GEN_897; // @[lut_35.scala 2407:105 lut_35.scala 2437:43]
  wire  _GEN_985 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 1'h0 : _GEN_898; // @[lut_35.scala 2407:105 lut_35.scala 2438:43]
  wire  _GEN_986 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 1'h0 : _GEN_899; // @[lut_35.scala 2407:105 lut_35.scala 2439:43]
  wire  _GEN_987 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 1'h0 : _GEN_900; // @[lut_35.scala 2407:105 lut_35.scala 2440:43]
  wire  _GEN_988 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 1'h0 : _GEN_901; // @[lut_35.scala 2407:105 lut_35.scala 2441:43]
  wire  _GEN_989 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 1'h0 : _GEN_902; // @[lut_35.scala 2407:105 lut_35.scala 2442:43]
  wire  _GEN_990 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 1'h0 : _GEN_903; // @[lut_35.scala 2407:105 lut_35.scala 2443:43]
  wire  _GEN_991 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 1'h0 : _GEN_904; // @[lut_35.scala 2407:105 lut_35.scala 2444:43]
  wire  _GEN_992 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 1'h0 : _GEN_905; // @[lut_35.scala 2407:105 lut_35.scala 2445:43]
  wire  _GEN_993 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 1'h0 : _GEN_906; // @[lut_35.scala 2407:105 lut_35.scala 2446:43]
  wire  _GEN_994 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] | _GEN_907; // @[lut_35.scala 2407:105 lut_35.scala 2447:38]
  wire  _GEN_998 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2407:105 lut_35.scala 216:26 lut_35.scala 2449:89]
  wire  _GEN_1001 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 1'h0 : _GEN_911; // @[lut_35.scala 2407:105 lut_35.scala 216:26]
  wire  _GEN_1004 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 1'h0 : _GEN_914; // @[lut_35.scala 2407:105 lut_35.scala 216:26]
  wire  _GEN_1007 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 1'h0 : _GEN_917; // @[lut_35.scala 2407:105 lut_35.scala 216:26]
  wire  _GEN_1010 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 1'h0 : _GEN_920; // @[lut_35.scala 2407:105 lut_35.scala 216:26]
  wire  _GEN_1013 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 1'h0 : _GEN_923; // @[lut_35.scala 2407:105 lut_35.scala 216:26]
  wire  _GEN_1016 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 1'h0 : _GEN_926; // @[lut_35.scala 2407:105 lut_35.scala 216:26]
  wire  _GEN_1019 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 1'h0 : _GEN_929; // @[lut_35.scala 2407:105 lut_35.scala 216:26]
  wire  _GEN_1022 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 1'h0 : _GEN_932; // @[lut_35.scala 2407:105 lut_35.scala 216:26]
  wire  _GEN_1025 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 1'h0 : _GEN_935; // @[lut_35.scala 2407:105 lut_35.scala 216:26]
  wire  _GEN_1028 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 1'h0 : _GEN_938; // @[lut_35.scala 2407:105 lut_35.scala 216:26]
  wire  _GEN_1031 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 1'h0 : _GEN_941; // @[lut_35.scala 2407:105 lut_35.scala 216:26]
  wire  _GEN_1034 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 1'h0 : _GEN_944; // @[lut_35.scala 2407:105 lut_35.scala 216:26]
  wire  _GEN_1037 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 1'h0 : _GEN_947; // @[lut_35.scala 2407:105 lut_35.scala 216:26]
  wire  _GEN_1040 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 1'h0 : _GEN_950; // @[lut_35.scala 2407:105 lut_35.scala 216:26]
  wire  _GEN_1043 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 1'h0 : _GEN_953; // @[lut_35.scala 2407:105 lut_35.scala 216:26]
  wire  _GEN_1046 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 1'h0 : _GEN_956; // @[lut_35.scala 2407:105 lut_35.scala 216:26]
  wire  _GEN_1049 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 1'h0 : _GEN_959; // @[lut_35.scala 2407:105 lut_35.scala 216:26]
  wire  _GEN_1052 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 1'h0 : _GEN_962; // @[lut_35.scala 2407:105 lut_35.scala 216:26]
  wire  _GEN_1055 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 1'h0 : _GEN_965; // @[lut_35.scala 2407:105 lut_35.scala 216:26]
  wire  _GEN_1058 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_83_data[32] ? 1'h0 : _GEN_968; // @[lut_35.scala 2407:105 lut_35.scala 216:26]
  wire [5:0] _GEN_1059 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 6'hc : _GEN_969; // @[lut_35.scala 2365:105 lut_35.scala 2366:42]
  wire [31:0] _GEN_1060 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? push_ray_id : _GEN_970; // @[lut_35.scala 2365:105 lut_35.scala 2367:42]
  wire  _GEN_1063 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _T_362; // @[lut_35.scala 2365:105 lut_35.scala 2383:43]
  wire  _GEN_1064 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _GEN_973; // @[lut_35.scala 2365:105 lut_35.scala 2384:43]
  wire  _GEN_1065 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _GEN_974; // @[lut_35.scala 2365:105 lut_35.scala 2385:43]
  wire  _GEN_1066 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _GEN_975; // @[lut_35.scala 2365:105 lut_35.scala 2386:43]
  wire  _GEN_1067 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _GEN_976; // @[lut_35.scala 2365:105 lut_35.scala 2387:43]
  wire  _GEN_1068 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _GEN_977; // @[lut_35.scala 2365:105 lut_35.scala 2388:43]
  wire  _GEN_1069 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _GEN_978; // @[lut_35.scala 2365:105 lut_35.scala 2389:43]
  wire  _GEN_1070 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _GEN_979; // @[lut_35.scala 2365:105 lut_35.scala 2390:43]
  wire  _GEN_1071 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _GEN_980; // @[lut_35.scala 2365:105 lut_35.scala 2391:43]
  wire  _GEN_1072 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _GEN_981; // @[lut_35.scala 2365:105 lut_35.scala 2392:43]
  wire  _GEN_1073 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _GEN_982; // @[lut_35.scala 2365:105 lut_35.scala 2393:43]
  wire  _GEN_1074 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _GEN_983; // @[lut_35.scala 2365:105 lut_35.scala 2394:43]
  wire  _GEN_1075 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _GEN_984; // @[lut_35.scala 2365:105 lut_35.scala 2395:43]
  wire  _GEN_1076 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _GEN_985; // @[lut_35.scala 2365:105 lut_35.scala 2396:43]
  wire  _GEN_1077 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _GEN_986; // @[lut_35.scala 2365:105 lut_35.scala 2397:43]
  wire  _GEN_1078 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _GEN_987; // @[lut_35.scala 2365:105 lut_35.scala 2398:43]
  wire  _GEN_1079 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _GEN_988; // @[lut_35.scala 2365:105 lut_35.scala 2399:43]
  wire  _GEN_1080 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _GEN_989; // @[lut_35.scala 2365:105 lut_35.scala 2400:43]
  wire  _GEN_1081 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _GEN_990; // @[lut_35.scala 2365:105 lut_35.scala 2401:43]
  wire  _GEN_1082 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _GEN_991; // @[lut_35.scala 2365:105 lut_35.scala 2402:43]
  wire  _GEN_1083 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _GEN_992; // @[lut_35.scala 2365:105 lut_35.scala 2403:43]
  wire  _GEN_1084 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _GEN_993; // @[lut_35.scala 2365:105 lut_35.scala 2404:43]
  wire  _GEN_1085 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] | _GEN_994; // @[lut_35.scala 2365:105 lut_35.scala 2405:38]
  wire  _GEN_1089 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2365:105 lut_35.scala 216:26 lut_35.scala 2407:89]
  wire  _GEN_1092 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _GEN_998; // @[lut_35.scala 2365:105 lut_35.scala 216:26]
  wire  _GEN_1095 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _GEN_1001; // @[lut_35.scala 2365:105 lut_35.scala 216:26]
  wire  _GEN_1098 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _GEN_1004; // @[lut_35.scala 2365:105 lut_35.scala 216:26]
  wire  _GEN_1101 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _GEN_1007; // @[lut_35.scala 2365:105 lut_35.scala 216:26]
  wire  _GEN_1104 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _GEN_1010; // @[lut_35.scala 2365:105 lut_35.scala 216:26]
  wire  _GEN_1107 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _GEN_1013; // @[lut_35.scala 2365:105 lut_35.scala 216:26]
  wire  _GEN_1110 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _GEN_1016; // @[lut_35.scala 2365:105 lut_35.scala 216:26]
  wire  _GEN_1113 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _GEN_1019; // @[lut_35.scala 2365:105 lut_35.scala 216:26]
  wire  _GEN_1116 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _GEN_1022; // @[lut_35.scala 2365:105 lut_35.scala 216:26]
  wire  _GEN_1119 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _GEN_1025; // @[lut_35.scala 2365:105 lut_35.scala 216:26]
  wire  _GEN_1122 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _GEN_1028; // @[lut_35.scala 2365:105 lut_35.scala 216:26]
  wire  _GEN_1125 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _GEN_1031; // @[lut_35.scala 2365:105 lut_35.scala 216:26]
  wire  _GEN_1128 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _GEN_1034; // @[lut_35.scala 2365:105 lut_35.scala 216:26]
  wire  _GEN_1131 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _GEN_1037; // @[lut_35.scala 2365:105 lut_35.scala 216:26]
  wire  _GEN_1134 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _GEN_1040; // @[lut_35.scala 2365:105 lut_35.scala 216:26]
  wire  _GEN_1137 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _GEN_1043; // @[lut_35.scala 2365:105 lut_35.scala 216:26]
  wire  _GEN_1140 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _GEN_1046; // @[lut_35.scala 2365:105 lut_35.scala 216:26]
  wire  _GEN_1143 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _GEN_1049; // @[lut_35.scala 2365:105 lut_35.scala 216:26]
  wire  _GEN_1146 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _GEN_1052; // @[lut_35.scala 2365:105 lut_35.scala 216:26]
  wire  _GEN_1149 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _GEN_1055; // @[lut_35.scala 2365:105 lut_35.scala 216:26]
  wire  _GEN_1152 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_82_data[32] ? 1'h0 : _GEN_1058; // @[lut_35.scala 2365:105 lut_35.scala 216:26]
  wire [5:0] _GEN_1153 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 6'hb : _GEN_1059; // @[lut_35.scala 2323:105 lut_35.scala 2324:42]
  wire [31:0] _GEN_1154 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? push_ray_id : _GEN_1060; // @[lut_35.scala 2323:105 lut_35.scala 2325:42]
  wire  _GEN_1157 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _T_354; // @[lut_35.scala 2323:105 lut_35.scala 2340:43]
  wire  _GEN_1158 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1063; // @[lut_35.scala 2323:105 lut_35.scala 2341:43]
  wire  _GEN_1159 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1064; // @[lut_35.scala 2323:105 lut_35.scala 2342:43]
  wire  _GEN_1160 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1065; // @[lut_35.scala 2323:105 lut_35.scala 2343:43]
  wire  _GEN_1161 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1066; // @[lut_35.scala 2323:105 lut_35.scala 2344:43]
  wire  _GEN_1162 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1067; // @[lut_35.scala 2323:105 lut_35.scala 2345:43]
  wire  _GEN_1163 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1068; // @[lut_35.scala 2323:105 lut_35.scala 2346:43]
  wire  _GEN_1164 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1069; // @[lut_35.scala 2323:105 lut_35.scala 2347:43]
  wire  _GEN_1165 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1070; // @[lut_35.scala 2323:105 lut_35.scala 2348:43]
  wire  _GEN_1166 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1071; // @[lut_35.scala 2323:105 lut_35.scala 2349:43]
  wire  _GEN_1167 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1072; // @[lut_35.scala 2323:105 lut_35.scala 2350:43]
  wire  _GEN_1168 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1073; // @[lut_35.scala 2323:105 lut_35.scala 2351:43]
  wire  _GEN_1169 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1074; // @[lut_35.scala 2323:105 lut_35.scala 2352:43]
  wire  _GEN_1170 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1075; // @[lut_35.scala 2323:105 lut_35.scala 2353:43]
  wire  _GEN_1171 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1076; // @[lut_35.scala 2323:105 lut_35.scala 2354:43]
  wire  _GEN_1172 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1077; // @[lut_35.scala 2323:105 lut_35.scala 2355:43]
  wire  _GEN_1173 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1078; // @[lut_35.scala 2323:105 lut_35.scala 2356:43]
  wire  _GEN_1174 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1079; // @[lut_35.scala 2323:105 lut_35.scala 2357:43]
  wire  _GEN_1175 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1080; // @[lut_35.scala 2323:105 lut_35.scala 2358:43]
  wire  _GEN_1176 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1081; // @[lut_35.scala 2323:105 lut_35.scala 2359:43]
  wire  _GEN_1177 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1082; // @[lut_35.scala 2323:105 lut_35.scala 2360:43]
  wire  _GEN_1178 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1083; // @[lut_35.scala 2323:105 lut_35.scala 2361:43]
  wire  _GEN_1179 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1084; // @[lut_35.scala 2323:105 lut_35.scala 2362:43]
  wire  _GEN_1180 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] | _GEN_1085; // @[lut_35.scala 2323:105 lut_35.scala 2363:38]
  wire  _GEN_1184 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2323:105 lut_35.scala 216:26 lut_35.scala 2365:89]
  wire  _GEN_1187 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1089; // @[lut_35.scala 2323:105 lut_35.scala 216:26]
  wire  _GEN_1190 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1092; // @[lut_35.scala 2323:105 lut_35.scala 216:26]
  wire  _GEN_1193 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1095; // @[lut_35.scala 2323:105 lut_35.scala 216:26]
  wire  _GEN_1196 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1098; // @[lut_35.scala 2323:105 lut_35.scala 216:26]
  wire  _GEN_1199 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1101; // @[lut_35.scala 2323:105 lut_35.scala 216:26]
  wire  _GEN_1202 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1104; // @[lut_35.scala 2323:105 lut_35.scala 216:26]
  wire  _GEN_1205 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1107; // @[lut_35.scala 2323:105 lut_35.scala 216:26]
  wire  _GEN_1208 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1110; // @[lut_35.scala 2323:105 lut_35.scala 216:26]
  wire  _GEN_1211 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1113; // @[lut_35.scala 2323:105 lut_35.scala 216:26]
  wire  _GEN_1214 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1116; // @[lut_35.scala 2323:105 lut_35.scala 216:26]
  wire  _GEN_1217 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1119; // @[lut_35.scala 2323:105 lut_35.scala 216:26]
  wire  _GEN_1220 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1122; // @[lut_35.scala 2323:105 lut_35.scala 216:26]
  wire  _GEN_1223 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1125; // @[lut_35.scala 2323:105 lut_35.scala 216:26]
  wire  _GEN_1226 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1128; // @[lut_35.scala 2323:105 lut_35.scala 216:26]
  wire  _GEN_1229 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1131; // @[lut_35.scala 2323:105 lut_35.scala 216:26]
  wire  _GEN_1232 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1134; // @[lut_35.scala 2323:105 lut_35.scala 216:26]
  wire  _GEN_1235 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1137; // @[lut_35.scala 2323:105 lut_35.scala 216:26]
  wire  _GEN_1238 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1140; // @[lut_35.scala 2323:105 lut_35.scala 216:26]
  wire  _GEN_1241 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1143; // @[lut_35.scala 2323:105 lut_35.scala 216:26]
  wire  _GEN_1244 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1146; // @[lut_35.scala 2323:105 lut_35.scala 216:26]
  wire  _GEN_1247 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1149; // @[lut_35.scala 2323:105 lut_35.scala 216:26]
  wire  _GEN_1250 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_81_data[32] ? 1'h0 : _GEN_1152; // @[lut_35.scala 2323:105 lut_35.scala 216:26]
  wire [5:0] _GEN_1251 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 6'ha : _GEN_1153; // @[lut_35.scala 2281:105 lut_35.scala 2282:42]
  wire [31:0] _GEN_1252 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? push_ray_id : _GEN_1154; // @[lut_35.scala 2281:105 lut_35.scala 2283:42]
  wire  _GEN_1255 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _T_346; // @[lut_35.scala 2281:105 lut_35.scala 2297:43]
  wire  _GEN_1256 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1157; // @[lut_35.scala 2281:105 lut_35.scala 2298:43]
  wire  _GEN_1257 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1158; // @[lut_35.scala 2281:105 lut_35.scala 2299:43]
  wire  _GEN_1258 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1159; // @[lut_35.scala 2281:105 lut_35.scala 2300:43]
  wire  _GEN_1259 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1160; // @[lut_35.scala 2281:105 lut_35.scala 2301:43]
  wire  _GEN_1260 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1161; // @[lut_35.scala 2281:105 lut_35.scala 2302:43]
  wire  _GEN_1261 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1162; // @[lut_35.scala 2281:105 lut_35.scala 2303:43]
  wire  _GEN_1262 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1163; // @[lut_35.scala 2281:105 lut_35.scala 2304:43]
  wire  _GEN_1263 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1164; // @[lut_35.scala 2281:105 lut_35.scala 2305:43]
  wire  _GEN_1264 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1165; // @[lut_35.scala 2281:105 lut_35.scala 2306:43]
  wire  _GEN_1265 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1166; // @[lut_35.scala 2281:105 lut_35.scala 2307:43]
  wire  _GEN_1266 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1167; // @[lut_35.scala 2281:105 lut_35.scala 2308:43]
  wire  _GEN_1267 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1168; // @[lut_35.scala 2281:105 lut_35.scala 2309:43]
  wire  _GEN_1268 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1169; // @[lut_35.scala 2281:105 lut_35.scala 2310:43]
  wire  _GEN_1269 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1170; // @[lut_35.scala 2281:105 lut_35.scala 2311:43]
  wire  _GEN_1270 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1171; // @[lut_35.scala 2281:105 lut_35.scala 2312:43]
  wire  _GEN_1271 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1172; // @[lut_35.scala 2281:105 lut_35.scala 2313:43]
  wire  _GEN_1272 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1173; // @[lut_35.scala 2281:105 lut_35.scala 2314:43]
  wire  _GEN_1273 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1174; // @[lut_35.scala 2281:105 lut_35.scala 2315:43]
  wire  _GEN_1274 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1175; // @[lut_35.scala 2281:105 lut_35.scala 2316:43]
  wire  _GEN_1275 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1176; // @[lut_35.scala 2281:105 lut_35.scala 2317:43]
  wire  _GEN_1276 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1177; // @[lut_35.scala 2281:105 lut_35.scala 2318:43]
  wire  _GEN_1277 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1178; // @[lut_35.scala 2281:105 lut_35.scala 2319:43]
  wire  _GEN_1278 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1179; // @[lut_35.scala 2281:105 lut_35.scala 2320:43]
  wire  _GEN_1279 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] | _GEN_1180; // @[lut_35.scala 2281:105 lut_35.scala 2321:38]
  wire  _GEN_1283 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2281:105 lut_35.scala 216:26 lut_35.scala 2323:89]
  wire  _GEN_1286 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1184; // @[lut_35.scala 2281:105 lut_35.scala 216:26]
  wire  _GEN_1289 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1187; // @[lut_35.scala 2281:105 lut_35.scala 216:26]
  wire  _GEN_1292 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1190; // @[lut_35.scala 2281:105 lut_35.scala 216:26]
  wire  _GEN_1295 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1193; // @[lut_35.scala 2281:105 lut_35.scala 216:26]
  wire  _GEN_1298 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1196; // @[lut_35.scala 2281:105 lut_35.scala 216:26]
  wire  _GEN_1301 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1199; // @[lut_35.scala 2281:105 lut_35.scala 216:26]
  wire  _GEN_1304 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1202; // @[lut_35.scala 2281:105 lut_35.scala 216:26]
  wire  _GEN_1307 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1205; // @[lut_35.scala 2281:105 lut_35.scala 216:26]
  wire  _GEN_1310 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1208; // @[lut_35.scala 2281:105 lut_35.scala 216:26]
  wire  _GEN_1313 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1211; // @[lut_35.scala 2281:105 lut_35.scala 216:26]
  wire  _GEN_1316 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1214; // @[lut_35.scala 2281:105 lut_35.scala 216:26]
  wire  _GEN_1319 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1217; // @[lut_35.scala 2281:105 lut_35.scala 216:26]
  wire  _GEN_1322 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1220; // @[lut_35.scala 2281:105 lut_35.scala 216:26]
  wire  _GEN_1325 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1223; // @[lut_35.scala 2281:105 lut_35.scala 216:26]
  wire  _GEN_1328 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1226; // @[lut_35.scala 2281:105 lut_35.scala 216:26]
  wire  _GEN_1331 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1229; // @[lut_35.scala 2281:105 lut_35.scala 216:26]
  wire  _GEN_1334 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1232; // @[lut_35.scala 2281:105 lut_35.scala 216:26]
  wire  _GEN_1337 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1235; // @[lut_35.scala 2281:105 lut_35.scala 216:26]
  wire  _GEN_1340 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1238; // @[lut_35.scala 2281:105 lut_35.scala 216:26]
  wire  _GEN_1343 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1241; // @[lut_35.scala 2281:105 lut_35.scala 216:26]
  wire  _GEN_1346 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1244; // @[lut_35.scala 2281:105 lut_35.scala 216:26]
  wire  _GEN_1349 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1247; // @[lut_35.scala 2281:105 lut_35.scala 216:26]
  wire  _GEN_1352 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_80_data[32] ? 1'h0 : _GEN_1250; // @[lut_35.scala 2281:105 lut_35.scala 216:26]
  wire [5:0] _GEN_1353 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 6'h9 : _GEN_1251; // @[lut_35.scala 2239:102 lut_35.scala 2240:42]
  wire [31:0] _GEN_1354 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? push_ray_id : _GEN_1252; // @[lut_35.scala 2239:102 lut_35.scala 2241:42]
  wire  _GEN_1357 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _T_338; // @[lut_35.scala 2239:102 lut_35.scala 2254:43]
  wire  _GEN_1358 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1255; // @[lut_35.scala 2239:102 lut_35.scala 2255:43]
  wire  _GEN_1359 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1256; // @[lut_35.scala 2239:102 lut_35.scala 2256:43]
  wire  _GEN_1360 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1257; // @[lut_35.scala 2239:102 lut_35.scala 2257:43]
  wire  _GEN_1361 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1258; // @[lut_35.scala 2239:102 lut_35.scala 2258:43]
  wire  _GEN_1362 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1259; // @[lut_35.scala 2239:102 lut_35.scala 2259:43]
  wire  _GEN_1363 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1260; // @[lut_35.scala 2239:102 lut_35.scala 2260:43]
  wire  _GEN_1364 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1261; // @[lut_35.scala 2239:102 lut_35.scala 2261:43]
  wire  _GEN_1365 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1262; // @[lut_35.scala 2239:102 lut_35.scala 2262:43]
  wire  _GEN_1366 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1263; // @[lut_35.scala 2239:102 lut_35.scala 2263:43]
  wire  _GEN_1367 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1264; // @[lut_35.scala 2239:102 lut_35.scala 2264:43]
  wire  _GEN_1368 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1265; // @[lut_35.scala 2239:102 lut_35.scala 2265:43]
  wire  _GEN_1369 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1266; // @[lut_35.scala 2239:102 lut_35.scala 2266:43]
  wire  _GEN_1370 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1267; // @[lut_35.scala 2239:102 lut_35.scala 2267:43]
  wire  _GEN_1371 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1268; // @[lut_35.scala 2239:102 lut_35.scala 2268:43]
  wire  _GEN_1372 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1269; // @[lut_35.scala 2239:102 lut_35.scala 2269:43]
  wire  _GEN_1373 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1270; // @[lut_35.scala 2239:102 lut_35.scala 2270:43]
  wire  _GEN_1374 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1271; // @[lut_35.scala 2239:102 lut_35.scala 2271:43]
  wire  _GEN_1375 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1272; // @[lut_35.scala 2239:102 lut_35.scala 2272:43]
  wire  _GEN_1376 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1273; // @[lut_35.scala 2239:102 lut_35.scala 2273:43]
  wire  _GEN_1377 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1274; // @[lut_35.scala 2239:102 lut_35.scala 2274:43]
  wire  _GEN_1378 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1275; // @[lut_35.scala 2239:102 lut_35.scala 2275:43]
  wire  _GEN_1379 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1276; // @[lut_35.scala 2239:102 lut_35.scala 2276:43]
  wire  _GEN_1380 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1277; // @[lut_35.scala 2239:102 lut_35.scala 2277:43]
  wire  _GEN_1381 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1278; // @[lut_35.scala 2239:102 lut_35.scala 2278:43]
  wire  _GEN_1382 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] | _GEN_1279; // @[lut_35.scala 2239:102 lut_35.scala 2279:38]
  wire  _GEN_1386 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2239:102 lut_35.scala 216:26 lut_35.scala 2281:89]
  wire  _GEN_1389 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1283; // @[lut_35.scala 2239:102 lut_35.scala 216:26]
  wire  _GEN_1392 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1286; // @[lut_35.scala 2239:102 lut_35.scala 216:26]
  wire  _GEN_1395 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1289; // @[lut_35.scala 2239:102 lut_35.scala 216:26]
  wire  _GEN_1398 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1292; // @[lut_35.scala 2239:102 lut_35.scala 216:26]
  wire  _GEN_1401 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1295; // @[lut_35.scala 2239:102 lut_35.scala 216:26]
  wire  _GEN_1404 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1298; // @[lut_35.scala 2239:102 lut_35.scala 216:26]
  wire  _GEN_1407 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1301; // @[lut_35.scala 2239:102 lut_35.scala 216:26]
  wire  _GEN_1410 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1304; // @[lut_35.scala 2239:102 lut_35.scala 216:26]
  wire  _GEN_1413 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1307; // @[lut_35.scala 2239:102 lut_35.scala 216:26]
  wire  _GEN_1416 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1310; // @[lut_35.scala 2239:102 lut_35.scala 216:26]
  wire  _GEN_1419 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1313; // @[lut_35.scala 2239:102 lut_35.scala 216:26]
  wire  _GEN_1422 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1316; // @[lut_35.scala 2239:102 lut_35.scala 216:26]
  wire  _GEN_1425 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1319; // @[lut_35.scala 2239:102 lut_35.scala 216:26]
  wire  _GEN_1428 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1322; // @[lut_35.scala 2239:102 lut_35.scala 216:26]
  wire  _GEN_1431 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1325; // @[lut_35.scala 2239:102 lut_35.scala 216:26]
  wire  _GEN_1434 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1328; // @[lut_35.scala 2239:102 lut_35.scala 216:26]
  wire  _GEN_1437 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1331; // @[lut_35.scala 2239:102 lut_35.scala 216:26]
  wire  _GEN_1440 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1334; // @[lut_35.scala 2239:102 lut_35.scala 216:26]
  wire  _GEN_1443 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1337; // @[lut_35.scala 2239:102 lut_35.scala 216:26]
  wire  _GEN_1446 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1340; // @[lut_35.scala 2239:102 lut_35.scala 216:26]
  wire  _GEN_1449 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1343; // @[lut_35.scala 2239:102 lut_35.scala 216:26]
  wire  _GEN_1452 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1346; // @[lut_35.scala 2239:102 lut_35.scala 216:26]
  wire  _GEN_1455 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1349; // @[lut_35.scala 2239:102 lut_35.scala 216:26]
  wire  _GEN_1458 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_79_data[32] ? 1'h0 : _GEN_1352; // @[lut_35.scala 2239:102 lut_35.scala 216:26]
  wire [5:0] _GEN_1459 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 6'h8 : _GEN_1353; // @[lut_35.scala 2197:102 lut_35.scala 2198:42]
  wire [31:0] _GEN_1460 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? push_ray_id : _GEN_1354; // @[lut_35.scala 2197:102 lut_35.scala 2199:42]
  wire  _GEN_1463 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _T_330; // @[lut_35.scala 2197:102 lut_35.scala 2211:42]
  wire  _GEN_1464 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1357; // @[lut_35.scala 2197:102 lut_35.scala 2212:43]
  wire  _GEN_1465 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1358; // @[lut_35.scala 2197:102 lut_35.scala 2213:43]
  wire  _GEN_1466 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1359; // @[lut_35.scala 2197:102 lut_35.scala 2214:43]
  wire  _GEN_1467 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1360; // @[lut_35.scala 2197:102 lut_35.scala 2215:43]
  wire  _GEN_1468 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1361; // @[lut_35.scala 2197:102 lut_35.scala 2216:43]
  wire  _GEN_1469 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1362; // @[lut_35.scala 2197:102 lut_35.scala 2217:43]
  wire  _GEN_1470 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1363; // @[lut_35.scala 2197:102 lut_35.scala 2218:43]
  wire  _GEN_1471 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1364; // @[lut_35.scala 2197:102 lut_35.scala 2219:43]
  wire  _GEN_1472 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1365; // @[lut_35.scala 2197:102 lut_35.scala 2220:43]
  wire  _GEN_1473 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1366; // @[lut_35.scala 2197:102 lut_35.scala 2221:43]
  wire  _GEN_1474 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1367; // @[lut_35.scala 2197:102 lut_35.scala 2222:43]
  wire  _GEN_1475 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1368; // @[lut_35.scala 2197:102 lut_35.scala 2223:43]
  wire  _GEN_1476 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1369; // @[lut_35.scala 2197:102 lut_35.scala 2224:43]
  wire  _GEN_1477 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1370; // @[lut_35.scala 2197:102 lut_35.scala 2225:43]
  wire  _GEN_1478 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1371; // @[lut_35.scala 2197:102 lut_35.scala 2226:43]
  wire  _GEN_1479 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1372; // @[lut_35.scala 2197:102 lut_35.scala 2227:43]
  wire  _GEN_1480 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1373; // @[lut_35.scala 2197:102 lut_35.scala 2228:43]
  wire  _GEN_1481 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1374; // @[lut_35.scala 2197:102 lut_35.scala 2229:43]
  wire  _GEN_1482 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1375; // @[lut_35.scala 2197:102 lut_35.scala 2230:43]
  wire  _GEN_1483 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1376; // @[lut_35.scala 2197:102 lut_35.scala 2231:43]
  wire  _GEN_1484 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1377; // @[lut_35.scala 2197:102 lut_35.scala 2232:43]
  wire  _GEN_1485 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1378; // @[lut_35.scala 2197:102 lut_35.scala 2233:43]
  wire  _GEN_1486 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1379; // @[lut_35.scala 2197:102 lut_35.scala 2234:43]
  wire  _GEN_1487 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1380; // @[lut_35.scala 2197:102 lut_35.scala 2235:43]
  wire  _GEN_1488 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1381; // @[lut_35.scala 2197:102 lut_35.scala 2236:43]
  wire  _GEN_1489 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] | _GEN_1382; // @[lut_35.scala 2197:102 lut_35.scala 2237:38]
  wire  _GEN_1493 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2197:102 lut_35.scala 216:26 lut_35.scala 2239:87]
  wire  _GEN_1496 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1386; // @[lut_35.scala 2197:102 lut_35.scala 216:26]
  wire  _GEN_1499 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1389; // @[lut_35.scala 2197:102 lut_35.scala 216:26]
  wire  _GEN_1502 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1392; // @[lut_35.scala 2197:102 lut_35.scala 216:26]
  wire  _GEN_1505 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1395; // @[lut_35.scala 2197:102 lut_35.scala 216:26]
  wire  _GEN_1508 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1398; // @[lut_35.scala 2197:102 lut_35.scala 216:26]
  wire  _GEN_1511 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1401; // @[lut_35.scala 2197:102 lut_35.scala 216:26]
  wire  _GEN_1514 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1404; // @[lut_35.scala 2197:102 lut_35.scala 216:26]
  wire  _GEN_1517 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1407; // @[lut_35.scala 2197:102 lut_35.scala 216:26]
  wire  _GEN_1520 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1410; // @[lut_35.scala 2197:102 lut_35.scala 216:26]
  wire  _GEN_1523 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1413; // @[lut_35.scala 2197:102 lut_35.scala 216:26]
  wire  _GEN_1526 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1416; // @[lut_35.scala 2197:102 lut_35.scala 216:26]
  wire  _GEN_1529 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1419; // @[lut_35.scala 2197:102 lut_35.scala 216:26]
  wire  _GEN_1532 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1422; // @[lut_35.scala 2197:102 lut_35.scala 216:26]
  wire  _GEN_1535 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1425; // @[lut_35.scala 2197:102 lut_35.scala 216:26]
  wire  _GEN_1538 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1428; // @[lut_35.scala 2197:102 lut_35.scala 216:26]
  wire  _GEN_1541 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1431; // @[lut_35.scala 2197:102 lut_35.scala 216:26]
  wire  _GEN_1544 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1434; // @[lut_35.scala 2197:102 lut_35.scala 216:26]
  wire  _GEN_1547 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1437; // @[lut_35.scala 2197:102 lut_35.scala 216:26]
  wire  _GEN_1550 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1440; // @[lut_35.scala 2197:102 lut_35.scala 216:26]
  wire  _GEN_1553 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1443; // @[lut_35.scala 2197:102 lut_35.scala 216:26]
  wire  _GEN_1556 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1446; // @[lut_35.scala 2197:102 lut_35.scala 216:26]
  wire  _GEN_1559 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1449; // @[lut_35.scala 2197:102 lut_35.scala 216:26]
  wire  _GEN_1562 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1452; // @[lut_35.scala 2197:102 lut_35.scala 216:26]
  wire  _GEN_1565 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1455; // @[lut_35.scala 2197:102 lut_35.scala 216:26]
  wire  _GEN_1568 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_78_data[32] ? 1'h0 : _GEN_1458; // @[lut_35.scala 2197:102 lut_35.scala 216:26]
  wire [5:0] _GEN_1569 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 6'h7 : _GEN_1459; // @[lut_35.scala 2155:102 lut_35.scala 2156:42]
  wire [31:0] _GEN_1570 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? push_ray_id : _GEN_1460; // @[lut_35.scala 2155:102 lut_35.scala 2157:42]
  wire  _GEN_1573 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _T_322; // @[lut_35.scala 2155:102 lut_35.scala 2168:42]
  wire  _GEN_1574 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1463; // @[lut_35.scala 2155:102 lut_35.scala 2169:42]
  wire  _GEN_1575 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1464; // @[lut_35.scala 2155:102 lut_35.scala 2170:43]
  wire  _GEN_1576 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1465; // @[lut_35.scala 2155:102 lut_35.scala 2171:43]
  wire  _GEN_1577 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1466; // @[lut_35.scala 2155:102 lut_35.scala 2172:43]
  wire  _GEN_1578 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1467; // @[lut_35.scala 2155:102 lut_35.scala 2173:43]
  wire  _GEN_1579 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1468; // @[lut_35.scala 2155:102 lut_35.scala 2174:43]
  wire  _GEN_1580 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1469; // @[lut_35.scala 2155:102 lut_35.scala 2175:43]
  wire  _GEN_1581 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1470; // @[lut_35.scala 2155:102 lut_35.scala 2176:43]
  wire  _GEN_1582 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1471; // @[lut_35.scala 2155:102 lut_35.scala 2177:43]
  wire  _GEN_1583 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1472; // @[lut_35.scala 2155:102 lut_35.scala 2178:43]
  wire  _GEN_1584 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1473; // @[lut_35.scala 2155:102 lut_35.scala 2179:43]
  wire  _GEN_1585 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1474; // @[lut_35.scala 2155:102 lut_35.scala 2180:43]
  wire  _GEN_1586 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1475; // @[lut_35.scala 2155:102 lut_35.scala 2181:43]
  wire  _GEN_1587 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1476; // @[lut_35.scala 2155:102 lut_35.scala 2182:43]
  wire  _GEN_1588 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1477; // @[lut_35.scala 2155:102 lut_35.scala 2183:43]
  wire  _GEN_1589 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1478; // @[lut_35.scala 2155:102 lut_35.scala 2184:43]
  wire  _GEN_1590 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1479; // @[lut_35.scala 2155:102 lut_35.scala 2185:43]
  wire  _GEN_1591 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1480; // @[lut_35.scala 2155:102 lut_35.scala 2186:43]
  wire  _GEN_1592 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1481; // @[lut_35.scala 2155:102 lut_35.scala 2187:43]
  wire  _GEN_1593 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1482; // @[lut_35.scala 2155:102 lut_35.scala 2188:43]
  wire  _GEN_1594 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1483; // @[lut_35.scala 2155:102 lut_35.scala 2189:43]
  wire  _GEN_1595 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1484; // @[lut_35.scala 2155:102 lut_35.scala 2190:43]
  wire  _GEN_1596 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1485; // @[lut_35.scala 2155:102 lut_35.scala 2191:43]
  wire  _GEN_1597 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1486; // @[lut_35.scala 2155:102 lut_35.scala 2192:43]
  wire  _GEN_1598 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1487; // @[lut_35.scala 2155:102 lut_35.scala 2193:43]
  wire  _GEN_1599 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1488; // @[lut_35.scala 2155:102 lut_35.scala 2194:43]
  wire  _GEN_1600 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] | _GEN_1489; // @[lut_35.scala 2155:102 lut_35.scala 2195:38]
  wire  _GEN_1604 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2155:102 lut_35.scala 216:26 lut_35.scala 2197:87]
  wire  _GEN_1607 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1493; // @[lut_35.scala 2155:102 lut_35.scala 216:26]
  wire  _GEN_1610 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1496; // @[lut_35.scala 2155:102 lut_35.scala 216:26]
  wire  _GEN_1613 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1499; // @[lut_35.scala 2155:102 lut_35.scala 216:26]
  wire  _GEN_1616 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1502; // @[lut_35.scala 2155:102 lut_35.scala 216:26]
  wire  _GEN_1619 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1505; // @[lut_35.scala 2155:102 lut_35.scala 216:26]
  wire  _GEN_1622 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1508; // @[lut_35.scala 2155:102 lut_35.scala 216:26]
  wire  _GEN_1625 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1511; // @[lut_35.scala 2155:102 lut_35.scala 216:26]
  wire  _GEN_1628 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1514; // @[lut_35.scala 2155:102 lut_35.scala 216:26]
  wire  _GEN_1631 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1517; // @[lut_35.scala 2155:102 lut_35.scala 216:26]
  wire  _GEN_1634 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1520; // @[lut_35.scala 2155:102 lut_35.scala 216:26]
  wire  _GEN_1637 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1523; // @[lut_35.scala 2155:102 lut_35.scala 216:26]
  wire  _GEN_1640 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1526; // @[lut_35.scala 2155:102 lut_35.scala 216:26]
  wire  _GEN_1643 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1529; // @[lut_35.scala 2155:102 lut_35.scala 216:26]
  wire  _GEN_1646 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1532; // @[lut_35.scala 2155:102 lut_35.scala 216:26]
  wire  _GEN_1649 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1535; // @[lut_35.scala 2155:102 lut_35.scala 216:26]
  wire  _GEN_1652 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1538; // @[lut_35.scala 2155:102 lut_35.scala 216:26]
  wire  _GEN_1655 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1541; // @[lut_35.scala 2155:102 lut_35.scala 216:26]
  wire  _GEN_1658 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1544; // @[lut_35.scala 2155:102 lut_35.scala 216:26]
  wire  _GEN_1661 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1547; // @[lut_35.scala 2155:102 lut_35.scala 216:26]
  wire  _GEN_1664 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1550; // @[lut_35.scala 2155:102 lut_35.scala 216:26]
  wire  _GEN_1667 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1553; // @[lut_35.scala 2155:102 lut_35.scala 216:26]
  wire  _GEN_1670 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1556; // @[lut_35.scala 2155:102 lut_35.scala 216:26]
  wire  _GEN_1673 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1559; // @[lut_35.scala 2155:102 lut_35.scala 216:26]
  wire  _GEN_1676 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1562; // @[lut_35.scala 2155:102 lut_35.scala 216:26]
  wire  _GEN_1679 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1565; // @[lut_35.scala 2155:102 lut_35.scala 216:26]
  wire  _GEN_1682 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_77_data[32] ? 1'h0 : _GEN_1568; // @[lut_35.scala 2155:102 lut_35.scala 216:26]
  wire [5:0] _GEN_1683 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 6'h6 : _GEN_1569; // @[lut_35.scala 2113:102 lut_35.scala 2114:42]
  wire [31:0] _GEN_1684 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? push_ray_id : _GEN_1570; // @[lut_35.scala 2113:102 lut_35.scala 2115:42]
  wire  _GEN_1687 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _T_314; // @[lut_35.scala 2113:102 lut_35.scala 2125:42]
  wire  _GEN_1688 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1573; // @[lut_35.scala 2113:102 lut_35.scala 2126:42]
  wire  _GEN_1689 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1574; // @[lut_35.scala 2113:102 lut_35.scala 2127:42]
  wire  _GEN_1690 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1575; // @[lut_35.scala 2113:102 lut_35.scala 2128:43]
  wire  _GEN_1691 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1576; // @[lut_35.scala 2113:102 lut_35.scala 2129:43]
  wire  _GEN_1692 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1577; // @[lut_35.scala 2113:102 lut_35.scala 2130:43]
  wire  _GEN_1693 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1578; // @[lut_35.scala 2113:102 lut_35.scala 2131:43]
  wire  _GEN_1694 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1579; // @[lut_35.scala 2113:102 lut_35.scala 2132:43]
  wire  _GEN_1695 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1580; // @[lut_35.scala 2113:102 lut_35.scala 2133:43]
  wire  _GEN_1696 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1581; // @[lut_35.scala 2113:102 lut_35.scala 2134:43]
  wire  _GEN_1697 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1582; // @[lut_35.scala 2113:102 lut_35.scala 2135:43]
  wire  _GEN_1698 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1583; // @[lut_35.scala 2113:102 lut_35.scala 2136:43]
  wire  _GEN_1699 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1584; // @[lut_35.scala 2113:102 lut_35.scala 2137:43]
  wire  _GEN_1700 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1585; // @[lut_35.scala 2113:102 lut_35.scala 2138:43]
  wire  _GEN_1701 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1586; // @[lut_35.scala 2113:102 lut_35.scala 2139:43]
  wire  _GEN_1702 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1587; // @[lut_35.scala 2113:102 lut_35.scala 2140:43]
  wire  _GEN_1703 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1588; // @[lut_35.scala 2113:102 lut_35.scala 2141:43]
  wire  _GEN_1704 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1589; // @[lut_35.scala 2113:102 lut_35.scala 2142:43]
  wire  _GEN_1705 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1590; // @[lut_35.scala 2113:102 lut_35.scala 2143:43]
  wire  _GEN_1706 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1591; // @[lut_35.scala 2113:102 lut_35.scala 2144:43]
  wire  _GEN_1707 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1592; // @[lut_35.scala 2113:102 lut_35.scala 2145:43]
  wire  _GEN_1708 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1593; // @[lut_35.scala 2113:102 lut_35.scala 2146:43]
  wire  _GEN_1709 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1594; // @[lut_35.scala 2113:102 lut_35.scala 2147:43]
  wire  _GEN_1710 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1595; // @[lut_35.scala 2113:102 lut_35.scala 2148:43]
  wire  _GEN_1711 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1596; // @[lut_35.scala 2113:102 lut_35.scala 2149:43]
  wire  _GEN_1712 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1597; // @[lut_35.scala 2113:102 lut_35.scala 2150:43]
  wire  _GEN_1713 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1598; // @[lut_35.scala 2113:102 lut_35.scala 2151:43]
  wire  _GEN_1714 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1599; // @[lut_35.scala 2113:102 lut_35.scala 2152:43]
  wire  _GEN_1715 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] | _GEN_1600; // @[lut_35.scala 2113:102 lut_35.scala 2153:38]
  wire  _GEN_1719 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2113:102 lut_35.scala 216:26 lut_35.scala 2155:87]
  wire  _GEN_1722 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1604; // @[lut_35.scala 2113:102 lut_35.scala 216:26]
  wire  _GEN_1725 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1607; // @[lut_35.scala 2113:102 lut_35.scala 216:26]
  wire  _GEN_1728 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1610; // @[lut_35.scala 2113:102 lut_35.scala 216:26]
  wire  _GEN_1731 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1613; // @[lut_35.scala 2113:102 lut_35.scala 216:26]
  wire  _GEN_1734 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1616; // @[lut_35.scala 2113:102 lut_35.scala 216:26]
  wire  _GEN_1737 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1619; // @[lut_35.scala 2113:102 lut_35.scala 216:26]
  wire  _GEN_1740 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1622; // @[lut_35.scala 2113:102 lut_35.scala 216:26]
  wire  _GEN_1743 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1625; // @[lut_35.scala 2113:102 lut_35.scala 216:26]
  wire  _GEN_1746 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1628; // @[lut_35.scala 2113:102 lut_35.scala 216:26]
  wire  _GEN_1749 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1631; // @[lut_35.scala 2113:102 lut_35.scala 216:26]
  wire  _GEN_1752 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1634; // @[lut_35.scala 2113:102 lut_35.scala 216:26]
  wire  _GEN_1755 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1637; // @[lut_35.scala 2113:102 lut_35.scala 216:26]
  wire  _GEN_1758 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1640; // @[lut_35.scala 2113:102 lut_35.scala 216:26]
  wire  _GEN_1761 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1643; // @[lut_35.scala 2113:102 lut_35.scala 216:26]
  wire  _GEN_1764 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1646; // @[lut_35.scala 2113:102 lut_35.scala 216:26]
  wire  _GEN_1767 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1649; // @[lut_35.scala 2113:102 lut_35.scala 216:26]
  wire  _GEN_1770 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1652; // @[lut_35.scala 2113:102 lut_35.scala 216:26]
  wire  _GEN_1773 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1655; // @[lut_35.scala 2113:102 lut_35.scala 216:26]
  wire  _GEN_1776 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1658; // @[lut_35.scala 2113:102 lut_35.scala 216:26]
  wire  _GEN_1779 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1661; // @[lut_35.scala 2113:102 lut_35.scala 216:26]
  wire  _GEN_1782 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1664; // @[lut_35.scala 2113:102 lut_35.scala 216:26]
  wire  _GEN_1785 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1667; // @[lut_35.scala 2113:102 lut_35.scala 216:26]
  wire  _GEN_1788 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1670; // @[lut_35.scala 2113:102 lut_35.scala 216:26]
  wire  _GEN_1791 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1673; // @[lut_35.scala 2113:102 lut_35.scala 216:26]
  wire  _GEN_1794 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1676; // @[lut_35.scala 2113:102 lut_35.scala 216:26]
  wire  _GEN_1797 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1679; // @[lut_35.scala 2113:102 lut_35.scala 216:26]
  wire  _GEN_1800 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_76_data[32] ? 1'h0 : _GEN_1682; // @[lut_35.scala 2113:102 lut_35.scala 216:26]
  wire [5:0] _GEN_1801 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 6'h5 : _GEN_1683; // @[lut_35.scala 2071:102 lut_35.scala 2072:42]
  wire [31:0] _GEN_1802 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? push_ray_id : _GEN_1684; // @[lut_35.scala 2071:102 lut_35.scala 2073:42]
  wire  _GEN_1805 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _T_306; // @[lut_35.scala 2071:102 lut_35.scala 2082:42]
  wire  _GEN_1806 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1687; // @[lut_35.scala 2071:102 lut_35.scala 2083:42]
  wire  _GEN_1807 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1688; // @[lut_35.scala 2071:102 lut_35.scala 2084:42]
  wire  _GEN_1808 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1689; // @[lut_35.scala 2071:102 lut_35.scala 2085:42]
  wire  _GEN_1809 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1690; // @[lut_35.scala 2071:102 lut_35.scala 2086:43]
  wire  _GEN_1810 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1691; // @[lut_35.scala 2071:102 lut_35.scala 2087:43]
  wire  _GEN_1811 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1692; // @[lut_35.scala 2071:102 lut_35.scala 2088:43]
  wire  _GEN_1812 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1693; // @[lut_35.scala 2071:102 lut_35.scala 2089:43]
  wire  _GEN_1813 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1694; // @[lut_35.scala 2071:102 lut_35.scala 2090:43]
  wire  _GEN_1814 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1695; // @[lut_35.scala 2071:102 lut_35.scala 2091:43]
  wire  _GEN_1815 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1696; // @[lut_35.scala 2071:102 lut_35.scala 2092:43]
  wire  _GEN_1816 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1697; // @[lut_35.scala 2071:102 lut_35.scala 2093:43]
  wire  _GEN_1817 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1698; // @[lut_35.scala 2071:102 lut_35.scala 2094:43]
  wire  _GEN_1818 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1699; // @[lut_35.scala 2071:102 lut_35.scala 2095:43]
  wire  _GEN_1819 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1700; // @[lut_35.scala 2071:102 lut_35.scala 2096:43]
  wire  _GEN_1820 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1701; // @[lut_35.scala 2071:102 lut_35.scala 2097:43]
  wire  _GEN_1821 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1702; // @[lut_35.scala 2071:102 lut_35.scala 2098:43]
  wire  _GEN_1822 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1703; // @[lut_35.scala 2071:102 lut_35.scala 2099:43]
  wire  _GEN_1823 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1704; // @[lut_35.scala 2071:102 lut_35.scala 2100:43]
  wire  _GEN_1824 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1705; // @[lut_35.scala 2071:102 lut_35.scala 2101:43]
  wire  _GEN_1825 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1706; // @[lut_35.scala 2071:102 lut_35.scala 2102:43]
  wire  _GEN_1826 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1707; // @[lut_35.scala 2071:102 lut_35.scala 2103:43]
  wire  _GEN_1827 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1708; // @[lut_35.scala 2071:102 lut_35.scala 2104:43]
  wire  _GEN_1828 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1709; // @[lut_35.scala 2071:102 lut_35.scala 2105:43]
  wire  _GEN_1829 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1710; // @[lut_35.scala 2071:102 lut_35.scala 2106:43]
  wire  _GEN_1830 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1711; // @[lut_35.scala 2071:102 lut_35.scala 2107:43]
  wire  _GEN_1831 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1712; // @[lut_35.scala 2071:102 lut_35.scala 2108:43]
  wire  _GEN_1832 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1713; // @[lut_35.scala 2071:102 lut_35.scala 2109:43]
  wire  _GEN_1833 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1714; // @[lut_35.scala 2071:102 lut_35.scala 2110:43]
  wire  _GEN_1834 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] | _GEN_1715; // @[lut_35.scala 2071:102 lut_35.scala 2111:38]
  wire  _GEN_1838 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2071:102 lut_35.scala 216:26 lut_35.scala 2113:87]
  wire  _GEN_1841 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1719; // @[lut_35.scala 2071:102 lut_35.scala 216:26]
  wire  _GEN_1844 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1722; // @[lut_35.scala 2071:102 lut_35.scala 216:26]
  wire  _GEN_1847 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1725; // @[lut_35.scala 2071:102 lut_35.scala 216:26]
  wire  _GEN_1850 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1728; // @[lut_35.scala 2071:102 lut_35.scala 216:26]
  wire  _GEN_1853 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1731; // @[lut_35.scala 2071:102 lut_35.scala 216:26]
  wire  _GEN_1856 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1734; // @[lut_35.scala 2071:102 lut_35.scala 216:26]
  wire  _GEN_1859 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1737; // @[lut_35.scala 2071:102 lut_35.scala 216:26]
  wire  _GEN_1862 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1740; // @[lut_35.scala 2071:102 lut_35.scala 216:26]
  wire  _GEN_1865 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1743; // @[lut_35.scala 2071:102 lut_35.scala 216:26]
  wire  _GEN_1868 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1746; // @[lut_35.scala 2071:102 lut_35.scala 216:26]
  wire  _GEN_1871 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1749; // @[lut_35.scala 2071:102 lut_35.scala 216:26]
  wire  _GEN_1874 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1752; // @[lut_35.scala 2071:102 lut_35.scala 216:26]
  wire  _GEN_1877 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1755; // @[lut_35.scala 2071:102 lut_35.scala 216:26]
  wire  _GEN_1880 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1758; // @[lut_35.scala 2071:102 lut_35.scala 216:26]
  wire  _GEN_1883 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1761; // @[lut_35.scala 2071:102 lut_35.scala 216:26]
  wire  _GEN_1886 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1764; // @[lut_35.scala 2071:102 lut_35.scala 216:26]
  wire  _GEN_1889 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1767; // @[lut_35.scala 2071:102 lut_35.scala 216:26]
  wire  _GEN_1892 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1770; // @[lut_35.scala 2071:102 lut_35.scala 216:26]
  wire  _GEN_1895 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1773; // @[lut_35.scala 2071:102 lut_35.scala 216:26]
  wire  _GEN_1898 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1776; // @[lut_35.scala 2071:102 lut_35.scala 216:26]
  wire  _GEN_1901 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1779; // @[lut_35.scala 2071:102 lut_35.scala 216:26]
  wire  _GEN_1904 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1782; // @[lut_35.scala 2071:102 lut_35.scala 216:26]
  wire  _GEN_1907 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1785; // @[lut_35.scala 2071:102 lut_35.scala 216:26]
  wire  _GEN_1910 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1788; // @[lut_35.scala 2071:102 lut_35.scala 216:26]
  wire  _GEN_1913 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1791; // @[lut_35.scala 2071:102 lut_35.scala 216:26]
  wire  _GEN_1916 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1794; // @[lut_35.scala 2071:102 lut_35.scala 216:26]
  wire  _GEN_1919 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1797; // @[lut_35.scala 2071:102 lut_35.scala 216:26]
  wire  _GEN_1922 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_75_data[32] ? 1'h0 : _GEN_1800; // @[lut_35.scala 2071:102 lut_35.scala 216:26]
  wire [5:0] _GEN_1923 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 6'h4 : _GEN_1801; // @[lut_35.scala 2029:102 lut_35.scala 2030:42]
  wire [31:0] _GEN_1924 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? push_ray_id : _GEN_1802; // @[lut_35.scala 2029:102 lut_35.scala 2031:42]
  wire  _GEN_1927 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _T_298; // @[lut_35.scala 2029:102 lut_35.scala 2039:42]
  wire  _GEN_1928 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1805; // @[lut_35.scala 2029:102 lut_35.scala 2040:42]
  wire  _GEN_1929 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1806; // @[lut_35.scala 2029:102 lut_35.scala 2041:42]
  wire  _GEN_1930 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1807; // @[lut_35.scala 2029:102 lut_35.scala 2042:42]
  wire  _GEN_1931 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1808; // @[lut_35.scala 2029:102 lut_35.scala 2043:42]
  wire  _GEN_1932 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1809; // @[lut_35.scala 2029:102 lut_35.scala 2044:43]
  wire  _GEN_1933 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1810; // @[lut_35.scala 2029:102 lut_35.scala 2045:43]
  wire  _GEN_1934 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1811; // @[lut_35.scala 2029:102 lut_35.scala 2046:43]
  wire  _GEN_1935 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1812; // @[lut_35.scala 2029:102 lut_35.scala 2047:43]
  wire  _GEN_1936 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1813; // @[lut_35.scala 2029:102 lut_35.scala 2048:43]
  wire  _GEN_1937 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1814; // @[lut_35.scala 2029:102 lut_35.scala 2049:43]
  wire  _GEN_1938 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1815; // @[lut_35.scala 2029:102 lut_35.scala 2050:43]
  wire  _GEN_1939 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1816; // @[lut_35.scala 2029:102 lut_35.scala 2051:43]
  wire  _GEN_1940 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1817; // @[lut_35.scala 2029:102 lut_35.scala 2052:43]
  wire  _GEN_1941 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1818; // @[lut_35.scala 2029:102 lut_35.scala 2053:43]
  wire  _GEN_1942 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1819; // @[lut_35.scala 2029:102 lut_35.scala 2054:43]
  wire  _GEN_1943 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1820; // @[lut_35.scala 2029:102 lut_35.scala 2055:43]
  wire  _GEN_1944 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1821; // @[lut_35.scala 2029:102 lut_35.scala 2056:43]
  wire  _GEN_1945 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1822; // @[lut_35.scala 2029:102 lut_35.scala 2057:43]
  wire  _GEN_1946 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1823; // @[lut_35.scala 2029:102 lut_35.scala 2058:43]
  wire  _GEN_1947 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1824; // @[lut_35.scala 2029:102 lut_35.scala 2059:43]
  wire  _GEN_1948 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1825; // @[lut_35.scala 2029:102 lut_35.scala 2060:43]
  wire  _GEN_1949 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1826; // @[lut_35.scala 2029:102 lut_35.scala 2061:43]
  wire  _GEN_1950 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1827; // @[lut_35.scala 2029:102 lut_35.scala 2062:43]
  wire  _GEN_1951 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1828; // @[lut_35.scala 2029:102 lut_35.scala 2063:43]
  wire  _GEN_1952 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1829; // @[lut_35.scala 2029:102 lut_35.scala 2064:43]
  wire  _GEN_1953 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1830; // @[lut_35.scala 2029:102 lut_35.scala 2065:43]
  wire  _GEN_1954 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1831; // @[lut_35.scala 2029:102 lut_35.scala 2066:43]
  wire  _GEN_1955 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1832; // @[lut_35.scala 2029:102 lut_35.scala 2067:43]
  wire  _GEN_1956 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1833; // @[lut_35.scala 2029:102 lut_35.scala 2068:43]
  wire  _GEN_1957 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] | _GEN_1834; // @[lut_35.scala 2029:102 lut_35.scala 2069:38]
  wire  _GEN_1961 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2029:102 lut_35.scala 216:26 lut_35.scala 2071:87]
  wire  _GEN_1964 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1838; // @[lut_35.scala 2029:102 lut_35.scala 216:26]
  wire  _GEN_1967 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1841; // @[lut_35.scala 2029:102 lut_35.scala 216:26]
  wire  _GEN_1970 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1844; // @[lut_35.scala 2029:102 lut_35.scala 216:26]
  wire  _GEN_1973 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1847; // @[lut_35.scala 2029:102 lut_35.scala 216:26]
  wire  _GEN_1976 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1850; // @[lut_35.scala 2029:102 lut_35.scala 216:26]
  wire  _GEN_1979 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1853; // @[lut_35.scala 2029:102 lut_35.scala 216:26]
  wire  _GEN_1982 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1856; // @[lut_35.scala 2029:102 lut_35.scala 216:26]
  wire  _GEN_1985 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1859; // @[lut_35.scala 2029:102 lut_35.scala 216:26]
  wire  _GEN_1988 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1862; // @[lut_35.scala 2029:102 lut_35.scala 216:26]
  wire  _GEN_1991 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1865; // @[lut_35.scala 2029:102 lut_35.scala 216:26]
  wire  _GEN_1994 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1868; // @[lut_35.scala 2029:102 lut_35.scala 216:26]
  wire  _GEN_1997 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1871; // @[lut_35.scala 2029:102 lut_35.scala 216:26]
  wire  _GEN_2000 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1874; // @[lut_35.scala 2029:102 lut_35.scala 216:26]
  wire  _GEN_2003 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1877; // @[lut_35.scala 2029:102 lut_35.scala 216:26]
  wire  _GEN_2006 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1880; // @[lut_35.scala 2029:102 lut_35.scala 216:26]
  wire  _GEN_2009 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1883; // @[lut_35.scala 2029:102 lut_35.scala 216:26]
  wire  _GEN_2012 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1886; // @[lut_35.scala 2029:102 lut_35.scala 216:26]
  wire  _GEN_2015 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1889; // @[lut_35.scala 2029:102 lut_35.scala 216:26]
  wire  _GEN_2018 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1892; // @[lut_35.scala 2029:102 lut_35.scala 216:26]
  wire  _GEN_2021 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1895; // @[lut_35.scala 2029:102 lut_35.scala 216:26]
  wire  _GEN_2024 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1898; // @[lut_35.scala 2029:102 lut_35.scala 216:26]
  wire  _GEN_2027 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1901; // @[lut_35.scala 2029:102 lut_35.scala 216:26]
  wire  _GEN_2030 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1904; // @[lut_35.scala 2029:102 lut_35.scala 216:26]
  wire  _GEN_2033 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1907; // @[lut_35.scala 2029:102 lut_35.scala 216:26]
  wire  _GEN_2036 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1910; // @[lut_35.scala 2029:102 lut_35.scala 216:26]
  wire  _GEN_2039 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1913; // @[lut_35.scala 2029:102 lut_35.scala 216:26]
  wire  _GEN_2042 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1916; // @[lut_35.scala 2029:102 lut_35.scala 216:26]
  wire  _GEN_2045 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1919; // @[lut_35.scala 2029:102 lut_35.scala 216:26]
  wire  _GEN_2048 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_74_data[32] ? 1'h0 : _GEN_1922; // @[lut_35.scala 2029:102 lut_35.scala 216:26]
  wire [5:0] _GEN_2049 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 6'h3 : _GEN_1923; // @[lut_35.scala 1987:102 lut_35.scala 1988:42]
  wire [31:0] _GEN_2050 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? push_ray_id : _GEN_1924; // @[lut_35.scala 1987:102 lut_35.scala 1989:42]
  wire  _GEN_2053 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _T_290; // @[lut_35.scala 1987:102 lut_35.scala 1996:42]
  wire  _GEN_2054 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1927; // @[lut_35.scala 1987:102 lut_35.scala 1997:42]
  wire  _GEN_2055 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1928; // @[lut_35.scala 1987:102 lut_35.scala 1998:42]
  wire  _GEN_2056 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1929; // @[lut_35.scala 1987:102 lut_35.scala 1999:42]
  wire  _GEN_2057 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1930; // @[lut_35.scala 1987:102 lut_35.scala 2000:42]
  wire  _GEN_2058 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1931; // @[lut_35.scala 1987:102 lut_35.scala 2001:42]
  wire  _GEN_2059 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1932; // @[lut_35.scala 1987:102 lut_35.scala 2002:43]
  wire  _GEN_2060 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1933; // @[lut_35.scala 1987:102 lut_35.scala 2003:43]
  wire  _GEN_2061 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1934; // @[lut_35.scala 1987:102 lut_35.scala 2004:43]
  wire  _GEN_2062 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1935; // @[lut_35.scala 1987:102 lut_35.scala 2005:43]
  wire  _GEN_2063 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1936; // @[lut_35.scala 1987:102 lut_35.scala 2006:43]
  wire  _GEN_2064 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1937; // @[lut_35.scala 1987:102 lut_35.scala 2007:43]
  wire  _GEN_2065 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1938; // @[lut_35.scala 1987:102 lut_35.scala 2008:43]
  wire  _GEN_2066 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1939; // @[lut_35.scala 1987:102 lut_35.scala 2009:43]
  wire  _GEN_2067 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1940; // @[lut_35.scala 1987:102 lut_35.scala 2010:43]
  wire  _GEN_2068 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1941; // @[lut_35.scala 1987:102 lut_35.scala 2011:43]
  wire  _GEN_2069 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1942; // @[lut_35.scala 1987:102 lut_35.scala 2012:43]
  wire  _GEN_2070 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1943; // @[lut_35.scala 1987:102 lut_35.scala 2013:43]
  wire  _GEN_2071 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1944; // @[lut_35.scala 1987:102 lut_35.scala 2014:43]
  wire  _GEN_2072 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1945; // @[lut_35.scala 1987:102 lut_35.scala 2015:43]
  wire  _GEN_2073 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1946; // @[lut_35.scala 1987:102 lut_35.scala 2016:43]
  wire  _GEN_2074 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1947; // @[lut_35.scala 1987:102 lut_35.scala 2017:43]
  wire  _GEN_2075 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1948; // @[lut_35.scala 1987:102 lut_35.scala 2018:43]
  wire  _GEN_2076 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1949; // @[lut_35.scala 1987:102 lut_35.scala 2019:43]
  wire  _GEN_2077 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1950; // @[lut_35.scala 1987:102 lut_35.scala 2020:43]
  wire  _GEN_2078 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1951; // @[lut_35.scala 1987:102 lut_35.scala 2021:43]
  wire  _GEN_2079 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1952; // @[lut_35.scala 1987:102 lut_35.scala 2022:43]
  wire  _GEN_2080 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1953; // @[lut_35.scala 1987:102 lut_35.scala 2023:43]
  wire  _GEN_2081 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1954; // @[lut_35.scala 1987:102 lut_35.scala 2024:43]
  wire  _GEN_2082 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1955; // @[lut_35.scala 1987:102 lut_35.scala 2025:43]
  wire  _GEN_2083 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1956; // @[lut_35.scala 1987:102 lut_35.scala 2026:43]
  wire  _GEN_2084 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] | _GEN_1957; // @[lut_35.scala 1987:102 lut_35.scala 2027:38]
  wire  _GEN_2088 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 1987:102 lut_35.scala 216:26 lut_35.scala 2029:87]
  wire  _GEN_2091 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1961; // @[lut_35.scala 1987:102 lut_35.scala 216:26]
  wire  _GEN_2094 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1964; // @[lut_35.scala 1987:102 lut_35.scala 216:26]
  wire  _GEN_2097 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1967; // @[lut_35.scala 1987:102 lut_35.scala 216:26]
  wire  _GEN_2100 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1970; // @[lut_35.scala 1987:102 lut_35.scala 216:26]
  wire  _GEN_2103 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1973; // @[lut_35.scala 1987:102 lut_35.scala 216:26]
  wire  _GEN_2106 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1976; // @[lut_35.scala 1987:102 lut_35.scala 216:26]
  wire  _GEN_2109 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1979; // @[lut_35.scala 1987:102 lut_35.scala 216:26]
  wire  _GEN_2112 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1982; // @[lut_35.scala 1987:102 lut_35.scala 216:26]
  wire  _GEN_2115 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1985; // @[lut_35.scala 1987:102 lut_35.scala 216:26]
  wire  _GEN_2118 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1988; // @[lut_35.scala 1987:102 lut_35.scala 216:26]
  wire  _GEN_2121 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1991; // @[lut_35.scala 1987:102 lut_35.scala 216:26]
  wire  _GEN_2124 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1994; // @[lut_35.scala 1987:102 lut_35.scala 216:26]
  wire  _GEN_2127 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_1997; // @[lut_35.scala 1987:102 lut_35.scala 216:26]
  wire  _GEN_2130 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_2000; // @[lut_35.scala 1987:102 lut_35.scala 216:26]
  wire  _GEN_2133 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_2003; // @[lut_35.scala 1987:102 lut_35.scala 216:26]
  wire  _GEN_2136 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_2006; // @[lut_35.scala 1987:102 lut_35.scala 216:26]
  wire  _GEN_2139 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_2009; // @[lut_35.scala 1987:102 lut_35.scala 216:26]
  wire  _GEN_2142 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_2012; // @[lut_35.scala 1987:102 lut_35.scala 216:26]
  wire  _GEN_2145 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_2015; // @[lut_35.scala 1987:102 lut_35.scala 216:26]
  wire  _GEN_2148 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_2018; // @[lut_35.scala 1987:102 lut_35.scala 216:26]
  wire  _GEN_2151 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_2021; // @[lut_35.scala 1987:102 lut_35.scala 216:26]
  wire  _GEN_2154 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_2024; // @[lut_35.scala 1987:102 lut_35.scala 216:26]
  wire  _GEN_2157 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_2027; // @[lut_35.scala 1987:102 lut_35.scala 216:26]
  wire  _GEN_2160 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_2030; // @[lut_35.scala 1987:102 lut_35.scala 216:26]
  wire  _GEN_2163 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_2033; // @[lut_35.scala 1987:102 lut_35.scala 216:26]
  wire  _GEN_2166 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_2036; // @[lut_35.scala 1987:102 lut_35.scala 216:26]
  wire  _GEN_2169 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_2039; // @[lut_35.scala 1987:102 lut_35.scala 216:26]
  wire  _GEN_2172 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_2042; // @[lut_35.scala 1987:102 lut_35.scala 216:26]
  wire  _GEN_2175 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_2045; // @[lut_35.scala 1987:102 lut_35.scala 216:26]
  wire  _GEN_2178 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_73_data[32] ? 1'h0 : _GEN_2048; // @[lut_35.scala 1987:102 lut_35.scala 216:26]
  wire [5:0] _GEN_2179 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 6'h2 : _GEN_2049; // @[lut_35.scala 1945:102 lut_35.scala 1946:42]
  wire [31:0] _GEN_2180 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? push_ray_id : _GEN_2050; // @[lut_35.scala 1945:102 lut_35.scala 1947:42]
  wire  _GEN_2183 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _T_282; // @[lut_35.scala 1945:102 lut_35.scala 1953:42]
  wire  _GEN_2184 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2053; // @[lut_35.scala 1945:102 lut_35.scala 1954:42]
  wire  _GEN_2185 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2054; // @[lut_35.scala 1945:102 lut_35.scala 1955:42]
  wire  _GEN_2186 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2055; // @[lut_35.scala 1945:102 lut_35.scala 1956:42]
  wire  _GEN_2187 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2056; // @[lut_35.scala 1945:102 lut_35.scala 1957:42]
  wire  _GEN_2188 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2057; // @[lut_35.scala 1945:102 lut_35.scala 1958:42]
  wire  _GEN_2189 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2058; // @[lut_35.scala 1945:102 lut_35.scala 1959:42]
  wire  _GEN_2190 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2059; // @[lut_35.scala 1945:102 lut_35.scala 1960:43]
  wire  _GEN_2191 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2060; // @[lut_35.scala 1945:102 lut_35.scala 1961:43]
  wire  _GEN_2192 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2061; // @[lut_35.scala 1945:102 lut_35.scala 1962:43]
  wire  _GEN_2193 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2062; // @[lut_35.scala 1945:102 lut_35.scala 1963:43]
  wire  _GEN_2194 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2063; // @[lut_35.scala 1945:102 lut_35.scala 1964:43]
  wire  _GEN_2195 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2064; // @[lut_35.scala 1945:102 lut_35.scala 1965:43]
  wire  _GEN_2196 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2065; // @[lut_35.scala 1945:102 lut_35.scala 1966:43]
  wire  _GEN_2197 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2066; // @[lut_35.scala 1945:102 lut_35.scala 1967:43]
  wire  _GEN_2198 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2067; // @[lut_35.scala 1945:102 lut_35.scala 1968:43]
  wire  _GEN_2199 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2068; // @[lut_35.scala 1945:102 lut_35.scala 1969:43]
  wire  _GEN_2200 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2069; // @[lut_35.scala 1945:102 lut_35.scala 1970:43]
  wire  _GEN_2201 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2070; // @[lut_35.scala 1945:102 lut_35.scala 1971:43]
  wire  _GEN_2202 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2071; // @[lut_35.scala 1945:102 lut_35.scala 1972:43]
  wire  _GEN_2203 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2072; // @[lut_35.scala 1945:102 lut_35.scala 1973:43]
  wire  _GEN_2204 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2073; // @[lut_35.scala 1945:102 lut_35.scala 1974:43]
  wire  _GEN_2205 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2074; // @[lut_35.scala 1945:102 lut_35.scala 1975:43]
  wire  _GEN_2206 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2075; // @[lut_35.scala 1945:102 lut_35.scala 1976:43]
  wire  _GEN_2207 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2076; // @[lut_35.scala 1945:102 lut_35.scala 1977:43]
  wire  _GEN_2208 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2077; // @[lut_35.scala 1945:102 lut_35.scala 1978:43]
  wire  _GEN_2209 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2078; // @[lut_35.scala 1945:102 lut_35.scala 1979:43]
  wire  _GEN_2210 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2079; // @[lut_35.scala 1945:102 lut_35.scala 1980:43]
  wire  _GEN_2211 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2080; // @[lut_35.scala 1945:102 lut_35.scala 1981:43]
  wire  _GEN_2212 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2081; // @[lut_35.scala 1945:102 lut_35.scala 1982:43]
  wire  _GEN_2213 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2082; // @[lut_35.scala 1945:102 lut_35.scala 1983:43]
  wire  _GEN_2214 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2083; // @[lut_35.scala 1945:102 lut_35.scala 1984:43]
  wire  _GEN_2215 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] | _GEN_2084; // @[lut_35.scala 1945:102 lut_35.scala 1985:38]
  wire  _GEN_2219 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 1945:102 lut_35.scala 216:26 lut_35.scala 1987:87]
  wire  _GEN_2222 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2088; // @[lut_35.scala 1945:102 lut_35.scala 216:26]
  wire  _GEN_2225 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2091; // @[lut_35.scala 1945:102 lut_35.scala 216:26]
  wire  _GEN_2228 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2094; // @[lut_35.scala 1945:102 lut_35.scala 216:26]
  wire  _GEN_2231 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2097; // @[lut_35.scala 1945:102 lut_35.scala 216:26]
  wire  _GEN_2234 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2100; // @[lut_35.scala 1945:102 lut_35.scala 216:26]
  wire  _GEN_2237 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2103; // @[lut_35.scala 1945:102 lut_35.scala 216:26]
  wire  _GEN_2240 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2106; // @[lut_35.scala 1945:102 lut_35.scala 216:26]
  wire  _GEN_2243 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2109; // @[lut_35.scala 1945:102 lut_35.scala 216:26]
  wire  _GEN_2246 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2112; // @[lut_35.scala 1945:102 lut_35.scala 216:26]
  wire  _GEN_2249 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2115; // @[lut_35.scala 1945:102 lut_35.scala 216:26]
  wire  _GEN_2252 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2118; // @[lut_35.scala 1945:102 lut_35.scala 216:26]
  wire  _GEN_2255 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2121; // @[lut_35.scala 1945:102 lut_35.scala 216:26]
  wire  _GEN_2258 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2124; // @[lut_35.scala 1945:102 lut_35.scala 216:26]
  wire  _GEN_2261 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2127; // @[lut_35.scala 1945:102 lut_35.scala 216:26]
  wire  _GEN_2264 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2130; // @[lut_35.scala 1945:102 lut_35.scala 216:26]
  wire  _GEN_2267 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2133; // @[lut_35.scala 1945:102 lut_35.scala 216:26]
  wire  _GEN_2270 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2136; // @[lut_35.scala 1945:102 lut_35.scala 216:26]
  wire  _GEN_2273 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2139; // @[lut_35.scala 1945:102 lut_35.scala 216:26]
  wire  _GEN_2276 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2142; // @[lut_35.scala 1945:102 lut_35.scala 216:26]
  wire  _GEN_2279 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2145; // @[lut_35.scala 1945:102 lut_35.scala 216:26]
  wire  _GEN_2282 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2148; // @[lut_35.scala 1945:102 lut_35.scala 216:26]
  wire  _GEN_2285 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2151; // @[lut_35.scala 1945:102 lut_35.scala 216:26]
  wire  _GEN_2288 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2154; // @[lut_35.scala 1945:102 lut_35.scala 216:26]
  wire  _GEN_2291 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2157; // @[lut_35.scala 1945:102 lut_35.scala 216:26]
  wire  _GEN_2294 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2160; // @[lut_35.scala 1945:102 lut_35.scala 216:26]
  wire  _GEN_2297 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2163; // @[lut_35.scala 1945:102 lut_35.scala 216:26]
  wire  _GEN_2300 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2166; // @[lut_35.scala 1945:102 lut_35.scala 216:26]
  wire  _GEN_2303 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2169; // @[lut_35.scala 1945:102 lut_35.scala 216:26]
  wire  _GEN_2306 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2172; // @[lut_35.scala 1945:102 lut_35.scala 216:26]
  wire  _GEN_2309 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2175; // @[lut_35.scala 1945:102 lut_35.scala 216:26]
  wire  _GEN_2312 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_72_data[32] ? 1'h0 : _GEN_2178; // @[lut_35.scala 1945:102 lut_35.scala 216:26]
  wire [5:0] _GEN_2313 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 6'h1 : _GEN_2179; // @[lut_35.scala 1903:102 lut_35.scala 1904:42]
  wire [31:0] _GEN_2314 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? push_ray_id : _GEN_2180; // @[lut_35.scala 1903:102 lut_35.scala 1905:42]
  wire  _GEN_2317 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _T_274; // @[lut_35.scala 1903:102 lut_35.scala 1910:42]
  wire  _GEN_2318 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2183; // @[lut_35.scala 1903:102 lut_35.scala 1911:42]
  wire  _GEN_2319 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2184; // @[lut_35.scala 1903:102 lut_35.scala 1912:42]
  wire  _GEN_2320 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2185; // @[lut_35.scala 1903:102 lut_35.scala 1913:42]
  wire  _GEN_2321 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2186; // @[lut_35.scala 1903:102 lut_35.scala 1914:42]
  wire  _GEN_2322 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2187; // @[lut_35.scala 1903:102 lut_35.scala 1915:42]
  wire  _GEN_2323 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2188; // @[lut_35.scala 1903:102 lut_35.scala 1916:42]
  wire  _GEN_2324 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2189; // @[lut_35.scala 1903:102 lut_35.scala 1917:42]
  wire  _GEN_2325 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2190; // @[lut_35.scala 1903:102 lut_35.scala 1918:43]
  wire  _GEN_2326 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2191; // @[lut_35.scala 1903:102 lut_35.scala 1919:43]
  wire  _GEN_2327 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2192; // @[lut_35.scala 1903:102 lut_35.scala 1920:43]
  wire  _GEN_2328 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2193; // @[lut_35.scala 1903:102 lut_35.scala 1921:43]
  wire  _GEN_2329 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2194; // @[lut_35.scala 1903:102 lut_35.scala 1922:43]
  wire  _GEN_2330 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2195; // @[lut_35.scala 1903:102 lut_35.scala 1923:43]
  wire  _GEN_2331 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2196; // @[lut_35.scala 1903:102 lut_35.scala 1924:43]
  wire  _GEN_2332 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2197; // @[lut_35.scala 1903:102 lut_35.scala 1925:43]
  wire  _GEN_2333 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2198; // @[lut_35.scala 1903:102 lut_35.scala 1926:43]
  wire  _GEN_2334 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2199; // @[lut_35.scala 1903:102 lut_35.scala 1927:43]
  wire  _GEN_2335 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2200; // @[lut_35.scala 1903:102 lut_35.scala 1928:43]
  wire  _GEN_2336 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2201; // @[lut_35.scala 1903:102 lut_35.scala 1929:43]
  wire  _GEN_2337 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2202; // @[lut_35.scala 1903:102 lut_35.scala 1930:43]
  wire  _GEN_2338 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2203; // @[lut_35.scala 1903:102 lut_35.scala 1931:43]
  wire  _GEN_2339 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2204; // @[lut_35.scala 1903:102 lut_35.scala 1932:43]
  wire  _GEN_2340 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2205; // @[lut_35.scala 1903:102 lut_35.scala 1933:43]
  wire  _GEN_2341 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2206; // @[lut_35.scala 1903:102 lut_35.scala 1934:43]
  wire  _GEN_2342 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2207; // @[lut_35.scala 1903:102 lut_35.scala 1935:43]
  wire  _GEN_2343 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2208; // @[lut_35.scala 1903:102 lut_35.scala 1936:43]
  wire  _GEN_2344 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2209; // @[lut_35.scala 1903:102 lut_35.scala 1937:43]
  wire  _GEN_2345 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2210; // @[lut_35.scala 1903:102 lut_35.scala 1938:43]
  wire  _GEN_2346 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2211; // @[lut_35.scala 1903:102 lut_35.scala 1939:43]
  wire  _GEN_2347 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2212; // @[lut_35.scala 1903:102 lut_35.scala 1940:43]
  wire  _GEN_2348 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2213; // @[lut_35.scala 1903:102 lut_35.scala 1941:43]
  wire  _GEN_2349 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2214; // @[lut_35.scala 1903:102 lut_35.scala 1942:43]
  wire  _GEN_2350 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] | _GEN_2215; // @[lut_35.scala 1903:102 lut_35.scala 1943:38]
  wire  _GEN_2354 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 1903:102 lut_35.scala 216:26 lut_35.scala 1945:87]
  wire  _GEN_2357 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2219; // @[lut_35.scala 1903:102 lut_35.scala 216:26]
  wire  _GEN_2360 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2222; // @[lut_35.scala 1903:102 lut_35.scala 216:26]
  wire  _GEN_2363 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2225; // @[lut_35.scala 1903:102 lut_35.scala 216:26]
  wire  _GEN_2366 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2228; // @[lut_35.scala 1903:102 lut_35.scala 216:26]
  wire  _GEN_2369 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2231; // @[lut_35.scala 1903:102 lut_35.scala 216:26]
  wire  _GEN_2372 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2234; // @[lut_35.scala 1903:102 lut_35.scala 216:26]
  wire  _GEN_2375 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2237; // @[lut_35.scala 1903:102 lut_35.scala 216:26]
  wire  _GEN_2378 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2240; // @[lut_35.scala 1903:102 lut_35.scala 216:26]
  wire  _GEN_2381 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2243; // @[lut_35.scala 1903:102 lut_35.scala 216:26]
  wire  _GEN_2384 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2246; // @[lut_35.scala 1903:102 lut_35.scala 216:26]
  wire  _GEN_2387 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2249; // @[lut_35.scala 1903:102 lut_35.scala 216:26]
  wire  _GEN_2390 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2252; // @[lut_35.scala 1903:102 lut_35.scala 216:26]
  wire  _GEN_2393 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2255; // @[lut_35.scala 1903:102 lut_35.scala 216:26]
  wire  _GEN_2396 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2258; // @[lut_35.scala 1903:102 lut_35.scala 216:26]
  wire  _GEN_2399 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2261; // @[lut_35.scala 1903:102 lut_35.scala 216:26]
  wire  _GEN_2402 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2264; // @[lut_35.scala 1903:102 lut_35.scala 216:26]
  wire  _GEN_2405 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2267; // @[lut_35.scala 1903:102 lut_35.scala 216:26]
  wire  _GEN_2408 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2270; // @[lut_35.scala 1903:102 lut_35.scala 216:26]
  wire  _GEN_2411 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2273; // @[lut_35.scala 1903:102 lut_35.scala 216:26]
  wire  _GEN_2414 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2276; // @[lut_35.scala 1903:102 lut_35.scala 216:26]
  wire  _GEN_2417 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2279; // @[lut_35.scala 1903:102 lut_35.scala 216:26]
  wire  _GEN_2420 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2282; // @[lut_35.scala 1903:102 lut_35.scala 216:26]
  wire  _GEN_2423 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2285; // @[lut_35.scala 1903:102 lut_35.scala 216:26]
  wire  _GEN_2426 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2288; // @[lut_35.scala 1903:102 lut_35.scala 216:26]
  wire  _GEN_2429 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2291; // @[lut_35.scala 1903:102 lut_35.scala 216:26]
  wire  _GEN_2432 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2294; // @[lut_35.scala 1903:102 lut_35.scala 216:26]
  wire  _GEN_2435 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2297; // @[lut_35.scala 1903:102 lut_35.scala 216:26]
  wire  _GEN_2438 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2300; // @[lut_35.scala 1903:102 lut_35.scala 216:26]
  wire  _GEN_2441 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2303; // @[lut_35.scala 1903:102 lut_35.scala 216:26]
  wire  _GEN_2444 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2306; // @[lut_35.scala 1903:102 lut_35.scala 216:26]
  wire  _GEN_2447 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2309; // @[lut_35.scala 1903:102 lut_35.scala 216:26]
  wire  _GEN_2450 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_71_data[32] ? 1'h0 : _GEN_2312; // @[lut_35.scala 1903:102 lut_35.scala 216:26]
  wire [5:0] _GEN_2451 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 6'h0 : _GEN_2313; // @[lut_35.scala 1861:103 lut_35.scala 1862:42]
  wire [31:0] _GEN_2452 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? push_ray_id : _GEN_2314; // @[lut_35.scala 1861:103 lut_35.scala 1863:42]
  wire  _GEN_2454 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _T_266; // @[lut_35.scala 1861:103 lut_35.scala 1867:42]
  wire  _GEN_2455 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2317; // @[lut_35.scala 1861:103 lut_35.scala 1868:42]
  wire  _GEN_2456 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2318; // @[lut_35.scala 1861:103 lut_35.scala 1869:42]
  wire  _GEN_2457 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2319; // @[lut_35.scala 1861:103 lut_35.scala 1870:42]
  wire  _GEN_2458 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2320; // @[lut_35.scala 1861:103 lut_35.scala 1871:42]
  wire  _GEN_2459 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2321; // @[lut_35.scala 1861:103 lut_35.scala 1872:42]
  wire  _GEN_2460 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2322; // @[lut_35.scala 1861:103 lut_35.scala 1873:42]
  wire  _GEN_2461 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2323; // @[lut_35.scala 1861:103 lut_35.scala 1874:42]
  wire  _GEN_2462 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2324; // @[lut_35.scala 1861:103 lut_35.scala 1875:42]
  wire  _GEN_2463 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2325; // @[lut_35.scala 1861:103 lut_35.scala 1876:43]
  wire  _GEN_2464 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2326; // @[lut_35.scala 1861:103 lut_35.scala 1877:43]
  wire  _GEN_2465 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2327; // @[lut_35.scala 1861:103 lut_35.scala 1878:43]
  wire  _GEN_2466 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2328; // @[lut_35.scala 1861:103 lut_35.scala 1879:43]
  wire  _GEN_2467 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2329; // @[lut_35.scala 1861:103 lut_35.scala 1880:43]
  wire  _GEN_2468 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2330; // @[lut_35.scala 1861:103 lut_35.scala 1881:43]
  wire  _GEN_2469 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2331; // @[lut_35.scala 1861:103 lut_35.scala 1882:43]
  wire  _GEN_2470 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2332; // @[lut_35.scala 1861:103 lut_35.scala 1883:43]
  wire  _GEN_2471 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2333; // @[lut_35.scala 1861:103 lut_35.scala 1884:43]
  wire  _GEN_2472 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2334; // @[lut_35.scala 1861:103 lut_35.scala 1885:43]
  wire  _GEN_2473 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2335; // @[lut_35.scala 1861:103 lut_35.scala 1886:43]
  wire  _GEN_2474 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2336; // @[lut_35.scala 1861:103 lut_35.scala 1887:43]
  wire  _GEN_2475 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2337; // @[lut_35.scala 1861:103 lut_35.scala 1888:43]
  wire  _GEN_2476 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2338; // @[lut_35.scala 1861:103 lut_35.scala 1889:43]
  wire  _GEN_2477 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2339; // @[lut_35.scala 1861:103 lut_35.scala 1890:43]
  wire  _GEN_2478 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2340; // @[lut_35.scala 1861:103 lut_35.scala 1891:43]
  wire  _GEN_2479 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2341; // @[lut_35.scala 1861:103 lut_35.scala 1892:43]
  wire  _GEN_2480 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2342; // @[lut_35.scala 1861:103 lut_35.scala 1893:43]
  wire  _GEN_2481 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2343; // @[lut_35.scala 1861:103 lut_35.scala 1894:43]
  wire  _GEN_2482 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2344; // @[lut_35.scala 1861:103 lut_35.scala 1895:43]
  wire  _GEN_2483 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2345; // @[lut_35.scala 1861:103 lut_35.scala 1896:43]
  wire  _GEN_2484 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2346; // @[lut_35.scala 1861:103 lut_35.scala 1897:43]
  wire  _GEN_2485 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2347; // @[lut_35.scala 1861:103 lut_35.scala 1898:43]
  wire  _GEN_2486 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2348; // @[lut_35.scala 1861:103 lut_35.scala 1899:43]
  wire  _GEN_2487 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2349; // @[lut_35.scala 1861:103 lut_35.scala 1900:43]
  wire  _GEN_2488 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] | _GEN_2350; // @[lut_35.scala 1861:103 lut_35.scala 1901:38]
  wire  _GEN_2492 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 1861:103 lut_35.scala 216:26 lut_35.scala 1903:87]
  wire  _GEN_2495 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2354; // @[lut_35.scala 1861:103 lut_35.scala 216:26]
  wire  _GEN_2498 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2357; // @[lut_35.scala 1861:103 lut_35.scala 216:26]
  wire  _GEN_2501 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2360; // @[lut_35.scala 1861:103 lut_35.scala 216:26]
  wire  _GEN_2504 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2363; // @[lut_35.scala 1861:103 lut_35.scala 216:26]
  wire  _GEN_2507 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2366; // @[lut_35.scala 1861:103 lut_35.scala 216:26]
  wire  _GEN_2510 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2369; // @[lut_35.scala 1861:103 lut_35.scala 216:26]
  wire  _GEN_2513 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2372; // @[lut_35.scala 1861:103 lut_35.scala 216:26]
  wire  _GEN_2516 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2375; // @[lut_35.scala 1861:103 lut_35.scala 216:26]
  wire  _GEN_2519 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2378; // @[lut_35.scala 1861:103 lut_35.scala 216:26]
  wire  _GEN_2522 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2381; // @[lut_35.scala 1861:103 lut_35.scala 216:26]
  wire  _GEN_2525 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2384; // @[lut_35.scala 1861:103 lut_35.scala 216:26]
  wire  _GEN_2528 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2387; // @[lut_35.scala 1861:103 lut_35.scala 216:26]
  wire  _GEN_2531 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2390; // @[lut_35.scala 1861:103 lut_35.scala 216:26]
  wire  _GEN_2534 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2393; // @[lut_35.scala 1861:103 lut_35.scala 216:26]
  wire  _GEN_2537 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2396; // @[lut_35.scala 1861:103 lut_35.scala 216:26]
  wire  _GEN_2540 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2399; // @[lut_35.scala 1861:103 lut_35.scala 216:26]
  wire  _GEN_2543 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2402; // @[lut_35.scala 1861:103 lut_35.scala 216:26]
  wire  _GEN_2546 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2405; // @[lut_35.scala 1861:103 lut_35.scala 216:26]
  wire  _GEN_2549 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2408; // @[lut_35.scala 1861:103 lut_35.scala 216:26]
  wire  _GEN_2552 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2411; // @[lut_35.scala 1861:103 lut_35.scala 216:26]
  wire  _GEN_2555 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2414; // @[lut_35.scala 1861:103 lut_35.scala 216:26]
  wire  _GEN_2558 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2417; // @[lut_35.scala 1861:103 lut_35.scala 216:26]
  wire  _GEN_2561 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2420; // @[lut_35.scala 1861:103 lut_35.scala 216:26]
  wire  _GEN_2564 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2423; // @[lut_35.scala 1861:103 lut_35.scala 216:26]
  wire  _GEN_2567 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2426; // @[lut_35.scala 1861:103 lut_35.scala 216:26]
  wire  _GEN_2570 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2429; // @[lut_35.scala 1861:103 lut_35.scala 216:26]
  wire  _GEN_2573 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2432; // @[lut_35.scala 1861:103 lut_35.scala 216:26]
  wire  _GEN_2576 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2435; // @[lut_35.scala 1861:103 lut_35.scala 216:26]
  wire  _GEN_2579 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2438; // @[lut_35.scala 1861:103 lut_35.scala 216:26]
  wire  _GEN_2582 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2441; // @[lut_35.scala 1861:103 lut_35.scala 216:26]
  wire  _GEN_2585 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2444; // @[lut_35.scala 1861:103 lut_35.scala 216:26]
  wire  _GEN_2588 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2447; // @[lut_35.scala 1861:103 lut_35.scala 216:26]
  wire  _GEN_2591 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_70_data[32] ? 1'h0 : _GEN_2450; // @[lut_35.scala 1861:103 lut_35.scala 216:26]
  wire [5:0] _GEN_2595 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 !=
    push_ray_id & push_valid ? _GEN_2451 : 6'h23; // @[lut_35.scala 1860:125 lut_35.scala 3373:42]
  wire [31:0] _GEN_2596 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 !=
    push_ray_id & push_valid ? _GEN_2452 : 32'h0; // @[lut_35.scala 1860:125 lut_35.scala 3374:42]
  wire  _GEN_2597 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _T_258; // @[lut_35.scala 1860:125 lut_35.scala 3375:32]
  wire  _GEN_2598 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2454; // @[lut_35.scala 1860:125 lut_35.scala 3376:32]
  wire  _GEN_2599 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2455; // @[lut_35.scala 1860:125 lut_35.scala 3377:32]
  wire  _GEN_2600 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2456; // @[lut_35.scala 1860:125 lut_35.scala 3378:32]
  wire  _GEN_2601 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2457; // @[lut_35.scala 1860:125 lut_35.scala 3379:32]
  wire  _GEN_2602 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2458; // @[lut_35.scala 1860:125 lut_35.scala 3380:32]
  wire  _GEN_2603 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2459; // @[lut_35.scala 1860:125 lut_35.scala 3381:32]
  wire  _GEN_2604 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2460; // @[lut_35.scala 1860:125 lut_35.scala 3382:32]
  wire  _GEN_2605 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2461; // @[lut_35.scala 1860:125 lut_35.scala 3383:42]
  wire  _GEN_2606 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2462; // @[lut_35.scala 1860:125 lut_35.scala 3384:42]
  wire  _GEN_2607 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2463; // @[lut_35.scala 1860:125 lut_35.scala 3385:43]
  wire  _GEN_2608 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2464; // @[lut_35.scala 1860:125 lut_35.scala 3386:43]
  wire  _GEN_2609 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2465; // @[lut_35.scala 1860:125 lut_35.scala 3387:43]
  wire  _GEN_2610 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2466; // @[lut_35.scala 1860:125 lut_35.scala 3388:43]
  wire  _GEN_2611 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2467; // @[lut_35.scala 1860:125 lut_35.scala 3389:43]
  wire  _GEN_2612 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2468; // @[lut_35.scala 1860:125 lut_35.scala 3390:43]
  wire  _GEN_2613 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2469; // @[lut_35.scala 1860:125 lut_35.scala 3391:43]
  wire  _GEN_2614 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2470; // @[lut_35.scala 1860:125 lut_35.scala 3392:43]
  wire  _GEN_2615 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2471; // @[lut_35.scala 1860:125 lut_35.scala 3393:43]
  wire  _GEN_2616 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2472; // @[lut_35.scala 1860:125 lut_35.scala 3394:43]
  wire  _GEN_2617 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2473; // @[lut_35.scala 1860:125 lut_35.scala 3395:43]
  wire  _GEN_2618 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2474; // @[lut_35.scala 1860:125 lut_35.scala 3396:43]
  wire  _GEN_2619 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2475; // @[lut_35.scala 1860:125 lut_35.scala 3397:43]
  wire  _GEN_2620 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2476; // @[lut_35.scala 1860:125 lut_35.scala 3398:43]
  wire  _GEN_2621 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2477; // @[lut_35.scala 1860:125 lut_35.scala 3399:43]
  wire  _GEN_2622 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2478; // @[lut_35.scala 1860:125 lut_35.scala 3400:43]
  wire  _GEN_2623 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2479; // @[lut_35.scala 1860:125 lut_35.scala 3401:43]
  wire  _GEN_2624 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2480; // @[lut_35.scala 1860:125 lut_35.scala 3402:43]
  wire  _GEN_2625 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2481; // @[lut_35.scala 1860:125 lut_35.scala 3403:43]
  wire  _GEN_2626 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2482; // @[lut_35.scala 1860:125 lut_35.scala 3404:43]
  wire  _GEN_2627 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2483; // @[lut_35.scala 1860:125 lut_35.scala 3405:43]
  wire  _GEN_2628 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2484; // @[lut_35.scala 1860:125 lut_35.scala 3406:43]
  wire  _GEN_2629 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2485; // @[lut_35.scala 1860:125 lut_35.scala 3407:43]
  wire  _GEN_2630 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2486; // @[lut_35.scala 1860:125 lut_35.scala 3408:43]
  wire  _GEN_2631 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2487; // @[lut_35.scala 1860:125 lut_35.scala 3409:43]
  wire  _GEN_2632 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2488; // @[lut_35.scala 1860:125 lut_35.scala 3410:30]
  wire  _GEN_2636 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2492; // @[lut_35.scala 1860:125 lut_35.scala 216:26]
  wire  _GEN_2639 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2495; // @[lut_35.scala 1860:125 lut_35.scala 216:26]
  wire  _GEN_2642 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2498; // @[lut_35.scala 1860:125 lut_35.scala 216:26]
  wire  _GEN_2645 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2501; // @[lut_35.scala 1860:125 lut_35.scala 216:26]
  wire  _GEN_2648 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2504; // @[lut_35.scala 1860:125 lut_35.scala 216:26]
  wire  _GEN_2651 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2507; // @[lut_35.scala 1860:125 lut_35.scala 216:26]
  wire  _GEN_2654 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2510; // @[lut_35.scala 1860:125 lut_35.scala 216:26]
  wire  _GEN_2657 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2513; // @[lut_35.scala 1860:125 lut_35.scala 216:26]
  wire  _GEN_2660 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2516; // @[lut_35.scala 1860:125 lut_35.scala 216:26]
  wire  _GEN_2663 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2519; // @[lut_35.scala 1860:125 lut_35.scala 216:26]
  wire  _GEN_2666 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2522; // @[lut_35.scala 1860:125 lut_35.scala 216:26]
  wire  _GEN_2669 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2525; // @[lut_35.scala 1860:125 lut_35.scala 216:26]
  wire  _GEN_2672 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2528; // @[lut_35.scala 1860:125 lut_35.scala 216:26]
  wire  _GEN_2675 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2531; // @[lut_35.scala 1860:125 lut_35.scala 216:26]
  wire  _GEN_2678 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2534; // @[lut_35.scala 1860:125 lut_35.scala 216:26]
  wire  _GEN_2681 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2537; // @[lut_35.scala 1860:125 lut_35.scala 216:26]
  wire  _GEN_2684 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2540; // @[lut_35.scala 1860:125 lut_35.scala 216:26]
  wire  _GEN_2687 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2543; // @[lut_35.scala 1860:125 lut_35.scala 216:26]
  wire  _GEN_2690 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2546; // @[lut_35.scala 1860:125 lut_35.scala 216:26]
  wire  _GEN_2693 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2549; // @[lut_35.scala 1860:125 lut_35.scala 216:26]
  wire  _GEN_2696 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2552; // @[lut_35.scala 1860:125 lut_35.scala 216:26]
  wire  _GEN_2699 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2555; // @[lut_35.scala 1860:125 lut_35.scala 216:26]
  wire  _GEN_2702 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2558; // @[lut_35.scala 1860:125 lut_35.scala 216:26]
  wire  _GEN_2705 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2561; // @[lut_35.scala 1860:125 lut_35.scala 216:26]
  wire  _GEN_2708 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2564; // @[lut_35.scala 1860:125 lut_35.scala 216:26]
  wire  _GEN_2711 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2567; // @[lut_35.scala 1860:125 lut_35.scala 216:26]
  wire  _GEN_2714 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2570; // @[lut_35.scala 1860:125 lut_35.scala 216:26]
  wire  _GEN_2717 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2573; // @[lut_35.scala 1860:125 lut_35.scala 216:26]
  wire  _GEN_2720 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2576; // @[lut_35.scala 1860:125 lut_35.scala 216:26]
  wire  _GEN_2723 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2579; // @[lut_35.scala 1860:125 lut_35.scala 216:26]
  wire  _GEN_2726 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2582; // @[lut_35.scala 1860:125 lut_35.scala 216:26]
  wire  _GEN_2729 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2585; // @[lut_35.scala 1860:125 lut_35.scala 216:26]
  wire  _GEN_2732 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2588; // @[lut_35.scala 1860:125 lut_35.scala 216:26]
  wire  _GEN_2735 = _T_242 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_2591; // @[lut_35.scala 1860:125 lut_35.scala 216:26]
  wire  _GEN_2736 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2597; // @[lut_35.scala 1817:74 lut_35.scala 1818:38]
  wire  _GEN_2737 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2598; // @[lut_35.scala 1817:74 lut_35.scala 1819:38]
  wire  _GEN_2738 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2599; // @[lut_35.scala 1817:74 lut_35.scala 1820:38]
  wire  _GEN_2739 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2600; // @[lut_35.scala 1817:74 lut_35.scala 1821:38]
  wire  _GEN_2740 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2601; // @[lut_35.scala 1817:74 lut_35.scala 1822:38]
  wire  _GEN_2741 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2602; // @[lut_35.scala 1817:74 lut_35.scala 1823:38]
  wire  _GEN_2742 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2603; // @[lut_35.scala 1817:74 lut_35.scala 1824:38]
  wire  _GEN_2743 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2604; // @[lut_35.scala 1817:74 lut_35.scala 1825:38]
  wire  _GEN_2744 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2605; // @[lut_35.scala 1817:74 lut_35.scala 1826:38]
  wire  _GEN_2745 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2606; // @[lut_35.scala 1817:74 lut_35.scala 1827:38]
  wire  _GEN_2746 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2607; // @[lut_35.scala 1817:74 lut_35.scala 1828:39]
  wire  _GEN_2747 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2608; // @[lut_35.scala 1817:74 lut_35.scala 1829:39]
  wire  _GEN_2748 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2609; // @[lut_35.scala 1817:74 lut_35.scala 1830:39]
  wire  _GEN_2749 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2610; // @[lut_35.scala 1817:74 lut_35.scala 1831:39]
  wire  _GEN_2750 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2611; // @[lut_35.scala 1817:74 lut_35.scala 1832:39]
  wire  _GEN_2751 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2612; // @[lut_35.scala 1817:74 lut_35.scala 1833:39]
  wire  _GEN_2752 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2613; // @[lut_35.scala 1817:74 lut_35.scala 1834:39]
  wire  _GEN_2753 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2614; // @[lut_35.scala 1817:74 lut_35.scala 1835:39]
  wire  _GEN_2754 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2615; // @[lut_35.scala 1817:74 lut_35.scala 1836:39]
  wire  _GEN_2755 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2616; // @[lut_35.scala 1817:74 lut_35.scala 1837:39]
  wire  _GEN_2756 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2617; // @[lut_35.scala 1817:74 lut_35.scala 1838:39]
  wire  _GEN_2757 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2618; // @[lut_35.scala 1817:74 lut_35.scala 1839:39]
  wire  _GEN_2758 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2619; // @[lut_35.scala 1817:74 lut_35.scala 1840:39]
  wire  _GEN_2759 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2620; // @[lut_35.scala 1817:74 lut_35.scala 1841:39]
  wire  _GEN_2760 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2621; // @[lut_35.scala 1817:74 lut_35.scala 1842:39]
  wire  _GEN_2761 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2622; // @[lut_35.scala 1817:74 lut_35.scala 1843:39]
  wire  _GEN_2762 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2623; // @[lut_35.scala 1817:74 lut_35.scala 1844:39]
  wire  _GEN_2763 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2624; // @[lut_35.scala 1817:74 lut_35.scala 1845:39]
  wire  _GEN_2764 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2625; // @[lut_35.scala 1817:74 lut_35.scala 1846:39]
  wire  _GEN_2765 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2626; // @[lut_35.scala 1817:74 lut_35.scala 1847:39]
  wire  _GEN_2766 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2627; // @[lut_35.scala 1817:74 lut_35.scala 1848:39]
  wire  _GEN_2767 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2628; // @[lut_35.scala 1817:74 lut_35.scala 1849:39]
  wire  _GEN_2768 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2629; // @[lut_35.scala 1817:74 lut_35.scala 1850:39]
  wire  _GEN_2769 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2630; // @[lut_35.scala 1817:74 lut_35.scala 1851:39]
  wire  _GEN_2770 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid | _GEN_2631; // @[lut_35.scala 1817:74 lut_35.scala 1852:39]
  wire  _GEN_2771 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid | _GEN_2632; // @[lut_35.scala 1817:74 lut_35.scala 1853:34]
  wire  _GEN_2775 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _T_250; // @[lut_35.scala 1817:74 lut_35.scala 216:26]
  wire [5:0] _GEN_2776 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? push_mem_temp : _GEN_2595; // @[lut_35.scala 1817:74 lut_35.scala 521:39]
  wire [31:0] _GEN_2777 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? push_id_temp : _GEN_2596; // @[lut_35.scala 1817:74 lut_35.scala 522:39]
  wire  _GEN_2780 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2636; // @[lut_35.scala 1817:74 lut_35.scala 216:26]
  wire  _GEN_2783 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2639; // @[lut_35.scala 1817:74 lut_35.scala 216:26]
  wire  _GEN_2786 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2642; // @[lut_35.scala 1817:74 lut_35.scala 216:26]
  wire  _GEN_2789 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2645; // @[lut_35.scala 1817:74 lut_35.scala 216:26]
  wire  _GEN_2792 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2648; // @[lut_35.scala 1817:74 lut_35.scala 216:26]
  wire  _GEN_2795 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2651; // @[lut_35.scala 1817:74 lut_35.scala 216:26]
  wire  _GEN_2798 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2654; // @[lut_35.scala 1817:74 lut_35.scala 216:26]
  wire  _GEN_2801 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2657; // @[lut_35.scala 1817:74 lut_35.scala 216:26]
  wire  _GEN_2804 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2660; // @[lut_35.scala 1817:74 lut_35.scala 216:26]
  wire  _GEN_2807 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2663; // @[lut_35.scala 1817:74 lut_35.scala 216:26]
  wire  _GEN_2810 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2666; // @[lut_35.scala 1817:74 lut_35.scala 216:26]
  wire  _GEN_2813 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2669; // @[lut_35.scala 1817:74 lut_35.scala 216:26]
  wire  _GEN_2816 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2672; // @[lut_35.scala 1817:74 lut_35.scala 216:26]
  wire  _GEN_2819 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2675; // @[lut_35.scala 1817:74 lut_35.scala 216:26]
  wire  _GEN_2822 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2678; // @[lut_35.scala 1817:74 lut_35.scala 216:26]
  wire  _GEN_2825 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2681; // @[lut_35.scala 1817:74 lut_35.scala 216:26]
  wire  _GEN_2828 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2684; // @[lut_35.scala 1817:74 lut_35.scala 216:26]
  wire  _GEN_2831 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2687; // @[lut_35.scala 1817:74 lut_35.scala 216:26]
  wire  _GEN_2834 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2690; // @[lut_35.scala 1817:74 lut_35.scala 216:26]
  wire  _GEN_2837 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2693; // @[lut_35.scala 1817:74 lut_35.scala 216:26]
  wire  _GEN_2840 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2696; // @[lut_35.scala 1817:74 lut_35.scala 216:26]
  wire  _GEN_2843 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2699; // @[lut_35.scala 1817:74 lut_35.scala 216:26]
  wire  _GEN_2846 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2702; // @[lut_35.scala 1817:74 lut_35.scala 216:26]
  wire  _GEN_2849 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2705; // @[lut_35.scala 1817:74 lut_35.scala 216:26]
  wire  _GEN_2852 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2708; // @[lut_35.scala 1817:74 lut_35.scala 216:26]
  wire  _GEN_2855 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2711; // @[lut_35.scala 1817:74 lut_35.scala 216:26]
  wire  _GEN_2858 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2714; // @[lut_35.scala 1817:74 lut_35.scala 216:26]
  wire  _GEN_2861 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2717; // @[lut_35.scala 1817:74 lut_35.scala 216:26]
  wire  _GEN_2864 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2720; // @[lut_35.scala 1817:74 lut_35.scala 216:26]
  wire  _GEN_2867 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2723; // @[lut_35.scala 1817:74 lut_35.scala 216:26]
  wire  _GEN_2870 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2726; // @[lut_35.scala 1817:74 lut_35.scala 216:26]
  wire  _GEN_2873 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2729; // @[lut_35.scala 1817:74 lut_35.scala 216:26]
  wire  _GEN_2876 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2732; // @[lut_35.scala 1817:74 lut_35.scala 216:26]
  wire  _GEN_2879 = LUT_mem_MPORT_69_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2735; // @[lut_35.scala 1817:74 lut_35.scala 216:26]
  wire  _GEN_2880 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2736; // @[lut_35.scala 1779:74 lut_35.scala 1780:38]
  wire  _GEN_2881 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2737; // @[lut_35.scala 1779:74 lut_35.scala 1781:38]
  wire  _GEN_2882 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2738; // @[lut_35.scala 1779:74 lut_35.scala 1782:38]
  wire  _GEN_2883 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2739; // @[lut_35.scala 1779:74 lut_35.scala 1783:38]
  wire  _GEN_2884 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2740; // @[lut_35.scala 1779:74 lut_35.scala 1784:38]
  wire  _GEN_2885 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2741; // @[lut_35.scala 1779:74 lut_35.scala 1785:38]
  wire  _GEN_2886 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2742; // @[lut_35.scala 1779:74 lut_35.scala 1786:38]
  wire  _GEN_2887 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2743; // @[lut_35.scala 1779:74 lut_35.scala 1787:38]
  wire  _GEN_2888 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2744; // @[lut_35.scala 1779:74 lut_35.scala 1788:38]
  wire  _GEN_2889 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2745; // @[lut_35.scala 1779:74 lut_35.scala 1789:38]
  wire  _GEN_2890 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2746; // @[lut_35.scala 1779:74 lut_35.scala 1790:39]
  wire  _GEN_2891 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2747; // @[lut_35.scala 1779:74 lut_35.scala 1791:39]
  wire  _GEN_2892 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2748; // @[lut_35.scala 1779:74 lut_35.scala 1792:39]
  wire  _GEN_2893 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2749; // @[lut_35.scala 1779:74 lut_35.scala 1793:39]
  wire  _GEN_2894 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2750; // @[lut_35.scala 1779:74 lut_35.scala 1794:39]
  wire  _GEN_2895 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2751; // @[lut_35.scala 1779:74 lut_35.scala 1795:39]
  wire  _GEN_2896 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2752; // @[lut_35.scala 1779:74 lut_35.scala 1796:39]
  wire  _GEN_2897 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2753; // @[lut_35.scala 1779:74 lut_35.scala 1797:39]
  wire  _GEN_2898 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2754; // @[lut_35.scala 1779:74 lut_35.scala 1798:39]
  wire  _GEN_2899 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2755; // @[lut_35.scala 1779:74 lut_35.scala 1799:39]
  wire  _GEN_2900 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2756; // @[lut_35.scala 1779:74 lut_35.scala 1800:39]
  wire  _GEN_2901 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2757; // @[lut_35.scala 1779:74 lut_35.scala 1801:39]
  wire  _GEN_2902 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2758; // @[lut_35.scala 1779:74 lut_35.scala 1802:39]
  wire  _GEN_2903 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2759; // @[lut_35.scala 1779:74 lut_35.scala 1803:39]
  wire  _GEN_2904 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2760; // @[lut_35.scala 1779:74 lut_35.scala 1804:39]
  wire  _GEN_2905 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2761; // @[lut_35.scala 1779:74 lut_35.scala 1805:39]
  wire  _GEN_2906 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2762; // @[lut_35.scala 1779:74 lut_35.scala 1806:39]
  wire  _GEN_2907 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2763; // @[lut_35.scala 1779:74 lut_35.scala 1807:39]
  wire  _GEN_2908 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2764; // @[lut_35.scala 1779:74 lut_35.scala 1808:39]
  wire  _GEN_2909 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2765; // @[lut_35.scala 1779:74 lut_35.scala 1809:39]
  wire  _GEN_2910 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2766; // @[lut_35.scala 1779:74 lut_35.scala 1810:39]
  wire  _GEN_2911 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2767; // @[lut_35.scala 1779:74 lut_35.scala 1811:39]
  wire  _GEN_2912 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2768; // @[lut_35.scala 1779:74 lut_35.scala 1812:39]
  wire  _GEN_2913 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid | _GEN_2769; // @[lut_35.scala 1779:74 lut_35.scala 1813:39]
  wire  _GEN_2914 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2770; // @[lut_35.scala 1779:74 lut_35.scala 1814:39]
  wire  _GEN_2915 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid | _GEN_2771; // @[lut_35.scala 1779:74 lut_35.scala 1815:34]
  wire  _GEN_2919 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1779:74 lut_35.scala 216:26 lut_35.scala 1817:27]
  wire  _GEN_2922 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2775; // @[lut_35.scala 1779:74 lut_35.scala 216:26]
  wire [5:0] _GEN_2923 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? push_mem_temp : _GEN_2776; // @[lut_35.scala 1779:74 lut_35.scala 521:39]
  wire [31:0] _GEN_2924 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? push_id_temp : _GEN_2777; // @[lut_35.scala 1779:74 lut_35.scala 522:39]
  wire  _GEN_2927 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2780; // @[lut_35.scala 1779:74 lut_35.scala 216:26]
  wire  _GEN_2930 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2783; // @[lut_35.scala 1779:74 lut_35.scala 216:26]
  wire  _GEN_2933 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2786; // @[lut_35.scala 1779:74 lut_35.scala 216:26]
  wire  _GEN_2936 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2789; // @[lut_35.scala 1779:74 lut_35.scala 216:26]
  wire  _GEN_2939 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2792; // @[lut_35.scala 1779:74 lut_35.scala 216:26]
  wire  _GEN_2942 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2795; // @[lut_35.scala 1779:74 lut_35.scala 216:26]
  wire  _GEN_2945 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2798; // @[lut_35.scala 1779:74 lut_35.scala 216:26]
  wire  _GEN_2948 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2801; // @[lut_35.scala 1779:74 lut_35.scala 216:26]
  wire  _GEN_2951 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2804; // @[lut_35.scala 1779:74 lut_35.scala 216:26]
  wire  _GEN_2954 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2807; // @[lut_35.scala 1779:74 lut_35.scala 216:26]
  wire  _GEN_2957 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2810; // @[lut_35.scala 1779:74 lut_35.scala 216:26]
  wire  _GEN_2960 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2813; // @[lut_35.scala 1779:74 lut_35.scala 216:26]
  wire  _GEN_2963 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2816; // @[lut_35.scala 1779:74 lut_35.scala 216:26]
  wire  _GEN_2966 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2819; // @[lut_35.scala 1779:74 lut_35.scala 216:26]
  wire  _GEN_2969 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2822; // @[lut_35.scala 1779:74 lut_35.scala 216:26]
  wire  _GEN_2972 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2825; // @[lut_35.scala 1779:74 lut_35.scala 216:26]
  wire  _GEN_2975 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2828; // @[lut_35.scala 1779:74 lut_35.scala 216:26]
  wire  _GEN_2978 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2831; // @[lut_35.scala 1779:74 lut_35.scala 216:26]
  wire  _GEN_2981 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2834; // @[lut_35.scala 1779:74 lut_35.scala 216:26]
  wire  _GEN_2984 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2837; // @[lut_35.scala 1779:74 lut_35.scala 216:26]
  wire  _GEN_2987 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2840; // @[lut_35.scala 1779:74 lut_35.scala 216:26]
  wire  _GEN_2990 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2843; // @[lut_35.scala 1779:74 lut_35.scala 216:26]
  wire  _GEN_2993 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2846; // @[lut_35.scala 1779:74 lut_35.scala 216:26]
  wire  _GEN_2996 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2849; // @[lut_35.scala 1779:74 lut_35.scala 216:26]
  wire  _GEN_2999 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2852; // @[lut_35.scala 1779:74 lut_35.scala 216:26]
  wire  _GEN_3002 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2855; // @[lut_35.scala 1779:74 lut_35.scala 216:26]
  wire  _GEN_3005 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2858; // @[lut_35.scala 1779:74 lut_35.scala 216:26]
  wire  _GEN_3008 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2861; // @[lut_35.scala 1779:74 lut_35.scala 216:26]
  wire  _GEN_3011 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2864; // @[lut_35.scala 1779:74 lut_35.scala 216:26]
  wire  _GEN_3014 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2867; // @[lut_35.scala 1779:74 lut_35.scala 216:26]
  wire  _GEN_3017 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2870; // @[lut_35.scala 1779:74 lut_35.scala 216:26]
  wire  _GEN_3020 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2873; // @[lut_35.scala 1779:74 lut_35.scala 216:26]
  wire  _GEN_3023 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2876; // @[lut_35.scala 1779:74 lut_35.scala 216:26]
  wire  _GEN_3026 = LUT_mem_MPORT_68_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2879; // @[lut_35.scala 1779:74 lut_35.scala 216:26]
  wire  _GEN_3027 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2880; // @[lut_35.scala 1741:74 lut_35.scala 1742:38]
  wire  _GEN_3028 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2881; // @[lut_35.scala 1741:74 lut_35.scala 1743:38]
  wire  _GEN_3029 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2882; // @[lut_35.scala 1741:74 lut_35.scala 1744:38]
  wire  _GEN_3030 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2883; // @[lut_35.scala 1741:74 lut_35.scala 1745:38]
  wire  _GEN_3031 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2884; // @[lut_35.scala 1741:74 lut_35.scala 1746:38]
  wire  _GEN_3032 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2885; // @[lut_35.scala 1741:74 lut_35.scala 1747:38]
  wire  _GEN_3033 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2886; // @[lut_35.scala 1741:74 lut_35.scala 1748:38]
  wire  _GEN_3034 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2887; // @[lut_35.scala 1741:74 lut_35.scala 1749:38]
  wire  _GEN_3035 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2888; // @[lut_35.scala 1741:74 lut_35.scala 1750:38]
  wire  _GEN_3036 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2889; // @[lut_35.scala 1741:74 lut_35.scala 1751:38]
  wire  _GEN_3037 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2890; // @[lut_35.scala 1741:74 lut_35.scala 1752:39]
  wire  _GEN_3038 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2891; // @[lut_35.scala 1741:74 lut_35.scala 1753:39]
  wire  _GEN_3039 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2892; // @[lut_35.scala 1741:74 lut_35.scala 1754:39]
  wire  _GEN_3040 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2893; // @[lut_35.scala 1741:74 lut_35.scala 1755:39]
  wire  _GEN_3041 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2894; // @[lut_35.scala 1741:74 lut_35.scala 1756:39]
  wire  _GEN_3042 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2895; // @[lut_35.scala 1741:74 lut_35.scala 1757:39]
  wire  _GEN_3043 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2896; // @[lut_35.scala 1741:74 lut_35.scala 1758:39]
  wire  _GEN_3044 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2897; // @[lut_35.scala 1741:74 lut_35.scala 1759:39]
  wire  _GEN_3045 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2898; // @[lut_35.scala 1741:74 lut_35.scala 1760:39]
  wire  _GEN_3046 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2899; // @[lut_35.scala 1741:74 lut_35.scala 1761:39]
  wire  _GEN_3047 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2900; // @[lut_35.scala 1741:74 lut_35.scala 1762:39]
  wire  _GEN_3048 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2901; // @[lut_35.scala 1741:74 lut_35.scala 1763:39]
  wire  _GEN_3049 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2902; // @[lut_35.scala 1741:74 lut_35.scala 1764:39]
  wire  _GEN_3050 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2903; // @[lut_35.scala 1741:74 lut_35.scala 1765:39]
  wire  _GEN_3051 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2904; // @[lut_35.scala 1741:74 lut_35.scala 1766:39]
  wire  _GEN_3052 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2905; // @[lut_35.scala 1741:74 lut_35.scala 1767:39]
  wire  _GEN_3053 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2906; // @[lut_35.scala 1741:74 lut_35.scala 1768:39]
  wire  _GEN_3054 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2907; // @[lut_35.scala 1741:74 lut_35.scala 1769:39]
  wire  _GEN_3055 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2908; // @[lut_35.scala 1741:74 lut_35.scala 1770:39]
  wire  _GEN_3056 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2909; // @[lut_35.scala 1741:74 lut_35.scala 1771:39]
  wire  _GEN_3057 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2910; // @[lut_35.scala 1741:74 lut_35.scala 1772:39]
  wire  _GEN_3058 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2911; // @[lut_35.scala 1741:74 lut_35.scala 1773:39]
  wire  _GEN_3059 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid | _GEN_2912; // @[lut_35.scala 1741:74 lut_35.scala 1774:39]
  wire  _GEN_3060 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2913; // @[lut_35.scala 1741:74 lut_35.scala 1775:39]
  wire  _GEN_3061 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2914; // @[lut_35.scala 1741:74 lut_35.scala 1776:39]
  wire  _GEN_3062 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid | _GEN_2915; // @[lut_35.scala 1741:74 lut_35.scala 1777:34]
  wire  _GEN_3066 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1741:74 lut_35.scala 216:26 lut_35.scala 1779:27]
  wire  _GEN_3069 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2919; // @[lut_35.scala 1741:74 lut_35.scala 216:26]
  wire  _GEN_3072 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2922; // @[lut_35.scala 1741:74 lut_35.scala 216:26]
  wire [5:0] _GEN_3073 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? push_mem_temp : _GEN_2923; // @[lut_35.scala 1741:74 lut_35.scala 521:39]
  wire [31:0] _GEN_3074 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? push_id_temp : _GEN_2924; // @[lut_35.scala 1741:74 lut_35.scala 522:39]
  wire  _GEN_3077 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2927; // @[lut_35.scala 1741:74 lut_35.scala 216:26]
  wire  _GEN_3080 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2930; // @[lut_35.scala 1741:74 lut_35.scala 216:26]
  wire  _GEN_3083 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2933; // @[lut_35.scala 1741:74 lut_35.scala 216:26]
  wire  _GEN_3086 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2936; // @[lut_35.scala 1741:74 lut_35.scala 216:26]
  wire  _GEN_3089 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2939; // @[lut_35.scala 1741:74 lut_35.scala 216:26]
  wire  _GEN_3092 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2942; // @[lut_35.scala 1741:74 lut_35.scala 216:26]
  wire  _GEN_3095 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2945; // @[lut_35.scala 1741:74 lut_35.scala 216:26]
  wire  _GEN_3098 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2948; // @[lut_35.scala 1741:74 lut_35.scala 216:26]
  wire  _GEN_3101 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2951; // @[lut_35.scala 1741:74 lut_35.scala 216:26]
  wire  _GEN_3104 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2954; // @[lut_35.scala 1741:74 lut_35.scala 216:26]
  wire  _GEN_3107 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2957; // @[lut_35.scala 1741:74 lut_35.scala 216:26]
  wire  _GEN_3110 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2960; // @[lut_35.scala 1741:74 lut_35.scala 216:26]
  wire  _GEN_3113 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2963; // @[lut_35.scala 1741:74 lut_35.scala 216:26]
  wire  _GEN_3116 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2966; // @[lut_35.scala 1741:74 lut_35.scala 216:26]
  wire  _GEN_3119 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2969; // @[lut_35.scala 1741:74 lut_35.scala 216:26]
  wire  _GEN_3122 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2972; // @[lut_35.scala 1741:74 lut_35.scala 216:26]
  wire  _GEN_3125 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2975; // @[lut_35.scala 1741:74 lut_35.scala 216:26]
  wire  _GEN_3128 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2978; // @[lut_35.scala 1741:74 lut_35.scala 216:26]
  wire  _GEN_3131 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2981; // @[lut_35.scala 1741:74 lut_35.scala 216:26]
  wire  _GEN_3134 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2984; // @[lut_35.scala 1741:74 lut_35.scala 216:26]
  wire  _GEN_3137 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2987; // @[lut_35.scala 1741:74 lut_35.scala 216:26]
  wire  _GEN_3140 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2990; // @[lut_35.scala 1741:74 lut_35.scala 216:26]
  wire  _GEN_3143 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2993; // @[lut_35.scala 1741:74 lut_35.scala 216:26]
  wire  _GEN_3146 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2996; // @[lut_35.scala 1741:74 lut_35.scala 216:26]
  wire  _GEN_3149 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_2999; // @[lut_35.scala 1741:74 lut_35.scala 216:26]
  wire  _GEN_3152 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3002; // @[lut_35.scala 1741:74 lut_35.scala 216:26]
  wire  _GEN_3155 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3005; // @[lut_35.scala 1741:74 lut_35.scala 216:26]
  wire  _GEN_3158 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3008; // @[lut_35.scala 1741:74 lut_35.scala 216:26]
  wire  _GEN_3161 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3011; // @[lut_35.scala 1741:74 lut_35.scala 216:26]
  wire  _GEN_3164 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3014; // @[lut_35.scala 1741:74 lut_35.scala 216:26]
  wire  _GEN_3167 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3017; // @[lut_35.scala 1741:74 lut_35.scala 216:26]
  wire  _GEN_3170 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3020; // @[lut_35.scala 1741:74 lut_35.scala 216:26]
  wire  _GEN_3173 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3023; // @[lut_35.scala 1741:74 lut_35.scala 216:26]
  wire  _GEN_3176 = LUT_mem_MPORT_67_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3026; // @[lut_35.scala 1741:74 lut_35.scala 216:26]
  wire  _GEN_3177 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3027; // @[lut_35.scala 1703:74 lut_35.scala 1704:38]
  wire  _GEN_3178 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3028; // @[lut_35.scala 1703:74 lut_35.scala 1705:38]
  wire  _GEN_3179 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3029; // @[lut_35.scala 1703:74 lut_35.scala 1706:38]
  wire  _GEN_3180 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3030; // @[lut_35.scala 1703:74 lut_35.scala 1707:38]
  wire  _GEN_3181 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3031; // @[lut_35.scala 1703:74 lut_35.scala 1708:38]
  wire  _GEN_3182 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3032; // @[lut_35.scala 1703:74 lut_35.scala 1709:38]
  wire  _GEN_3183 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3033; // @[lut_35.scala 1703:74 lut_35.scala 1710:38]
  wire  _GEN_3184 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3034; // @[lut_35.scala 1703:74 lut_35.scala 1711:38]
  wire  _GEN_3185 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3035; // @[lut_35.scala 1703:74 lut_35.scala 1712:38]
  wire  _GEN_3186 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3036; // @[lut_35.scala 1703:74 lut_35.scala 1713:38]
  wire  _GEN_3187 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3037; // @[lut_35.scala 1703:74 lut_35.scala 1714:39]
  wire  _GEN_3188 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3038; // @[lut_35.scala 1703:74 lut_35.scala 1715:39]
  wire  _GEN_3189 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3039; // @[lut_35.scala 1703:74 lut_35.scala 1716:39]
  wire  _GEN_3190 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3040; // @[lut_35.scala 1703:74 lut_35.scala 1717:39]
  wire  _GEN_3191 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3041; // @[lut_35.scala 1703:74 lut_35.scala 1718:39]
  wire  _GEN_3192 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3042; // @[lut_35.scala 1703:74 lut_35.scala 1719:39]
  wire  _GEN_3193 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3043; // @[lut_35.scala 1703:74 lut_35.scala 1720:39]
  wire  _GEN_3194 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3044; // @[lut_35.scala 1703:74 lut_35.scala 1721:39]
  wire  _GEN_3195 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3045; // @[lut_35.scala 1703:74 lut_35.scala 1722:39]
  wire  _GEN_3196 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3046; // @[lut_35.scala 1703:74 lut_35.scala 1723:39]
  wire  _GEN_3197 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3047; // @[lut_35.scala 1703:74 lut_35.scala 1724:39]
  wire  _GEN_3198 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3048; // @[lut_35.scala 1703:74 lut_35.scala 1725:39]
  wire  _GEN_3199 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3049; // @[lut_35.scala 1703:74 lut_35.scala 1726:39]
  wire  _GEN_3200 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3050; // @[lut_35.scala 1703:74 lut_35.scala 1727:39]
  wire  _GEN_3201 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3051; // @[lut_35.scala 1703:74 lut_35.scala 1728:39]
  wire  _GEN_3202 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3052; // @[lut_35.scala 1703:74 lut_35.scala 1729:39]
  wire  _GEN_3203 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3053; // @[lut_35.scala 1703:74 lut_35.scala 1730:39]
  wire  _GEN_3204 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3054; // @[lut_35.scala 1703:74 lut_35.scala 1731:39]
  wire  _GEN_3205 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3055; // @[lut_35.scala 1703:74 lut_35.scala 1732:39]
  wire  _GEN_3206 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3056; // @[lut_35.scala 1703:74 lut_35.scala 1733:39]
  wire  _GEN_3207 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3057; // @[lut_35.scala 1703:74 lut_35.scala 1734:39]
  wire  _GEN_3208 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid | _GEN_3058; // @[lut_35.scala 1703:74 lut_35.scala 1735:39]
  wire  _GEN_3209 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3059; // @[lut_35.scala 1703:74 lut_35.scala 1736:39]
  wire  _GEN_3210 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3060; // @[lut_35.scala 1703:74 lut_35.scala 1737:39]
  wire  _GEN_3211 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3061; // @[lut_35.scala 1703:74 lut_35.scala 1738:39]
  wire  _GEN_3212 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid | _GEN_3062; // @[lut_35.scala 1703:74 lut_35.scala 1739:34]
  wire  _GEN_3216 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1703:74 lut_35.scala 216:26 lut_35.scala 1741:27]
  wire  _GEN_3219 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3066; // @[lut_35.scala 1703:74 lut_35.scala 216:26]
  wire  _GEN_3222 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3069; // @[lut_35.scala 1703:74 lut_35.scala 216:26]
  wire  _GEN_3225 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3072; // @[lut_35.scala 1703:74 lut_35.scala 216:26]
  wire [5:0] _GEN_3226 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? push_mem_temp : _GEN_3073; // @[lut_35.scala 1703:74 lut_35.scala 521:39]
  wire [31:0] _GEN_3227 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? push_id_temp : _GEN_3074; // @[lut_35.scala 1703:74 lut_35.scala 522:39]
  wire  _GEN_3230 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3077; // @[lut_35.scala 1703:74 lut_35.scala 216:26]
  wire  _GEN_3233 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3080; // @[lut_35.scala 1703:74 lut_35.scala 216:26]
  wire  _GEN_3236 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3083; // @[lut_35.scala 1703:74 lut_35.scala 216:26]
  wire  _GEN_3239 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3086; // @[lut_35.scala 1703:74 lut_35.scala 216:26]
  wire  _GEN_3242 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3089; // @[lut_35.scala 1703:74 lut_35.scala 216:26]
  wire  _GEN_3245 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3092; // @[lut_35.scala 1703:74 lut_35.scala 216:26]
  wire  _GEN_3248 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3095; // @[lut_35.scala 1703:74 lut_35.scala 216:26]
  wire  _GEN_3251 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3098; // @[lut_35.scala 1703:74 lut_35.scala 216:26]
  wire  _GEN_3254 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3101; // @[lut_35.scala 1703:74 lut_35.scala 216:26]
  wire  _GEN_3257 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3104; // @[lut_35.scala 1703:74 lut_35.scala 216:26]
  wire  _GEN_3260 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3107; // @[lut_35.scala 1703:74 lut_35.scala 216:26]
  wire  _GEN_3263 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3110; // @[lut_35.scala 1703:74 lut_35.scala 216:26]
  wire  _GEN_3266 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3113; // @[lut_35.scala 1703:74 lut_35.scala 216:26]
  wire  _GEN_3269 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3116; // @[lut_35.scala 1703:74 lut_35.scala 216:26]
  wire  _GEN_3272 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3119; // @[lut_35.scala 1703:74 lut_35.scala 216:26]
  wire  _GEN_3275 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3122; // @[lut_35.scala 1703:74 lut_35.scala 216:26]
  wire  _GEN_3278 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3125; // @[lut_35.scala 1703:74 lut_35.scala 216:26]
  wire  _GEN_3281 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3128; // @[lut_35.scala 1703:74 lut_35.scala 216:26]
  wire  _GEN_3284 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3131; // @[lut_35.scala 1703:74 lut_35.scala 216:26]
  wire  _GEN_3287 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3134; // @[lut_35.scala 1703:74 lut_35.scala 216:26]
  wire  _GEN_3290 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3137; // @[lut_35.scala 1703:74 lut_35.scala 216:26]
  wire  _GEN_3293 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3140; // @[lut_35.scala 1703:74 lut_35.scala 216:26]
  wire  _GEN_3296 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3143; // @[lut_35.scala 1703:74 lut_35.scala 216:26]
  wire  _GEN_3299 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3146; // @[lut_35.scala 1703:74 lut_35.scala 216:26]
  wire  _GEN_3302 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3149; // @[lut_35.scala 1703:74 lut_35.scala 216:26]
  wire  _GEN_3305 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3152; // @[lut_35.scala 1703:74 lut_35.scala 216:26]
  wire  _GEN_3308 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3155; // @[lut_35.scala 1703:74 lut_35.scala 216:26]
  wire  _GEN_3311 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3158; // @[lut_35.scala 1703:74 lut_35.scala 216:26]
  wire  _GEN_3314 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3161; // @[lut_35.scala 1703:74 lut_35.scala 216:26]
  wire  _GEN_3317 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3164; // @[lut_35.scala 1703:74 lut_35.scala 216:26]
  wire  _GEN_3320 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3167; // @[lut_35.scala 1703:74 lut_35.scala 216:26]
  wire  _GEN_3323 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3170; // @[lut_35.scala 1703:74 lut_35.scala 216:26]
  wire  _GEN_3326 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3173; // @[lut_35.scala 1703:74 lut_35.scala 216:26]
  wire  _GEN_3329 = LUT_mem_MPORT_66_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3176; // @[lut_35.scala 1703:74 lut_35.scala 216:26]
  wire  _GEN_3330 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3177; // @[lut_35.scala 1665:74 lut_35.scala 1666:38]
  wire  _GEN_3331 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3178; // @[lut_35.scala 1665:74 lut_35.scala 1667:38]
  wire  _GEN_3332 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3179; // @[lut_35.scala 1665:74 lut_35.scala 1668:38]
  wire  _GEN_3333 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3180; // @[lut_35.scala 1665:74 lut_35.scala 1669:38]
  wire  _GEN_3334 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3181; // @[lut_35.scala 1665:74 lut_35.scala 1670:38]
  wire  _GEN_3335 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3182; // @[lut_35.scala 1665:74 lut_35.scala 1671:38]
  wire  _GEN_3336 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3183; // @[lut_35.scala 1665:74 lut_35.scala 1672:38]
  wire  _GEN_3337 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3184; // @[lut_35.scala 1665:74 lut_35.scala 1673:38]
  wire  _GEN_3338 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3185; // @[lut_35.scala 1665:74 lut_35.scala 1674:38]
  wire  _GEN_3339 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3186; // @[lut_35.scala 1665:74 lut_35.scala 1675:38]
  wire  _GEN_3340 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3187; // @[lut_35.scala 1665:74 lut_35.scala 1676:39]
  wire  _GEN_3341 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3188; // @[lut_35.scala 1665:74 lut_35.scala 1677:39]
  wire  _GEN_3342 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3189; // @[lut_35.scala 1665:74 lut_35.scala 1678:39]
  wire  _GEN_3343 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3190; // @[lut_35.scala 1665:74 lut_35.scala 1679:39]
  wire  _GEN_3344 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3191; // @[lut_35.scala 1665:74 lut_35.scala 1680:39]
  wire  _GEN_3345 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3192; // @[lut_35.scala 1665:74 lut_35.scala 1681:39]
  wire  _GEN_3346 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3193; // @[lut_35.scala 1665:74 lut_35.scala 1682:39]
  wire  _GEN_3347 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3194; // @[lut_35.scala 1665:74 lut_35.scala 1683:39]
  wire  _GEN_3348 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3195; // @[lut_35.scala 1665:74 lut_35.scala 1684:39]
  wire  _GEN_3349 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3196; // @[lut_35.scala 1665:74 lut_35.scala 1685:39]
  wire  _GEN_3350 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3197; // @[lut_35.scala 1665:74 lut_35.scala 1686:39]
  wire  _GEN_3351 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3198; // @[lut_35.scala 1665:74 lut_35.scala 1687:39]
  wire  _GEN_3352 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3199; // @[lut_35.scala 1665:74 lut_35.scala 1688:39]
  wire  _GEN_3353 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3200; // @[lut_35.scala 1665:74 lut_35.scala 1689:39]
  wire  _GEN_3354 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3201; // @[lut_35.scala 1665:74 lut_35.scala 1690:39]
  wire  _GEN_3355 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3202; // @[lut_35.scala 1665:74 lut_35.scala 1691:39]
  wire  _GEN_3356 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3203; // @[lut_35.scala 1665:74 lut_35.scala 1692:39]
  wire  _GEN_3357 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3204; // @[lut_35.scala 1665:74 lut_35.scala 1693:39]
  wire  _GEN_3358 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3205; // @[lut_35.scala 1665:74 lut_35.scala 1694:39]
  wire  _GEN_3359 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3206; // @[lut_35.scala 1665:74 lut_35.scala 1695:39]
  wire  _GEN_3360 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid | _GEN_3207; // @[lut_35.scala 1665:74 lut_35.scala 1696:39]
  wire  _GEN_3361 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3208; // @[lut_35.scala 1665:74 lut_35.scala 1697:39]
  wire  _GEN_3362 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3209; // @[lut_35.scala 1665:74 lut_35.scala 1698:39]
  wire  _GEN_3363 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3210; // @[lut_35.scala 1665:74 lut_35.scala 1699:39]
  wire  _GEN_3364 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3211; // @[lut_35.scala 1665:74 lut_35.scala 1700:39]
  wire  _GEN_3365 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid | _GEN_3212; // @[lut_35.scala 1665:74 lut_35.scala 1701:34]
  wire  _GEN_3369 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1665:74 lut_35.scala 216:26 lut_35.scala 1703:27]
  wire  _GEN_3372 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3216; // @[lut_35.scala 1665:74 lut_35.scala 216:26]
  wire  _GEN_3375 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3219; // @[lut_35.scala 1665:74 lut_35.scala 216:26]
  wire  _GEN_3378 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3222; // @[lut_35.scala 1665:74 lut_35.scala 216:26]
  wire  _GEN_3381 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3225; // @[lut_35.scala 1665:74 lut_35.scala 216:26]
  wire [5:0] _GEN_3382 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? push_mem_temp : _GEN_3226; // @[lut_35.scala 1665:74 lut_35.scala 521:39]
  wire [31:0] _GEN_3383 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? push_id_temp : _GEN_3227; // @[lut_35.scala 1665:74 lut_35.scala 522:39]
  wire  _GEN_3386 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3230; // @[lut_35.scala 1665:74 lut_35.scala 216:26]
  wire  _GEN_3389 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3233; // @[lut_35.scala 1665:74 lut_35.scala 216:26]
  wire  _GEN_3392 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3236; // @[lut_35.scala 1665:74 lut_35.scala 216:26]
  wire  _GEN_3395 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3239; // @[lut_35.scala 1665:74 lut_35.scala 216:26]
  wire  _GEN_3398 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3242; // @[lut_35.scala 1665:74 lut_35.scala 216:26]
  wire  _GEN_3401 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3245; // @[lut_35.scala 1665:74 lut_35.scala 216:26]
  wire  _GEN_3404 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3248; // @[lut_35.scala 1665:74 lut_35.scala 216:26]
  wire  _GEN_3407 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3251; // @[lut_35.scala 1665:74 lut_35.scala 216:26]
  wire  _GEN_3410 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3254; // @[lut_35.scala 1665:74 lut_35.scala 216:26]
  wire  _GEN_3413 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3257; // @[lut_35.scala 1665:74 lut_35.scala 216:26]
  wire  _GEN_3416 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3260; // @[lut_35.scala 1665:74 lut_35.scala 216:26]
  wire  _GEN_3419 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3263; // @[lut_35.scala 1665:74 lut_35.scala 216:26]
  wire  _GEN_3422 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3266; // @[lut_35.scala 1665:74 lut_35.scala 216:26]
  wire  _GEN_3425 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3269; // @[lut_35.scala 1665:74 lut_35.scala 216:26]
  wire  _GEN_3428 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3272; // @[lut_35.scala 1665:74 lut_35.scala 216:26]
  wire  _GEN_3431 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3275; // @[lut_35.scala 1665:74 lut_35.scala 216:26]
  wire  _GEN_3434 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3278; // @[lut_35.scala 1665:74 lut_35.scala 216:26]
  wire  _GEN_3437 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3281; // @[lut_35.scala 1665:74 lut_35.scala 216:26]
  wire  _GEN_3440 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3284; // @[lut_35.scala 1665:74 lut_35.scala 216:26]
  wire  _GEN_3443 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3287; // @[lut_35.scala 1665:74 lut_35.scala 216:26]
  wire  _GEN_3446 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3290; // @[lut_35.scala 1665:74 lut_35.scala 216:26]
  wire  _GEN_3449 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3293; // @[lut_35.scala 1665:74 lut_35.scala 216:26]
  wire  _GEN_3452 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3296; // @[lut_35.scala 1665:74 lut_35.scala 216:26]
  wire  _GEN_3455 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3299; // @[lut_35.scala 1665:74 lut_35.scala 216:26]
  wire  _GEN_3458 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3302; // @[lut_35.scala 1665:74 lut_35.scala 216:26]
  wire  _GEN_3461 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3305; // @[lut_35.scala 1665:74 lut_35.scala 216:26]
  wire  _GEN_3464 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3308; // @[lut_35.scala 1665:74 lut_35.scala 216:26]
  wire  _GEN_3467 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3311; // @[lut_35.scala 1665:74 lut_35.scala 216:26]
  wire  _GEN_3470 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3314; // @[lut_35.scala 1665:74 lut_35.scala 216:26]
  wire  _GEN_3473 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3317; // @[lut_35.scala 1665:74 lut_35.scala 216:26]
  wire  _GEN_3476 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3320; // @[lut_35.scala 1665:74 lut_35.scala 216:26]
  wire  _GEN_3479 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3323; // @[lut_35.scala 1665:74 lut_35.scala 216:26]
  wire  _GEN_3482 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3326; // @[lut_35.scala 1665:74 lut_35.scala 216:26]
  wire  _GEN_3485 = LUT_mem_MPORT_65_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3329; // @[lut_35.scala 1665:74 lut_35.scala 216:26]
  wire  _GEN_3486 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3330; // @[lut_35.scala 1627:74 lut_35.scala 1628:38]
  wire  _GEN_3487 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3331; // @[lut_35.scala 1627:74 lut_35.scala 1629:38]
  wire  _GEN_3488 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3332; // @[lut_35.scala 1627:74 lut_35.scala 1630:38]
  wire  _GEN_3489 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3333; // @[lut_35.scala 1627:74 lut_35.scala 1631:38]
  wire  _GEN_3490 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3334; // @[lut_35.scala 1627:74 lut_35.scala 1632:38]
  wire  _GEN_3491 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3335; // @[lut_35.scala 1627:74 lut_35.scala 1633:38]
  wire  _GEN_3492 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3336; // @[lut_35.scala 1627:74 lut_35.scala 1634:38]
  wire  _GEN_3493 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3337; // @[lut_35.scala 1627:74 lut_35.scala 1635:38]
  wire  _GEN_3494 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3338; // @[lut_35.scala 1627:74 lut_35.scala 1636:38]
  wire  _GEN_3495 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3339; // @[lut_35.scala 1627:74 lut_35.scala 1637:38]
  wire  _GEN_3496 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3340; // @[lut_35.scala 1627:74 lut_35.scala 1638:39]
  wire  _GEN_3497 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3341; // @[lut_35.scala 1627:74 lut_35.scala 1639:39]
  wire  _GEN_3498 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3342; // @[lut_35.scala 1627:74 lut_35.scala 1640:39]
  wire  _GEN_3499 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3343; // @[lut_35.scala 1627:74 lut_35.scala 1641:39]
  wire  _GEN_3500 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3344; // @[lut_35.scala 1627:74 lut_35.scala 1642:39]
  wire  _GEN_3501 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3345; // @[lut_35.scala 1627:74 lut_35.scala 1643:39]
  wire  _GEN_3502 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3346; // @[lut_35.scala 1627:74 lut_35.scala 1644:39]
  wire  _GEN_3503 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3347; // @[lut_35.scala 1627:74 lut_35.scala 1645:39]
  wire  _GEN_3504 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3348; // @[lut_35.scala 1627:74 lut_35.scala 1646:39]
  wire  _GEN_3505 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3349; // @[lut_35.scala 1627:74 lut_35.scala 1647:39]
  wire  _GEN_3506 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3350; // @[lut_35.scala 1627:74 lut_35.scala 1648:39]
  wire  _GEN_3507 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3351; // @[lut_35.scala 1627:74 lut_35.scala 1649:39]
  wire  _GEN_3508 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3352; // @[lut_35.scala 1627:74 lut_35.scala 1650:39]
  wire  _GEN_3509 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3353; // @[lut_35.scala 1627:74 lut_35.scala 1651:39]
  wire  _GEN_3510 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3354; // @[lut_35.scala 1627:74 lut_35.scala 1652:39]
  wire  _GEN_3511 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3355; // @[lut_35.scala 1627:74 lut_35.scala 1653:39]
  wire  _GEN_3512 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3356; // @[lut_35.scala 1627:74 lut_35.scala 1654:39]
  wire  _GEN_3513 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3357; // @[lut_35.scala 1627:74 lut_35.scala 1655:39]
  wire  _GEN_3514 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3358; // @[lut_35.scala 1627:74 lut_35.scala 1656:39]
  wire  _GEN_3515 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid | _GEN_3359; // @[lut_35.scala 1627:74 lut_35.scala 1657:39]
  wire  _GEN_3516 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3360; // @[lut_35.scala 1627:74 lut_35.scala 1658:39]
  wire  _GEN_3517 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3361; // @[lut_35.scala 1627:74 lut_35.scala 1659:39]
  wire  _GEN_3518 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3362; // @[lut_35.scala 1627:74 lut_35.scala 1660:39]
  wire  _GEN_3519 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3363; // @[lut_35.scala 1627:74 lut_35.scala 1661:39]
  wire  _GEN_3520 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3364; // @[lut_35.scala 1627:74 lut_35.scala 1662:39]
  wire  _GEN_3521 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid | _GEN_3365; // @[lut_35.scala 1627:74 lut_35.scala 1663:34]
  wire  _GEN_3525 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1627:74 lut_35.scala 216:26 lut_35.scala 1665:27]
  wire  _GEN_3528 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3369; // @[lut_35.scala 1627:74 lut_35.scala 216:26]
  wire  _GEN_3531 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3372; // @[lut_35.scala 1627:74 lut_35.scala 216:26]
  wire  _GEN_3534 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3375; // @[lut_35.scala 1627:74 lut_35.scala 216:26]
  wire  _GEN_3537 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3378; // @[lut_35.scala 1627:74 lut_35.scala 216:26]
  wire  _GEN_3540 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3381; // @[lut_35.scala 1627:74 lut_35.scala 216:26]
  wire [5:0] _GEN_3541 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? push_mem_temp : _GEN_3382; // @[lut_35.scala 1627:74 lut_35.scala 521:39]
  wire [31:0] _GEN_3542 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? push_id_temp : _GEN_3383; // @[lut_35.scala 1627:74 lut_35.scala 522:39]
  wire  _GEN_3545 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3386; // @[lut_35.scala 1627:74 lut_35.scala 216:26]
  wire  _GEN_3548 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3389; // @[lut_35.scala 1627:74 lut_35.scala 216:26]
  wire  _GEN_3551 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3392; // @[lut_35.scala 1627:74 lut_35.scala 216:26]
  wire  _GEN_3554 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3395; // @[lut_35.scala 1627:74 lut_35.scala 216:26]
  wire  _GEN_3557 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3398; // @[lut_35.scala 1627:74 lut_35.scala 216:26]
  wire  _GEN_3560 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3401; // @[lut_35.scala 1627:74 lut_35.scala 216:26]
  wire  _GEN_3563 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3404; // @[lut_35.scala 1627:74 lut_35.scala 216:26]
  wire  _GEN_3566 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3407; // @[lut_35.scala 1627:74 lut_35.scala 216:26]
  wire  _GEN_3569 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3410; // @[lut_35.scala 1627:74 lut_35.scala 216:26]
  wire  _GEN_3572 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3413; // @[lut_35.scala 1627:74 lut_35.scala 216:26]
  wire  _GEN_3575 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3416; // @[lut_35.scala 1627:74 lut_35.scala 216:26]
  wire  _GEN_3578 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3419; // @[lut_35.scala 1627:74 lut_35.scala 216:26]
  wire  _GEN_3581 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3422; // @[lut_35.scala 1627:74 lut_35.scala 216:26]
  wire  _GEN_3584 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3425; // @[lut_35.scala 1627:74 lut_35.scala 216:26]
  wire  _GEN_3587 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3428; // @[lut_35.scala 1627:74 lut_35.scala 216:26]
  wire  _GEN_3590 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3431; // @[lut_35.scala 1627:74 lut_35.scala 216:26]
  wire  _GEN_3593 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3434; // @[lut_35.scala 1627:74 lut_35.scala 216:26]
  wire  _GEN_3596 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3437; // @[lut_35.scala 1627:74 lut_35.scala 216:26]
  wire  _GEN_3599 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3440; // @[lut_35.scala 1627:74 lut_35.scala 216:26]
  wire  _GEN_3602 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3443; // @[lut_35.scala 1627:74 lut_35.scala 216:26]
  wire  _GEN_3605 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3446; // @[lut_35.scala 1627:74 lut_35.scala 216:26]
  wire  _GEN_3608 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3449; // @[lut_35.scala 1627:74 lut_35.scala 216:26]
  wire  _GEN_3611 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3452; // @[lut_35.scala 1627:74 lut_35.scala 216:26]
  wire  _GEN_3614 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3455; // @[lut_35.scala 1627:74 lut_35.scala 216:26]
  wire  _GEN_3617 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3458; // @[lut_35.scala 1627:74 lut_35.scala 216:26]
  wire  _GEN_3620 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3461; // @[lut_35.scala 1627:74 lut_35.scala 216:26]
  wire  _GEN_3623 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3464; // @[lut_35.scala 1627:74 lut_35.scala 216:26]
  wire  _GEN_3626 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3467; // @[lut_35.scala 1627:74 lut_35.scala 216:26]
  wire  _GEN_3629 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3470; // @[lut_35.scala 1627:74 lut_35.scala 216:26]
  wire  _GEN_3632 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3473; // @[lut_35.scala 1627:74 lut_35.scala 216:26]
  wire  _GEN_3635 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3476; // @[lut_35.scala 1627:74 lut_35.scala 216:26]
  wire  _GEN_3638 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3479; // @[lut_35.scala 1627:74 lut_35.scala 216:26]
  wire  _GEN_3641 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3482; // @[lut_35.scala 1627:74 lut_35.scala 216:26]
  wire  _GEN_3644 = LUT_mem_MPORT_64_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3485; // @[lut_35.scala 1627:74 lut_35.scala 216:26]
  wire  _GEN_3645 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3486; // @[lut_35.scala 1589:74 lut_35.scala 1590:38]
  wire  _GEN_3646 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3487; // @[lut_35.scala 1589:74 lut_35.scala 1591:38]
  wire  _GEN_3647 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3488; // @[lut_35.scala 1589:74 lut_35.scala 1592:38]
  wire  _GEN_3648 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3489; // @[lut_35.scala 1589:74 lut_35.scala 1593:38]
  wire  _GEN_3649 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3490; // @[lut_35.scala 1589:74 lut_35.scala 1594:38]
  wire  _GEN_3650 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3491; // @[lut_35.scala 1589:74 lut_35.scala 1595:38]
  wire  _GEN_3651 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3492; // @[lut_35.scala 1589:74 lut_35.scala 1596:38]
  wire  _GEN_3652 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3493; // @[lut_35.scala 1589:74 lut_35.scala 1597:38]
  wire  _GEN_3653 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3494; // @[lut_35.scala 1589:74 lut_35.scala 1598:38]
  wire  _GEN_3654 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3495; // @[lut_35.scala 1589:74 lut_35.scala 1599:38]
  wire  _GEN_3655 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3496; // @[lut_35.scala 1589:74 lut_35.scala 1600:39]
  wire  _GEN_3656 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3497; // @[lut_35.scala 1589:74 lut_35.scala 1601:39]
  wire  _GEN_3657 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3498; // @[lut_35.scala 1589:74 lut_35.scala 1602:39]
  wire  _GEN_3658 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3499; // @[lut_35.scala 1589:74 lut_35.scala 1603:39]
  wire  _GEN_3659 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3500; // @[lut_35.scala 1589:74 lut_35.scala 1604:39]
  wire  _GEN_3660 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3501; // @[lut_35.scala 1589:74 lut_35.scala 1605:39]
  wire  _GEN_3661 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3502; // @[lut_35.scala 1589:74 lut_35.scala 1606:39]
  wire  _GEN_3662 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3503; // @[lut_35.scala 1589:74 lut_35.scala 1607:39]
  wire  _GEN_3663 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3504; // @[lut_35.scala 1589:74 lut_35.scala 1608:39]
  wire  _GEN_3664 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3505; // @[lut_35.scala 1589:74 lut_35.scala 1609:39]
  wire  _GEN_3665 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3506; // @[lut_35.scala 1589:74 lut_35.scala 1610:39]
  wire  _GEN_3666 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3507; // @[lut_35.scala 1589:74 lut_35.scala 1611:39]
  wire  _GEN_3667 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3508; // @[lut_35.scala 1589:74 lut_35.scala 1612:39]
  wire  _GEN_3668 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3509; // @[lut_35.scala 1589:74 lut_35.scala 1613:39]
  wire  _GEN_3669 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3510; // @[lut_35.scala 1589:74 lut_35.scala 1614:39]
  wire  _GEN_3670 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3511; // @[lut_35.scala 1589:74 lut_35.scala 1615:39]
  wire  _GEN_3671 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3512; // @[lut_35.scala 1589:74 lut_35.scala 1616:39]
  wire  _GEN_3672 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3513; // @[lut_35.scala 1589:74 lut_35.scala 1617:39]
  wire  _GEN_3673 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid | _GEN_3514; // @[lut_35.scala 1589:74 lut_35.scala 1618:39]
  wire  _GEN_3674 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3515; // @[lut_35.scala 1589:74 lut_35.scala 1619:39]
  wire  _GEN_3675 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3516; // @[lut_35.scala 1589:74 lut_35.scala 1620:39]
  wire  _GEN_3676 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3517; // @[lut_35.scala 1589:74 lut_35.scala 1621:39]
  wire  _GEN_3677 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3518; // @[lut_35.scala 1589:74 lut_35.scala 1622:39]
  wire  _GEN_3678 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3519; // @[lut_35.scala 1589:74 lut_35.scala 1623:39]
  wire  _GEN_3679 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3520; // @[lut_35.scala 1589:74 lut_35.scala 1624:39]
  wire  _GEN_3680 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid | _GEN_3521; // @[lut_35.scala 1589:74 lut_35.scala 1625:34]
  wire  _GEN_3684 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1589:74 lut_35.scala 216:26 lut_35.scala 1627:27]
  wire  _GEN_3687 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3525; // @[lut_35.scala 1589:74 lut_35.scala 216:26]
  wire  _GEN_3690 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3528; // @[lut_35.scala 1589:74 lut_35.scala 216:26]
  wire  _GEN_3693 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3531; // @[lut_35.scala 1589:74 lut_35.scala 216:26]
  wire  _GEN_3696 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3534; // @[lut_35.scala 1589:74 lut_35.scala 216:26]
  wire  _GEN_3699 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3537; // @[lut_35.scala 1589:74 lut_35.scala 216:26]
  wire  _GEN_3702 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3540; // @[lut_35.scala 1589:74 lut_35.scala 216:26]
  wire [5:0] _GEN_3703 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? push_mem_temp : _GEN_3541; // @[lut_35.scala 1589:74 lut_35.scala 521:39]
  wire [31:0] _GEN_3704 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? push_id_temp : _GEN_3542; // @[lut_35.scala 1589:74 lut_35.scala 522:39]
  wire  _GEN_3707 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3545; // @[lut_35.scala 1589:74 lut_35.scala 216:26]
  wire  _GEN_3710 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3548; // @[lut_35.scala 1589:74 lut_35.scala 216:26]
  wire  _GEN_3713 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3551; // @[lut_35.scala 1589:74 lut_35.scala 216:26]
  wire  _GEN_3716 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3554; // @[lut_35.scala 1589:74 lut_35.scala 216:26]
  wire  _GEN_3719 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3557; // @[lut_35.scala 1589:74 lut_35.scala 216:26]
  wire  _GEN_3722 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3560; // @[lut_35.scala 1589:74 lut_35.scala 216:26]
  wire  _GEN_3725 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3563; // @[lut_35.scala 1589:74 lut_35.scala 216:26]
  wire  _GEN_3728 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3566; // @[lut_35.scala 1589:74 lut_35.scala 216:26]
  wire  _GEN_3731 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3569; // @[lut_35.scala 1589:74 lut_35.scala 216:26]
  wire  _GEN_3734 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3572; // @[lut_35.scala 1589:74 lut_35.scala 216:26]
  wire  _GEN_3737 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3575; // @[lut_35.scala 1589:74 lut_35.scala 216:26]
  wire  _GEN_3740 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3578; // @[lut_35.scala 1589:74 lut_35.scala 216:26]
  wire  _GEN_3743 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3581; // @[lut_35.scala 1589:74 lut_35.scala 216:26]
  wire  _GEN_3746 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3584; // @[lut_35.scala 1589:74 lut_35.scala 216:26]
  wire  _GEN_3749 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3587; // @[lut_35.scala 1589:74 lut_35.scala 216:26]
  wire  _GEN_3752 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3590; // @[lut_35.scala 1589:74 lut_35.scala 216:26]
  wire  _GEN_3755 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3593; // @[lut_35.scala 1589:74 lut_35.scala 216:26]
  wire  _GEN_3758 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3596; // @[lut_35.scala 1589:74 lut_35.scala 216:26]
  wire  _GEN_3761 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3599; // @[lut_35.scala 1589:74 lut_35.scala 216:26]
  wire  _GEN_3764 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3602; // @[lut_35.scala 1589:74 lut_35.scala 216:26]
  wire  _GEN_3767 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3605; // @[lut_35.scala 1589:74 lut_35.scala 216:26]
  wire  _GEN_3770 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3608; // @[lut_35.scala 1589:74 lut_35.scala 216:26]
  wire  _GEN_3773 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3611; // @[lut_35.scala 1589:74 lut_35.scala 216:26]
  wire  _GEN_3776 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3614; // @[lut_35.scala 1589:74 lut_35.scala 216:26]
  wire  _GEN_3779 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3617; // @[lut_35.scala 1589:74 lut_35.scala 216:26]
  wire  _GEN_3782 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3620; // @[lut_35.scala 1589:74 lut_35.scala 216:26]
  wire  _GEN_3785 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3623; // @[lut_35.scala 1589:74 lut_35.scala 216:26]
  wire  _GEN_3788 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3626; // @[lut_35.scala 1589:74 lut_35.scala 216:26]
  wire  _GEN_3791 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3629; // @[lut_35.scala 1589:74 lut_35.scala 216:26]
  wire  _GEN_3794 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3632; // @[lut_35.scala 1589:74 lut_35.scala 216:26]
  wire  _GEN_3797 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3635; // @[lut_35.scala 1589:74 lut_35.scala 216:26]
  wire  _GEN_3800 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3638; // @[lut_35.scala 1589:74 lut_35.scala 216:26]
  wire  _GEN_3803 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3641; // @[lut_35.scala 1589:74 lut_35.scala 216:26]
  wire  _GEN_3806 = LUT_mem_MPORT_63_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3644; // @[lut_35.scala 1589:74 lut_35.scala 216:26]
  wire  _GEN_3807 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3645; // @[lut_35.scala 1551:74 lut_35.scala 1552:38]
  wire  _GEN_3808 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3646; // @[lut_35.scala 1551:74 lut_35.scala 1553:38]
  wire  _GEN_3809 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3647; // @[lut_35.scala 1551:74 lut_35.scala 1554:38]
  wire  _GEN_3810 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3648; // @[lut_35.scala 1551:74 lut_35.scala 1555:38]
  wire  _GEN_3811 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3649; // @[lut_35.scala 1551:74 lut_35.scala 1556:38]
  wire  _GEN_3812 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3650; // @[lut_35.scala 1551:74 lut_35.scala 1557:38]
  wire  _GEN_3813 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3651; // @[lut_35.scala 1551:74 lut_35.scala 1558:38]
  wire  _GEN_3814 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3652; // @[lut_35.scala 1551:74 lut_35.scala 1559:38]
  wire  _GEN_3815 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3653; // @[lut_35.scala 1551:74 lut_35.scala 1560:38]
  wire  _GEN_3816 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3654; // @[lut_35.scala 1551:74 lut_35.scala 1561:38]
  wire  _GEN_3817 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3655; // @[lut_35.scala 1551:74 lut_35.scala 1562:39]
  wire  _GEN_3818 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3656; // @[lut_35.scala 1551:74 lut_35.scala 1563:39]
  wire  _GEN_3819 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3657; // @[lut_35.scala 1551:74 lut_35.scala 1564:39]
  wire  _GEN_3820 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3658; // @[lut_35.scala 1551:74 lut_35.scala 1565:39]
  wire  _GEN_3821 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3659; // @[lut_35.scala 1551:74 lut_35.scala 1566:39]
  wire  _GEN_3822 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3660; // @[lut_35.scala 1551:74 lut_35.scala 1567:39]
  wire  _GEN_3823 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3661; // @[lut_35.scala 1551:74 lut_35.scala 1568:39]
  wire  _GEN_3824 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3662; // @[lut_35.scala 1551:74 lut_35.scala 1569:39]
  wire  _GEN_3825 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3663; // @[lut_35.scala 1551:74 lut_35.scala 1570:39]
  wire  _GEN_3826 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3664; // @[lut_35.scala 1551:74 lut_35.scala 1571:39]
  wire  _GEN_3827 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3665; // @[lut_35.scala 1551:74 lut_35.scala 1572:39]
  wire  _GEN_3828 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3666; // @[lut_35.scala 1551:74 lut_35.scala 1573:39]
  wire  _GEN_3829 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3667; // @[lut_35.scala 1551:74 lut_35.scala 1574:39]
  wire  _GEN_3830 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3668; // @[lut_35.scala 1551:74 lut_35.scala 1575:39]
  wire  _GEN_3831 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3669; // @[lut_35.scala 1551:74 lut_35.scala 1576:39]
  wire  _GEN_3832 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3670; // @[lut_35.scala 1551:74 lut_35.scala 1577:39]
  wire  _GEN_3833 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3671; // @[lut_35.scala 1551:74 lut_35.scala 1578:39]
  wire  _GEN_3834 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid | _GEN_3672; // @[lut_35.scala 1551:74 lut_35.scala 1579:39]
  wire  _GEN_3835 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3673; // @[lut_35.scala 1551:74 lut_35.scala 1580:39]
  wire  _GEN_3836 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3674; // @[lut_35.scala 1551:74 lut_35.scala 1581:39]
  wire  _GEN_3837 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3675; // @[lut_35.scala 1551:74 lut_35.scala 1582:39]
  wire  _GEN_3838 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3676; // @[lut_35.scala 1551:74 lut_35.scala 1583:39]
  wire  _GEN_3839 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3677; // @[lut_35.scala 1551:74 lut_35.scala 1584:39]
  wire  _GEN_3840 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3678; // @[lut_35.scala 1551:74 lut_35.scala 1585:39]
  wire  _GEN_3841 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3679; // @[lut_35.scala 1551:74 lut_35.scala 1586:39]
  wire  _GEN_3842 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid | _GEN_3680; // @[lut_35.scala 1551:74 lut_35.scala 1587:34]
  wire  _GEN_3846 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1551:74 lut_35.scala 216:26 lut_35.scala 1589:27]
  wire  _GEN_3849 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3684; // @[lut_35.scala 1551:74 lut_35.scala 216:26]
  wire  _GEN_3852 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3687; // @[lut_35.scala 1551:74 lut_35.scala 216:26]
  wire  _GEN_3855 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3690; // @[lut_35.scala 1551:74 lut_35.scala 216:26]
  wire  _GEN_3858 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3693; // @[lut_35.scala 1551:74 lut_35.scala 216:26]
  wire  _GEN_3861 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3696; // @[lut_35.scala 1551:74 lut_35.scala 216:26]
  wire  _GEN_3864 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3699; // @[lut_35.scala 1551:74 lut_35.scala 216:26]
  wire  _GEN_3867 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3702; // @[lut_35.scala 1551:74 lut_35.scala 216:26]
  wire [5:0] _GEN_3868 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? push_mem_temp : _GEN_3703; // @[lut_35.scala 1551:74 lut_35.scala 521:39]
  wire [31:0] _GEN_3869 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? push_id_temp : _GEN_3704; // @[lut_35.scala 1551:74 lut_35.scala 522:39]
  wire  _GEN_3872 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3707; // @[lut_35.scala 1551:74 lut_35.scala 216:26]
  wire  _GEN_3875 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3710; // @[lut_35.scala 1551:74 lut_35.scala 216:26]
  wire  _GEN_3878 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3713; // @[lut_35.scala 1551:74 lut_35.scala 216:26]
  wire  _GEN_3881 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3716; // @[lut_35.scala 1551:74 lut_35.scala 216:26]
  wire  _GEN_3884 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3719; // @[lut_35.scala 1551:74 lut_35.scala 216:26]
  wire  _GEN_3887 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3722; // @[lut_35.scala 1551:74 lut_35.scala 216:26]
  wire  _GEN_3890 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3725; // @[lut_35.scala 1551:74 lut_35.scala 216:26]
  wire  _GEN_3893 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3728; // @[lut_35.scala 1551:74 lut_35.scala 216:26]
  wire  _GEN_3896 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3731; // @[lut_35.scala 1551:74 lut_35.scala 216:26]
  wire  _GEN_3899 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3734; // @[lut_35.scala 1551:74 lut_35.scala 216:26]
  wire  _GEN_3902 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3737; // @[lut_35.scala 1551:74 lut_35.scala 216:26]
  wire  _GEN_3905 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3740; // @[lut_35.scala 1551:74 lut_35.scala 216:26]
  wire  _GEN_3908 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3743; // @[lut_35.scala 1551:74 lut_35.scala 216:26]
  wire  _GEN_3911 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3746; // @[lut_35.scala 1551:74 lut_35.scala 216:26]
  wire  _GEN_3914 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3749; // @[lut_35.scala 1551:74 lut_35.scala 216:26]
  wire  _GEN_3917 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3752; // @[lut_35.scala 1551:74 lut_35.scala 216:26]
  wire  _GEN_3920 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3755; // @[lut_35.scala 1551:74 lut_35.scala 216:26]
  wire  _GEN_3923 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3758; // @[lut_35.scala 1551:74 lut_35.scala 216:26]
  wire  _GEN_3926 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3761; // @[lut_35.scala 1551:74 lut_35.scala 216:26]
  wire  _GEN_3929 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3764; // @[lut_35.scala 1551:74 lut_35.scala 216:26]
  wire  _GEN_3932 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3767; // @[lut_35.scala 1551:74 lut_35.scala 216:26]
  wire  _GEN_3935 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3770; // @[lut_35.scala 1551:74 lut_35.scala 216:26]
  wire  _GEN_3938 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3773; // @[lut_35.scala 1551:74 lut_35.scala 216:26]
  wire  _GEN_3941 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3776; // @[lut_35.scala 1551:74 lut_35.scala 216:26]
  wire  _GEN_3944 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3779; // @[lut_35.scala 1551:74 lut_35.scala 216:26]
  wire  _GEN_3947 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3782; // @[lut_35.scala 1551:74 lut_35.scala 216:26]
  wire  _GEN_3950 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3785; // @[lut_35.scala 1551:74 lut_35.scala 216:26]
  wire  _GEN_3953 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3788; // @[lut_35.scala 1551:74 lut_35.scala 216:26]
  wire  _GEN_3956 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3791; // @[lut_35.scala 1551:74 lut_35.scala 216:26]
  wire  _GEN_3959 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3794; // @[lut_35.scala 1551:74 lut_35.scala 216:26]
  wire  _GEN_3962 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3797; // @[lut_35.scala 1551:74 lut_35.scala 216:26]
  wire  _GEN_3965 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3800; // @[lut_35.scala 1551:74 lut_35.scala 216:26]
  wire  _GEN_3968 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3803; // @[lut_35.scala 1551:74 lut_35.scala 216:26]
  wire  _GEN_3971 = LUT_mem_MPORT_62_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3806; // @[lut_35.scala 1551:74 lut_35.scala 216:26]
  wire  _GEN_3972 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3807; // @[lut_35.scala 1513:74 lut_35.scala 1514:38]
  wire  _GEN_3973 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3808; // @[lut_35.scala 1513:74 lut_35.scala 1515:38]
  wire  _GEN_3974 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3809; // @[lut_35.scala 1513:74 lut_35.scala 1516:38]
  wire  _GEN_3975 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3810; // @[lut_35.scala 1513:74 lut_35.scala 1517:38]
  wire  _GEN_3976 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3811; // @[lut_35.scala 1513:74 lut_35.scala 1518:38]
  wire  _GEN_3977 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3812; // @[lut_35.scala 1513:74 lut_35.scala 1519:38]
  wire  _GEN_3978 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3813; // @[lut_35.scala 1513:74 lut_35.scala 1520:38]
  wire  _GEN_3979 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3814; // @[lut_35.scala 1513:74 lut_35.scala 1521:38]
  wire  _GEN_3980 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3815; // @[lut_35.scala 1513:74 lut_35.scala 1522:38]
  wire  _GEN_3981 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3816; // @[lut_35.scala 1513:74 lut_35.scala 1523:38]
  wire  _GEN_3982 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3817; // @[lut_35.scala 1513:74 lut_35.scala 1524:39]
  wire  _GEN_3983 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3818; // @[lut_35.scala 1513:74 lut_35.scala 1525:39]
  wire  _GEN_3984 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3819; // @[lut_35.scala 1513:74 lut_35.scala 1526:39]
  wire  _GEN_3985 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3820; // @[lut_35.scala 1513:74 lut_35.scala 1527:39]
  wire  _GEN_3986 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3821; // @[lut_35.scala 1513:74 lut_35.scala 1528:39]
  wire  _GEN_3987 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3822; // @[lut_35.scala 1513:74 lut_35.scala 1529:39]
  wire  _GEN_3988 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3823; // @[lut_35.scala 1513:74 lut_35.scala 1530:39]
  wire  _GEN_3989 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3824; // @[lut_35.scala 1513:74 lut_35.scala 1531:39]
  wire  _GEN_3990 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3825; // @[lut_35.scala 1513:74 lut_35.scala 1532:39]
  wire  _GEN_3991 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3826; // @[lut_35.scala 1513:74 lut_35.scala 1533:39]
  wire  _GEN_3992 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3827; // @[lut_35.scala 1513:74 lut_35.scala 1534:39]
  wire  _GEN_3993 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3828; // @[lut_35.scala 1513:74 lut_35.scala 1535:39]
  wire  _GEN_3994 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3829; // @[lut_35.scala 1513:74 lut_35.scala 1536:39]
  wire  _GEN_3995 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3830; // @[lut_35.scala 1513:74 lut_35.scala 1537:39]
  wire  _GEN_3996 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3831; // @[lut_35.scala 1513:74 lut_35.scala 1538:39]
  wire  _GEN_3997 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3832; // @[lut_35.scala 1513:74 lut_35.scala 1539:39]
  wire  _GEN_3998 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid | _GEN_3833; // @[lut_35.scala 1513:74 lut_35.scala 1540:39]
  wire  _GEN_3999 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3834; // @[lut_35.scala 1513:74 lut_35.scala 1541:39]
  wire  _GEN_4000 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3835; // @[lut_35.scala 1513:74 lut_35.scala 1542:39]
  wire  _GEN_4001 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3836; // @[lut_35.scala 1513:74 lut_35.scala 1543:39]
  wire  _GEN_4002 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3837; // @[lut_35.scala 1513:74 lut_35.scala 1544:39]
  wire  _GEN_4003 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3838; // @[lut_35.scala 1513:74 lut_35.scala 1545:39]
  wire  _GEN_4004 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3839; // @[lut_35.scala 1513:74 lut_35.scala 1546:39]
  wire  _GEN_4005 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3840; // @[lut_35.scala 1513:74 lut_35.scala 1547:39]
  wire  _GEN_4006 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3841; // @[lut_35.scala 1513:74 lut_35.scala 1548:39]
  wire  _GEN_4007 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid | _GEN_3842; // @[lut_35.scala 1513:74 lut_35.scala 1549:34]
  wire  _GEN_4011 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1513:74 lut_35.scala 216:26 lut_35.scala 1551:27]
  wire  _GEN_4014 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3846; // @[lut_35.scala 1513:74 lut_35.scala 216:26]
  wire  _GEN_4017 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3849; // @[lut_35.scala 1513:74 lut_35.scala 216:26]
  wire  _GEN_4020 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3852; // @[lut_35.scala 1513:74 lut_35.scala 216:26]
  wire  _GEN_4023 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3855; // @[lut_35.scala 1513:74 lut_35.scala 216:26]
  wire  _GEN_4026 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3858; // @[lut_35.scala 1513:74 lut_35.scala 216:26]
  wire  _GEN_4029 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3861; // @[lut_35.scala 1513:74 lut_35.scala 216:26]
  wire  _GEN_4032 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3864; // @[lut_35.scala 1513:74 lut_35.scala 216:26]
  wire  _GEN_4035 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3867; // @[lut_35.scala 1513:74 lut_35.scala 216:26]
  wire [5:0] _GEN_4036 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? push_mem_temp : _GEN_3868; // @[lut_35.scala 1513:74 lut_35.scala 521:39]
  wire [31:0] _GEN_4037 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? push_id_temp : _GEN_3869; // @[lut_35.scala 1513:74 lut_35.scala 522:39]
  wire  _GEN_4040 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3872; // @[lut_35.scala 1513:74 lut_35.scala 216:26]
  wire  _GEN_4043 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3875; // @[lut_35.scala 1513:74 lut_35.scala 216:26]
  wire  _GEN_4046 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3878; // @[lut_35.scala 1513:74 lut_35.scala 216:26]
  wire  _GEN_4049 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3881; // @[lut_35.scala 1513:74 lut_35.scala 216:26]
  wire  _GEN_4052 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3884; // @[lut_35.scala 1513:74 lut_35.scala 216:26]
  wire  _GEN_4055 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3887; // @[lut_35.scala 1513:74 lut_35.scala 216:26]
  wire  _GEN_4058 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3890; // @[lut_35.scala 1513:74 lut_35.scala 216:26]
  wire  _GEN_4061 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3893; // @[lut_35.scala 1513:74 lut_35.scala 216:26]
  wire  _GEN_4064 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3896; // @[lut_35.scala 1513:74 lut_35.scala 216:26]
  wire  _GEN_4067 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3899; // @[lut_35.scala 1513:74 lut_35.scala 216:26]
  wire  _GEN_4070 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3902; // @[lut_35.scala 1513:74 lut_35.scala 216:26]
  wire  _GEN_4073 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3905; // @[lut_35.scala 1513:74 lut_35.scala 216:26]
  wire  _GEN_4076 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3908; // @[lut_35.scala 1513:74 lut_35.scala 216:26]
  wire  _GEN_4079 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3911; // @[lut_35.scala 1513:74 lut_35.scala 216:26]
  wire  _GEN_4082 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3914; // @[lut_35.scala 1513:74 lut_35.scala 216:26]
  wire  _GEN_4085 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3917; // @[lut_35.scala 1513:74 lut_35.scala 216:26]
  wire  _GEN_4088 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3920; // @[lut_35.scala 1513:74 lut_35.scala 216:26]
  wire  _GEN_4091 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3923; // @[lut_35.scala 1513:74 lut_35.scala 216:26]
  wire  _GEN_4094 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3926; // @[lut_35.scala 1513:74 lut_35.scala 216:26]
  wire  _GEN_4097 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3929; // @[lut_35.scala 1513:74 lut_35.scala 216:26]
  wire  _GEN_4100 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3932; // @[lut_35.scala 1513:74 lut_35.scala 216:26]
  wire  _GEN_4103 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3935; // @[lut_35.scala 1513:74 lut_35.scala 216:26]
  wire  _GEN_4106 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3938; // @[lut_35.scala 1513:74 lut_35.scala 216:26]
  wire  _GEN_4109 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3941; // @[lut_35.scala 1513:74 lut_35.scala 216:26]
  wire  _GEN_4112 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3944; // @[lut_35.scala 1513:74 lut_35.scala 216:26]
  wire  _GEN_4115 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3947; // @[lut_35.scala 1513:74 lut_35.scala 216:26]
  wire  _GEN_4118 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3950; // @[lut_35.scala 1513:74 lut_35.scala 216:26]
  wire  _GEN_4121 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3953; // @[lut_35.scala 1513:74 lut_35.scala 216:26]
  wire  _GEN_4124 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3956; // @[lut_35.scala 1513:74 lut_35.scala 216:26]
  wire  _GEN_4127 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3959; // @[lut_35.scala 1513:74 lut_35.scala 216:26]
  wire  _GEN_4130 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3962; // @[lut_35.scala 1513:74 lut_35.scala 216:26]
  wire  _GEN_4133 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3965; // @[lut_35.scala 1513:74 lut_35.scala 216:26]
  wire  _GEN_4136 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3968; // @[lut_35.scala 1513:74 lut_35.scala 216:26]
  wire  _GEN_4139 = LUT_mem_MPORT_61_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3971; // @[lut_35.scala 1513:74 lut_35.scala 216:26]
  wire  _GEN_4140 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3972; // @[lut_35.scala 1475:74 lut_35.scala 1476:38]
  wire  _GEN_4141 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3973; // @[lut_35.scala 1475:74 lut_35.scala 1477:38]
  wire  _GEN_4142 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3974; // @[lut_35.scala 1475:74 lut_35.scala 1478:38]
  wire  _GEN_4143 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3975; // @[lut_35.scala 1475:74 lut_35.scala 1479:38]
  wire  _GEN_4144 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3976; // @[lut_35.scala 1475:74 lut_35.scala 1480:38]
  wire  _GEN_4145 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3977; // @[lut_35.scala 1475:74 lut_35.scala 1481:38]
  wire  _GEN_4146 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3978; // @[lut_35.scala 1475:74 lut_35.scala 1482:38]
  wire  _GEN_4147 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3979; // @[lut_35.scala 1475:74 lut_35.scala 1483:38]
  wire  _GEN_4148 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3980; // @[lut_35.scala 1475:74 lut_35.scala 1484:38]
  wire  _GEN_4149 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3981; // @[lut_35.scala 1475:74 lut_35.scala 1485:38]
  wire  _GEN_4150 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3982; // @[lut_35.scala 1475:74 lut_35.scala 1486:39]
  wire  _GEN_4151 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3983; // @[lut_35.scala 1475:74 lut_35.scala 1487:39]
  wire  _GEN_4152 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3984; // @[lut_35.scala 1475:74 lut_35.scala 1488:39]
  wire  _GEN_4153 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3985; // @[lut_35.scala 1475:74 lut_35.scala 1489:39]
  wire  _GEN_4154 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3986; // @[lut_35.scala 1475:74 lut_35.scala 1490:39]
  wire  _GEN_4155 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3987; // @[lut_35.scala 1475:74 lut_35.scala 1491:39]
  wire  _GEN_4156 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3988; // @[lut_35.scala 1475:74 lut_35.scala 1492:39]
  wire  _GEN_4157 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3989; // @[lut_35.scala 1475:74 lut_35.scala 1493:39]
  wire  _GEN_4158 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3990; // @[lut_35.scala 1475:74 lut_35.scala 1494:39]
  wire  _GEN_4159 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3991; // @[lut_35.scala 1475:74 lut_35.scala 1495:39]
  wire  _GEN_4160 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3992; // @[lut_35.scala 1475:74 lut_35.scala 1496:39]
  wire  _GEN_4161 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3993; // @[lut_35.scala 1475:74 lut_35.scala 1497:39]
  wire  _GEN_4162 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3994; // @[lut_35.scala 1475:74 lut_35.scala 1498:39]
  wire  _GEN_4163 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3995; // @[lut_35.scala 1475:74 lut_35.scala 1499:39]
  wire  _GEN_4164 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3996; // @[lut_35.scala 1475:74 lut_35.scala 1500:39]
  wire  _GEN_4165 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid | _GEN_3997; // @[lut_35.scala 1475:74 lut_35.scala 1501:39]
  wire  _GEN_4166 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3998; // @[lut_35.scala 1475:74 lut_35.scala 1502:39]
  wire  _GEN_4167 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_3999; // @[lut_35.scala 1475:74 lut_35.scala 1503:39]
  wire  _GEN_4168 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4000; // @[lut_35.scala 1475:74 lut_35.scala 1504:39]
  wire  _GEN_4169 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4001; // @[lut_35.scala 1475:74 lut_35.scala 1505:39]
  wire  _GEN_4170 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4002; // @[lut_35.scala 1475:74 lut_35.scala 1506:39]
  wire  _GEN_4171 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4003; // @[lut_35.scala 1475:74 lut_35.scala 1507:39]
  wire  _GEN_4172 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4004; // @[lut_35.scala 1475:74 lut_35.scala 1508:39]
  wire  _GEN_4173 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4005; // @[lut_35.scala 1475:74 lut_35.scala 1509:39]
  wire  _GEN_4174 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4006; // @[lut_35.scala 1475:74 lut_35.scala 1510:39]
  wire  _GEN_4175 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid | _GEN_4007; // @[lut_35.scala 1475:74 lut_35.scala 1511:34]
  wire  _GEN_4179 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1475:74 lut_35.scala 216:26 lut_35.scala 1513:27]
  wire  _GEN_4182 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4011; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire  _GEN_4185 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4014; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire  _GEN_4188 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4017; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire  _GEN_4191 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4020; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire  _GEN_4194 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4023; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire  _GEN_4197 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4026; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire  _GEN_4200 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4029; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire  _GEN_4203 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4032; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire  _GEN_4206 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4035; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire [5:0] _GEN_4207 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? push_mem_temp : _GEN_4036; // @[lut_35.scala 1475:74 lut_35.scala 521:39]
  wire [31:0] _GEN_4208 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? push_id_temp : _GEN_4037; // @[lut_35.scala 1475:74 lut_35.scala 522:39]
  wire  _GEN_4211 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4040; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire  _GEN_4214 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4043; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire  _GEN_4217 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4046; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire  _GEN_4220 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4049; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire  _GEN_4223 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4052; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire  _GEN_4226 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4055; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire  _GEN_4229 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4058; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire  _GEN_4232 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4061; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire  _GEN_4235 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4064; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire  _GEN_4238 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4067; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire  _GEN_4241 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4070; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire  _GEN_4244 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4073; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire  _GEN_4247 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4076; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire  _GEN_4250 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4079; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire  _GEN_4253 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4082; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire  _GEN_4256 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4085; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire  _GEN_4259 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4088; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire  _GEN_4262 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4091; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire  _GEN_4265 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4094; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire  _GEN_4268 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4097; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire  _GEN_4271 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4100; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire  _GEN_4274 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4103; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire  _GEN_4277 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4106; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire  _GEN_4280 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4109; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire  _GEN_4283 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4112; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire  _GEN_4286 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4115; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire  _GEN_4289 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4118; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire  _GEN_4292 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4121; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire  _GEN_4295 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4124; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire  _GEN_4298 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4127; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire  _GEN_4301 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4130; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire  _GEN_4304 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4133; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire  _GEN_4307 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4136; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire  _GEN_4310 = LUT_mem_MPORT_60_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4139; // @[lut_35.scala 1475:74 lut_35.scala 216:26]
  wire  _GEN_4311 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4140; // @[lut_35.scala 1437:74 lut_35.scala 1438:38]
  wire  _GEN_4312 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4141; // @[lut_35.scala 1437:74 lut_35.scala 1439:38]
  wire  _GEN_4313 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4142; // @[lut_35.scala 1437:74 lut_35.scala 1440:38]
  wire  _GEN_4314 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4143; // @[lut_35.scala 1437:74 lut_35.scala 1441:38]
  wire  _GEN_4315 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4144; // @[lut_35.scala 1437:74 lut_35.scala 1442:38]
  wire  _GEN_4316 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4145; // @[lut_35.scala 1437:74 lut_35.scala 1443:38]
  wire  _GEN_4317 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4146; // @[lut_35.scala 1437:74 lut_35.scala 1444:38]
  wire  _GEN_4318 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4147; // @[lut_35.scala 1437:74 lut_35.scala 1445:38]
  wire  _GEN_4319 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4148; // @[lut_35.scala 1437:74 lut_35.scala 1446:38]
  wire  _GEN_4320 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4149; // @[lut_35.scala 1437:74 lut_35.scala 1447:38]
  wire  _GEN_4321 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4150; // @[lut_35.scala 1437:74 lut_35.scala 1448:39]
  wire  _GEN_4322 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4151; // @[lut_35.scala 1437:74 lut_35.scala 1449:39]
  wire  _GEN_4323 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4152; // @[lut_35.scala 1437:74 lut_35.scala 1450:39]
  wire  _GEN_4324 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4153; // @[lut_35.scala 1437:74 lut_35.scala 1451:39]
  wire  _GEN_4325 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4154; // @[lut_35.scala 1437:74 lut_35.scala 1452:39]
  wire  _GEN_4326 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4155; // @[lut_35.scala 1437:74 lut_35.scala 1453:39]
  wire  _GEN_4327 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4156; // @[lut_35.scala 1437:74 lut_35.scala 1454:39]
  wire  _GEN_4328 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4157; // @[lut_35.scala 1437:74 lut_35.scala 1455:39]
  wire  _GEN_4329 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4158; // @[lut_35.scala 1437:74 lut_35.scala 1456:39]
  wire  _GEN_4330 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4159; // @[lut_35.scala 1437:74 lut_35.scala 1457:39]
  wire  _GEN_4331 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4160; // @[lut_35.scala 1437:74 lut_35.scala 1458:39]
  wire  _GEN_4332 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4161; // @[lut_35.scala 1437:74 lut_35.scala 1459:39]
  wire  _GEN_4333 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4162; // @[lut_35.scala 1437:74 lut_35.scala 1460:39]
  wire  _GEN_4334 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4163; // @[lut_35.scala 1437:74 lut_35.scala 1461:39]
  wire  _GEN_4335 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid | _GEN_4164; // @[lut_35.scala 1437:74 lut_35.scala 1462:39]
  wire  _GEN_4336 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4165; // @[lut_35.scala 1437:74 lut_35.scala 1463:39]
  wire  _GEN_4337 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4166; // @[lut_35.scala 1437:74 lut_35.scala 1464:39]
  wire  _GEN_4338 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4167; // @[lut_35.scala 1437:74 lut_35.scala 1465:39]
  wire  _GEN_4339 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4168; // @[lut_35.scala 1437:74 lut_35.scala 1466:39]
  wire  _GEN_4340 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4169; // @[lut_35.scala 1437:74 lut_35.scala 1467:39]
  wire  _GEN_4341 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4170; // @[lut_35.scala 1437:74 lut_35.scala 1468:39]
  wire  _GEN_4342 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4171; // @[lut_35.scala 1437:74 lut_35.scala 1469:39]
  wire  _GEN_4343 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4172; // @[lut_35.scala 1437:74 lut_35.scala 1470:39]
  wire  _GEN_4344 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4173; // @[lut_35.scala 1437:74 lut_35.scala 1471:39]
  wire  _GEN_4345 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4174; // @[lut_35.scala 1437:74 lut_35.scala 1472:39]
  wire  _GEN_4346 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid | _GEN_4175; // @[lut_35.scala 1437:74 lut_35.scala 1473:34]
  wire  _GEN_4350 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1437:74 lut_35.scala 216:26 lut_35.scala 1475:27]
  wire  _GEN_4353 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4179; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4356 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4182; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4359 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4185; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4362 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4188; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4365 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4191; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4368 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4194; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4371 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4197; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4374 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4200; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4377 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4203; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4380 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4206; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire [5:0] _GEN_4381 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? push_mem_temp : _GEN_4207; // @[lut_35.scala 1437:74 lut_35.scala 521:39]
  wire [31:0] _GEN_4382 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? push_id_temp : _GEN_4208; // @[lut_35.scala 1437:74 lut_35.scala 522:39]
  wire  _GEN_4385 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4211; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4388 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4214; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4391 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4217; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4394 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4220; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4397 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4223; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4400 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4226; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4403 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4229; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4406 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4232; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4409 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4235; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4412 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4238; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4415 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4241; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4418 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4244; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4421 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4247; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4424 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4250; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4427 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4253; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4430 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4256; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4433 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4259; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4436 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4262; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4439 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4265; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4442 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4268; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4445 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4271; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4448 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4274; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4451 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4277; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4454 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4280; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4457 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4283; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4460 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4286; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4463 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4289; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4466 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4292; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4469 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4295; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4472 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4298; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4475 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4301; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4478 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4304; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4481 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4307; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4484 = LUT_mem_MPORT_59_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4310; // @[lut_35.scala 1437:74 lut_35.scala 216:26]
  wire  _GEN_4485 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4311; // @[lut_35.scala 1399:74 lut_35.scala 1400:38]
  wire  _GEN_4486 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4312; // @[lut_35.scala 1399:74 lut_35.scala 1401:38]
  wire  _GEN_4487 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4313; // @[lut_35.scala 1399:74 lut_35.scala 1402:38]
  wire  _GEN_4488 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4314; // @[lut_35.scala 1399:74 lut_35.scala 1403:38]
  wire  _GEN_4489 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4315; // @[lut_35.scala 1399:74 lut_35.scala 1404:38]
  wire  _GEN_4490 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4316; // @[lut_35.scala 1399:74 lut_35.scala 1405:38]
  wire  _GEN_4491 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4317; // @[lut_35.scala 1399:74 lut_35.scala 1406:38]
  wire  _GEN_4492 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4318; // @[lut_35.scala 1399:74 lut_35.scala 1407:38]
  wire  _GEN_4493 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4319; // @[lut_35.scala 1399:74 lut_35.scala 1408:38]
  wire  _GEN_4494 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4320; // @[lut_35.scala 1399:74 lut_35.scala 1409:38]
  wire  _GEN_4495 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4321; // @[lut_35.scala 1399:74 lut_35.scala 1410:39]
  wire  _GEN_4496 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4322; // @[lut_35.scala 1399:74 lut_35.scala 1411:39]
  wire  _GEN_4497 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4323; // @[lut_35.scala 1399:74 lut_35.scala 1412:39]
  wire  _GEN_4498 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4324; // @[lut_35.scala 1399:74 lut_35.scala 1413:39]
  wire  _GEN_4499 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4325; // @[lut_35.scala 1399:74 lut_35.scala 1414:39]
  wire  _GEN_4500 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4326; // @[lut_35.scala 1399:74 lut_35.scala 1415:39]
  wire  _GEN_4501 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4327; // @[lut_35.scala 1399:74 lut_35.scala 1416:39]
  wire  _GEN_4502 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4328; // @[lut_35.scala 1399:74 lut_35.scala 1417:39]
  wire  _GEN_4503 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4329; // @[lut_35.scala 1399:74 lut_35.scala 1418:39]
  wire  _GEN_4504 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4330; // @[lut_35.scala 1399:74 lut_35.scala 1419:39]
  wire  _GEN_4505 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4331; // @[lut_35.scala 1399:74 lut_35.scala 1420:39]
  wire  _GEN_4506 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4332; // @[lut_35.scala 1399:74 lut_35.scala 1421:39]
  wire  _GEN_4507 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4333; // @[lut_35.scala 1399:74 lut_35.scala 1422:39]
  wire  _GEN_4508 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid | _GEN_4334; // @[lut_35.scala 1399:74 lut_35.scala 1423:39]
  wire  _GEN_4509 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4335; // @[lut_35.scala 1399:74 lut_35.scala 1424:39]
  wire  _GEN_4510 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4336; // @[lut_35.scala 1399:74 lut_35.scala 1425:39]
  wire  _GEN_4511 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4337; // @[lut_35.scala 1399:74 lut_35.scala 1426:39]
  wire  _GEN_4512 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4338; // @[lut_35.scala 1399:74 lut_35.scala 1427:39]
  wire  _GEN_4513 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4339; // @[lut_35.scala 1399:74 lut_35.scala 1428:39]
  wire  _GEN_4514 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4340; // @[lut_35.scala 1399:74 lut_35.scala 1429:39]
  wire  _GEN_4515 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4341; // @[lut_35.scala 1399:74 lut_35.scala 1430:39]
  wire  _GEN_4516 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4342; // @[lut_35.scala 1399:74 lut_35.scala 1431:39]
  wire  _GEN_4517 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4343; // @[lut_35.scala 1399:74 lut_35.scala 1432:39]
  wire  _GEN_4518 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4344; // @[lut_35.scala 1399:74 lut_35.scala 1433:39]
  wire  _GEN_4519 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4345; // @[lut_35.scala 1399:74 lut_35.scala 1434:39]
  wire  _GEN_4520 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid | _GEN_4346; // @[lut_35.scala 1399:74 lut_35.scala 1435:34]
  wire  _GEN_4524 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1399:74 lut_35.scala 216:26 lut_35.scala 1437:27]
  wire  _GEN_4527 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4350; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4530 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4353; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4533 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4356; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4536 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4359; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4539 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4362; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4542 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4365; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4545 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4368; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4548 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4371; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4551 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4374; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4554 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4377; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4557 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4380; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire [5:0] _GEN_4558 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? push_mem_temp : _GEN_4381; // @[lut_35.scala 1399:74 lut_35.scala 521:39]
  wire [31:0] _GEN_4559 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? push_id_temp : _GEN_4382; // @[lut_35.scala 1399:74 lut_35.scala 522:39]
  wire  _GEN_4562 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4385; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4565 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4388; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4568 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4391; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4571 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4394; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4574 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4397; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4577 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4400; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4580 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4403; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4583 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4406; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4586 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4409; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4589 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4412; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4592 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4415; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4595 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4418; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4598 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4421; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4601 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4424; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4604 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4427; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4607 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4430; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4610 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4433; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4613 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4436; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4616 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4439; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4619 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4442; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4622 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4445; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4625 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4448; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4628 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4451; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4631 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4454; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4634 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4457; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4637 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4460; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4640 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4463; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4643 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4466; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4646 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4469; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4649 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4472; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4652 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4475; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4655 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4478; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4658 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4481; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4661 = LUT_mem_MPORT_58_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4484; // @[lut_35.scala 1399:74 lut_35.scala 216:26]
  wire  _GEN_4662 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4485; // @[lut_35.scala 1361:75 lut_35.scala 1362:38]
  wire  _GEN_4663 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4486; // @[lut_35.scala 1361:75 lut_35.scala 1363:38]
  wire  _GEN_4664 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4487; // @[lut_35.scala 1361:75 lut_35.scala 1364:38]
  wire  _GEN_4665 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4488; // @[lut_35.scala 1361:75 lut_35.scala 1365:38]
  wire  _GEN_4666 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4489; // @[lut_35.scala 1361:75 lut_35.scala 1366:38]
  wire  _GEN_4667 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4490; // @[lut_35.scala 1361:75 lut_35.scala 1367:38]
  wire  _GEN_4668 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4491; // @[lut_35.scala 1361:75 lut_35.scala 1368:38]
  wire  _GEN_4669 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4492; // @[lut_35.scala 1361:75 lut_35.scala 1369:38]
  wire  _GEN_4670 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4493; // @[lut_35.scala 1361:75 lut_35.scala 1370:38]
  wire  _GEN_4671 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4494; // @[lut_35.scala 1361:75 lut_35.scala 1371:38]
  wire  _GEN_4672 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4495; // @[lut_35.scala 1361:75 lut_35.scala 1372:39]
  wire  _GEN_4673 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4496; // @[lut_35.scala 1361:75 lut_35.scala 1373:39]
  wire  _GEN_4674 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4497; // @[lut_35.scala 1361:75 lut_35.scala 1374:39]
  wire  _GEN_4675 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4498; // @[lut_35.scala 1361:75 lut_35.scala 1375:39]
  wire  _GEN_4676 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4499; // @[lut_35.scala 1361:75 lut_35.scala 1376:39]
  wire  _GEN_4677 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4500; // @[lut_35.scala 1361:75 lut_35.scala 1377:39]
  wire  _GEN_4678 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4501; // @[lut_35.scala 1361:75 lut_35.scala 1378:39]
  wire  _GEN_4679 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4502; // @[lut_35.scala 1361:75 lut_35.scala 1379:39]
  wire  _GEN_4680 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4503; // @[lut_35.scala 1361:75 lut_35.scala 1380:39]
  wire  _GEN_4681 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4504; // @[lut_35.scala 1361:75 lut_35.scala 1381:39]
  wire  _GEN_4682 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4505; // @[lut_35.scala 1361:75 lut_35.scala 1382:39]
  wire  _GEN_4683 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4506; // @[lut_35.scala 1361:75 lut_35.scala 1383:39]
  wire  _GEN_4684 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid | _GEN_4507; // @[lut_35.scala 1361:75 lut_35.scala 1384:39]
  wire  _GEN_4685 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4508; // @[lut_35.scala 1361:75 lut_35.scala 1385:39]
  wire  _GEN_4686 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4509; // @[lut_35.scala 1361:75 lut_35.scala 1386:39]
  wire  _GEN_4687 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4510; // @[lut_35.scala 1361:75 lut_35.scala 1387:39]
  wire  _GEN_4688 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4511; // @[lut_35.scala 1361:75 lut_35.scala 1388:39]
  wire  _GEN_4689 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4512; // @[lut_35.scala 1361:75 lut_35.scala 1389:39]
  wire  _GEN_4690 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4513; // @[lut_35.scala 1361:75 lut_35.scala 1390:39]
  wire  _GEN_4691 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4514; // @[lut_35.scala 1361:75 lut_35.scala 1391:39]
  wire  _GEN_4692 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4515; // @[lut_35.scala 1361:75 lut_35.scala 1392:39]
  wire  _GEN_4693 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4516; // @[lut_35.scala 1361:75 lut_35.scala 1393:39]
  wire  _GEN_4694 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4517; // @[lut_35.scala 1361:75 lut_35.scala 1394:39]
  wire  _GEN_4695 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4518; // @[lut_35.scala 1361:75 lut_35.scala 1395:39]
  wire  _GEN_4696 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4519; // @[lut_35.scala 1361:75 lut_35.scala 1396:39]
  wire  _GEN_4697 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid | _GEN_4520; // @[lut_35.scala 1361:75 lut_35.scala 1397:34]
  wire  _GEN_4701 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1361:75 lut_35.scala 216:26 lut_35.scala 1399:27]
  wire  _GEN_4704 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4524; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4707 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4527; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4710 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4530; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4713 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4533; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4716 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4536; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4719 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4539; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4722 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4542; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4725 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4545; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4728 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4548; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4731 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4551; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4734 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4554; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4737 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4557; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire [5:0] _GEN_4738 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? push_mem_temp : _GEN_4558; // @[lut_35.scala 1361:75 lut_35.scala 521:39]
  wire [31:0] _GEN_4739 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? push_id_temp : _GEN_4559; // @[lut_35.scala 1361:75 lut_35.scala 522:39]
  wire  _GEN_4742 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4562; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4745 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4565; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4748 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4568; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4751 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4571; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4754 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4574; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4757 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4577; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4760 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4580; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4763 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4583; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4766 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4586; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4769 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4589; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4772 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4592; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4775 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4595; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4778 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4598; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4781 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4601; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4784 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4604; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4787 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4607; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4790 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4610; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4793 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4613; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4796 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4616; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4799 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4619; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4802 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4622; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4805 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4625; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4808 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4628; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4811 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4631; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4814 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4634; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4817 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4637; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4820 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4640; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4823 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4643; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4826 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4646; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4829 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4649; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4832 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4652; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4835 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4655; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4838 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4658; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4841 = LUT_mem_MPORT_57_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4661; // @[lut_35.scala 1361:75 lut_35.scala 216:26]
  wire  _GEN_4842 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4662; // @[lut_35.scala 1323:74 lut_35.scala 1324:38]
  wire  _GEN_4843 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4663; // @[lut_35.scala 1323:74 lut_35.scala 1325:38]
  wire  _GEN_4844 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4664; // @[lut_35.scala 1323:74 lut_35.scala 1326:38]
  wire  _GEN_4845 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4665; // @[lut_35.scala 1323:74 lut_35.scala 1327:38]
  wire  _GEN_4846 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4666; // @[lut_35.scala 1323:74 lut_35.scala 1328:38]
  wire  _GEN_4847 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4667; // @[lut_35.scala 1323:74 lut_35.scala 1329:38]
  wire  _GEN_4848 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4668; // @[lut_35.scala 1323:74 lut_35.scala 1330:38]
  wire  _GEN_4849 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4669; // @[lut_35.scala 1323:74 lut_35.scala 1331:38]
  wire  _GEN_4850 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4670; // @[lut_35.scala 1323:74 lut_35.scala 1332:38]
  wire  _GEN_4851 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4671; // @[lut_35.scala 1323:74 lut_35.scala 1333:38]
  wire  _GEN_4852 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4672; // @[lut_35.scala 1323:74 lut_35.scala 1334:39]
  wire  _GEN_4853 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4673; // @[lut_35.scala 1323:74 lut_35.scala 1335:39]
  wire  _GEN_4854 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4674; // @[lut_35.scala 1323:74 lut_35.scala 1336:39]
  wire  _GEN_4855 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4675; // @[lut_35.scala 1323:74 lut_35.scala 1337:39]
  wire  _GEN_4856 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4676; // @[lut_35.scala 1323:74 lut_35.scala 1338:39]
  wire  _GEN_4857 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4677; // @[lut_35.scala 1323:74 lut_35.scala 1339:39]
  wire  _GEN_4858 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4678; // @[lut_35.scala 1323:74 lut_35.scala 1340:39]
  wire  _GEN_4859 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4679; // @[lut_35.scala 1323:74 lut_35.scala 1341:39]
  wire  _GEN_4860 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4680; // @[lut_35.scala 1323:74 lut_35.scala 1342:39]
  wire  _GEN_4861 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4681; // @[lut_35.scala 1323:74 lut_35.scala 1343:39]
  wire  _GEN_4862 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4682; // @[lut_35.scala 1323:74 lut_35.scala 1344:39]
  wire  _GEN_4863 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid | _GEN_4683; // @[lut_35.scala 1323:74 lut_35.scala 1345:39]
  wire  _GEN_4864 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4684; // @[lut_35.scala 1323:74 lut_35.scala 1346:39]
  wire  _GEN_4865 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4685; // @[lut_35.scala 1323:74 lut_35.scala 1347:39]
  wire  _GEN_4866 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4686; // @[lut_35.scala 1323:74 lut_35.scala 1348:39]
  wire  _GEN_4867 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4687; // @[lut_35.scala 1323:74 lut_35.scala 1349:39]
  wire  _GEN_4868 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4688; // @[lut_35.scala 1323:74 lut_35.scala 1350:39]
  wire  _GEN_4869 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4689; // @[lut_35.scala 1323:74 lut_35.scala 1351:39]
  wire  _GEN_4870 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4690; // @[lut_35.scala 1323:74 lut_35.scala 1352:39]
  wire  _GEN_4871 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4691; // @[lut_35.scala 1323:74 lut_35.scala 1353:39]
  wire  _GEN_4872 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4692; // @[lut_35.scala 1323:74 lut_35.scala 1354:39]
  wire  _GEN_4873 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4693; // @[lut_35.scala 1323:74 lut_35.scala 1355:39]
  wire  _GEN_4874 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4694; // @[lut_35.scala 1323:74 lut_35.scala 1356:39]
  wire  _GEN_4875 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4695; // @[lut_35.scala 1323:74 lut_35.scala 1357:39]
  wire  _GEN_4876 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4696; // @[lut_35.scala 1323:74 lut_35.scala 1358:39]
  wire  _GEN_4877 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid | _GEN_4697; // @[lut_35.scala 1323:74 lut_35.scala 1359:34]
  wire  _GEN_4881 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1323:74 lut_35.scala 216:26 lut_35.scala 1361:28]
  wire  _GEN_4884 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4701; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_4887 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4704; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_4890 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4707; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_4893 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4710; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_4896 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4713; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_4899 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4716; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_4902 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4719; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_4905 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4722; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_4908 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4725; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_4911 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4728; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_4914 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4731; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_4917 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4734; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_4920 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4737; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire [5:0] _GEN_4921 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? push_mem_temp : _GEN_4738; // @[lut_35.scala 1323:74 lut_35.scala 521:39]
  wire [31:0] _GEN_4922 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? push_id_temp : _GEN_4739; // @[lut_35.scala 1323:74 lut_35.scala 522:39]
  wire  _GEN_4925 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4742; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_4928 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4745; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_4931 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4748; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_4934 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4751; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_4937 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4754; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_4940 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4757; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_4943 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4760; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_4946 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4763; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_4949 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4766; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_4952 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4769; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_4955 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4772; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_4958 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4775; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_4961 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4778; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_4964 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4781; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_4967 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4784; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_4970 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4787; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_4973 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4790; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_4976 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4793; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_4979 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4796; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_4982 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4799; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_4985 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4802; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_4988 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4805; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_4991 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4808; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_4994 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4811; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_4997 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4814; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_5000 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4817; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_5003 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4820; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_5006 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4823; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_5009 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4826; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_5012 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4829; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_5015 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4832; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_5018 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4835; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_5021 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4838; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_5024 = LUT_mem_MPORT_56_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4841; // @[lut_35.scala 1323:74 lut_35.scala 216:26]
  wire  _GEN_5025 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4842; // @[lut_35.scala 1285:74 lut_35.scala 1286:38]
  wire  _GEN_5026 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4843; // @[lut_35.scala 1285:74 lut_35.scala 1287:38]
  wire  _GEN_5027 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4844; // @[lut_35.scala 1285:74 lut_35.scala 1288:38]
  wire  _GEN_5028 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4845; // @[lut_35.scala 1285:74 lut_35.scala 1289:38]
  wire  _GEN_5029 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4846; // @[lut_35.scala 1285:74 lut_35.scala 1290:38]
  wire  _GEN_5030 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4847; // @[lut_35.scala 1285:74 lut_35.scala 1291:38]
  wire  _GEN_5031 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4848; // @[lut_35.scala 1285:74 lut_35.scala 1292:38]
  wire  _GEN_5032 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4849; // @[lut_35.scala 1285:74 lut_35.scala 1293:38]
  wire  _GEN_5033 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4850; // @[lut_35.scala 1285:74 lut_35.scala 1294:38]
  wire  _GEN_5034 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4851; // @[lut_35.scala 1285:74 lut_35.scala 1295:38]
  wire  _GEN_5035 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4852; // @[lut_35.scala 1285:74 lut_35.scala 1296:39]
  wire  _GEN_5036 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4853; // @[lut_35.scala 1285:74 lut_35.scala 1297:39]
  wire  _GEN_5037 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4854; // @[lut_35.scala 1285:74 lut_35.scala 1298:39]
  wire  _GEN_5038 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4855; // @[lut_35.scala 1285:74 lut_35.scala 1299:39]
  wire  _GEN_5039 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4856; // @[lut_35.scala 1285:74 lut_35.scala 1300:39]
  wire  _GEN_5040 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4857; // @[lut_35.scala 1285:74 lut_35.scala 1301:39]
  wire  _GEN_5041 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4858; // @[lut_35.scala 1285:74 lut_35.scala 1302:39]
  wire  _GEN_5042 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4859; // @[lut_35.scala 1285:74 lut_35.scala 1303:39]
  wire  _GEN_5043 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4860; // @[lut_35.scala 1285:74 lut_35.scala 1304:39]
  wire  _GEN_5044 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4861; // @[lut_35.scala 1285:74 lut_35.scala 1305:39]
  wire  _GEN_5045 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid | _GEN_4862; // @[lut_35.scala 1285:74 lut_35.scala 1306:39]
  wire  _GEN_5046 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4863; // @[lut_35.scala 1285:74 lut_35.scala 1307:39]
  wire  _GEN_5047 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4864; // @[lut_35.scala 1285:74 lut_35.scala 1308:39]
  wire  _GEN_5048 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4865; // @[lut_35.scala 1285:74 lut_35.scala 1309:39]
  wire  _GEN_5049 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4866; // @[lut_35.scala 1285:74 lut_35.scala 1310:39]
  wire  _GEN_5050 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4867; // @[lut_35.scala 1285:74 lut_35.scala 1311:39]
  wire  _GEN_5051 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4868; // @[lut_35.scala 1285:74 lut_35.scala 1312:39]
  wire  _GEN_5052 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4869; // @[lut_35.scala 1285:74 lut_35.scala 1313:39]
  wire  _GEN_5053 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4870; // @[lut_35.scala 1285:74 lut_35.scala 1314:39]
  wire  _GEN_5054 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4871; // @[lut_35.scala 1285:74 lut_35.scala 1315:39]
  wire  _GEN_5055 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4872; // @[lut_35.scala 1285:74 lut_35.scala 1316:39]
  wire  _GEN_5056 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4873; // @[lut_35.scala 1285:74 lut_35.scala 1317:39]
  wire  _GEN_5057 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4874; // @[lut_35.scala 1285:74 lut_35.scala 1318:39]
  wire  _GEN_5058 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4875; // @[lut_35.scala 1285:74 lut_35.scala 1319:39]
  wire  _GEN_5059 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4876; // @[lut_35.scala 1285:74 lut_35.scala 1320:39]
  wire  _GEN_5060 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid | _GEN_4877; // @[lut_35.scala 1285:74 lut_35.scala 1321:34]
  wire  _GEN_5064 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1285:74 lut_35.scala 216:26 lut_35.scala 1323:27]
  wire  _GEN_5067 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4881; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5070 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4884; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5073 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4887; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5076 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4890; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5079 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4893; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5082 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4896; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5085 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4899; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5088 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4902; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5091 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4905; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5094 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4908; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5097 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4911; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5100 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4914; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5103 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4917; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5106 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4920; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire [5:0] _GEN_5107 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? push_mem_temp : _GEN_4921; // @[lut_35.scala 1285:74 lut_35.scala 521:39]
  wire [31:0] _GEN_5108 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? push_id_temp : _GEN_4922; // @[lut_35.scala 1285:74 lut_35.scala 522:39]
  wire  _GEN_5111 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4925; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5114 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4928; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5117 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4931; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5120 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4934; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5123 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4937; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5126 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4940; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5129 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4943; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5132 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4946; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5135 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4949; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5138 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4952; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5141 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4955; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5144 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4958; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5147 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4961; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5150 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4964; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5153 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4967; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5156 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4970; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5159 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4973; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5162 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4976; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5165 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4979; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5168 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4982; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5171 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4985; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5174 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4988; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5177 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4991; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5180 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4994; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5183 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_4997; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5186 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5000; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5189 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5003; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5192 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5006; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5195 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5009; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5198 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5012; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5201 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5015; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5204 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5018; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5207 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5021; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5210 = LUT_mem_MPORT_55_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5024; // @[lut_35.scala 1285:74 lut_35.scala 216:26]
  wire  _GEN_5211 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5025; // @[lut_35.scala 1247:74 lut_35.scala 1248:38]
  wire  _GEN_5212 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5026; // @[lut_35.scala 1247:74 lut_35.scala 1249:38]
  wire  _GEN_5213 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5027; // @[lut_35.scala 1247:74 lut_35.scala 1250:38]
  wire  _GEN_5214 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5028; // @[lut_35.scala 1247:74 lut_35.scala 1251:38]
  wire  _GEN_5215 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5029; // @[lut_35.scala 1247:74 lut_35.scala 1252:38]
  wire  _GEN_5216 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5030; // @[lut_35.scala 1247:74 lut_35.scala 1253:38]
  wire  _GEN_5217 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5031; // @[lut_35.scala 1247:74 lut_35.scala 1254:38]
  wire  _GEN_5218 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5032; // @[lut_35.scala 1247:74 lut_35.scala 1255:38]
  wire  _GEN_5219 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5033; // @[lut_35.scala 1247:74 lut_35.scala 1256:38]
  wire  _GEN_5220 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5034; // @[lut_35.scala 1247:74 lut_35.scala 1257:38]
  wire  _GEN_5221 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5035; // @[lut_35.scala 1247:74 lut_35.scala 1258:39]
  wire  _GEN_5222 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5036; // @[lut_35.scala 1247:74 lut_35.scala 1259:39]
  wire  _GEN_5223 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5037; // @[lut_35.scala 1247:74 lut_35.scala 1260:39]
  wire  _GEN_5224 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5038; // @[lut_35.scala 1247:74 lut_35.scala 1261:39]
  wire  _GEN_5225 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5039; // @[lut_35.scala 1247:74 lut_35.scala 1262:39]
  wire  _GEN_5226 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5040; // @[lut_35.scala 1247:74 lut_35.scala 1263:39]
  wire  _GEN_5227 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5041; // @[lut_35.scala 1247:74 lut_35.scala 1264:39]
  wire  _GEN_5228 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5042; // @[lut_35.scala 1247:74 lut_35.scala 1265:39]
  wire  _GEN_5229 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5043; // @[lut_35.scala 1247:74 lut_35.scala 1266:39]
  wire  _GEN_5230 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid | _GEN_5044; // @[lut_35.scala 1247:74 lut_35.scala 1267:39]
  wire  _GEN_5231 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5045; // @[lut_35.scala 1247:74 lut_35.scala 1268:39]
  wire  _GEN_5232 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5046; // @[lut_35.scala 1247:74 lut_35.scala 1269:39]
  wire  _GEN_5233 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5047; // @[lut_35.scala 1247:74 lut_35.scala 1270:39]
  wire  _GEN_5234 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5048; // @[lut_35.scala 1247:74 lut_35.scala 1271:39]
  wire  _GEN_5235 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5049; // @[lut_35.scala 1247:74 lut_35.scala 1272:39]
  wire  _GEN_5236 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5050; // @[lut_35.scala 1247:74 lut_35.scala 1273:39]
  wire  _GEN_5237 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5051; // @[lut_35.scala 1247:74 lut_35.scala 1274:39]
  wire  _GEN_5238 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5052; // @[lut_35.scala 1247:74 lut_35.scala 1275:39]
  wire  _GEN_5239 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5053; // @[lut_35.scala 1247:74 lut_35.scala 1276:39]
  wire  _GEN_5240 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5054; // @[lut_35.scala 1247:74 lut_35.scala 1277:39]
  wire  _GEN_5241 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5055; // @[lut_35.scala 1247:74 lut_35.scala 1278:39]
  wire  _GEN_5242 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5056; // @[lut_35.scala 1247:74 lut_35.scala 1279:39]
  wire  _GEN_5243 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5057; // @[lut_35.scala 1247:74 lut_35.scala 1280:39]
  wire  _GEN_5244 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5058; // @[lut_35.scala 1247:74 lut_35.scala 1281:39]
  wire  _GEN_5245 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5059; // @[lut_35.scala 1247:74 lut_35.scala 1282:39]
  wire  _GEN_5246 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid | _GEN_5060; // @[lut_35.scala 1247:74 lut_35.scala 1283:34]
  wire  _GEN_5250 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1247:74 lut_35.scala 216:26 lut_35.scala 1285:27]
  wire  _GEN_5253 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5064; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5256 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5067; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5259 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5070; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5262 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5073; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5265 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5076; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5268 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5079; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5271 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5082; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5274 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5085; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5277 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5088; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5280 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5091; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5283 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5094; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5286 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5097; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5289 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5100; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5292 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5103; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5295 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5106; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire [5:0] _GEN_5296 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? push_mem_temp : _GEN_5107; // @[lut_35.scala 1247:74 lut_35.scala 521:39]
  wire [31:0] _GEN_5297 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? push_id_temp : _GEN_5108; // @[lut_35.scala 1247:74 lut_35.scala 522:39]
  wire  _GEN_5300 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5111; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5303 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5114; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5306 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5117; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5309 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5120; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5312 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5123; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5315 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5126; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5318 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5129; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5321 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5132; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5324 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5135; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5327 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5138; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5330 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5141; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5333 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5144; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5336 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5147; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5339 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5150; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5342 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5153; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5345 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5156; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5348 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5159; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5351 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5162; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5354 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5165; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5357 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5168; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5360 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5171; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5363 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5174; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5366 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5177; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5369 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5180; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5372 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5183; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5375 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5186; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5378 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5189; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5381 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5192; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5384 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5195; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5387 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5198; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5390 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5201; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5393 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5204; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5396 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5207; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5399 = LUT_mem_MPORT_54_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5210; // @[lut_35.scala 1247:74 lut_35.scala 216:26]
  wire  _GEN_5400 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5211; // @[lut_35.scala 1209:74 lut_35.scala 1210:38]
  wire  _GEN_5401 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5212; // @[lut_35.scala 1209:74 lut_35.scala 1211:38]
  wire  _GEN_5402 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5213; // @[lut_35.scala 1209:74 lut_35.scala 1212:38]
  wire  _GEN_5403 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5214; // @[lut_35.scala 1209:74 lut_35.scala 1213:38]
  wire  _GEN_5404 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5215; // @[lut_35.scala 1209:74 lut_35.scala 1214:38]
  wire  _GEN_5405 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5216; // @[lut_35.scala 1209:74 lut_35.scala 1215:38]
  wire  _GEN_5406 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5217; // @[lut_35.scala 1209:74 lut_35.scala 1216:38]
  wire  _GEN_5407 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5218; // @[lut_35.scala 1209:74 lut_35.scala 1217:38]
  wire  _GEN_5408 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5219; // @[lut_35.scala 1209:74 lut_35.scala 1218:38]
  wire  _GEN_5409 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5220; // @[lut_35.scala 1209:74 lut_35.scala 1219:38]
  wire  _GEN_5410 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5221; // @[lut_35.scala 1209:74 lut_35.scala 1220:39]
  wire  _GEN_5411 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5222; // @[lut_35.scala 1209:74 lut_35.scala 1221:39]
  wire  _GEN_5412 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5223; // @[lut_35.scala 1209:74 lut_35.scala 1222:39]
  wire  _GEN_5413 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5224; // @[lut_35.scala 1209:74 lut_35.scala 1223:39]
  wire  _GEN_5414 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5225; // @[lut_35.scala 1209:74 lut_35.scala 1224:39]
  wire  _GEN_5415 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5226; // @[lut_35.scala 1209:74 lut_35.scala 1225:39]
  wire  _GEN_5416 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5227; // @[lut_35.scala 1209:74 lut_35.scala 1226:39]
  wire  _GEN_5417 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5228; // @[lut_35.scala 1209:74 lut_35.scala 1227:39]
  wire  _GEN_5418 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid | _GEN_5229; // @[lut_35.scala 1209:74 lut_35.scala 1228:39]
  wire  _GEN_5419 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5230; // @[lut_35.scala 1209:74 lut_35.scala 1229:39]
  wire  _GEN_5420 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5231; // @[lut_35.scala 1209:74 lut_35.scala 1230:39]
  wire  _GEN_5421 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5232; // @[lut_35.scala 1209:74 lut_35.scala 1231:39]
  wire  _GEN_5422 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5233; // @[lut_35.scala 1209:74 lut_35.scala 1232:39]
  wire  _GEN_5423 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5234; // @[lut_35.scala 1209:74 lut_35.scala 1233:39]
  wire  _GEN_5424 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5235; // @[lut_35.scala 1209:74 lut_35.scala 1234:39]
  wire  _GEN_5425 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5236; // @[lut_35.scala 1209:74 lut_35.scala 1235:39]
  wire  _GEN_5426 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5237; // @[lut_35.scala 1209:74 lut_35.scala 1236:39]
  wire  _GEN_5427 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5238; // @[lut_35.scala 1209:74 lut_35.scala 1237:39]
  wire  _GEN_5428 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5239; // @[lut_35.scala 1209:74 lut_35.scala 1238:39]
  wire  _GEN_5429 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5240; // @[lut_35.scala 1209:74 lut_35.scala 1239:39]
  wire  _GEN_5430 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5241; // @[lut_35.scala 1209:74 lut_35.scala 1240:39]
  wire  _GEN_5431 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5242; // @[lut_35.scala 1209:74 lut_35.scala 1241:39]
  wire  _GEN_5432 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5243; // @[lut_35.scala 1209:74 lut_35.scala 1242:39]
  wire  _GEN_5433 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5244; // @[lut_35.scala 1209:74 lut_35.scala 1243:39]
  wire  _GEN_5434 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5245; // @[lut_35.scala 1209:74 lut_35.scala 1244:39]
  wire  _GEN_5435 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid | _GEN_5246; // @[lut_35.scala 1209:74 lut_35.scala 1245:34]
  wire  _GEN_5439 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1209:74 lut_35.scala 216:26 lut_35.scala 1247:27]
  wire  _GEN_5442 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5250; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5445 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5253; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5448 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5256; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5451 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5259; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5454 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5262; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5457 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5265; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5460 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5268; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5463 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5271; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5466 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5274; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5469 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5277; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5472 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5280; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5475 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5283; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5478 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5286; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5481 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5289; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5484 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5292; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5487 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5295; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire [5:0] _GEN_5488 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? push_mem_temp : _GEN_5296; // @[lut_35.scala 1209:74 lut_35.scala 521:39]
  wire [31:0] _GEN_5489 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? push_id_temp : _GEN_5297; // @[lut_35.scala 1209:74 lut_35.scala 522:39]
  wire  _GEN_5492 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5300; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5495 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5303; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5498 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5306; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5501 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5309; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5504 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5312; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5507 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5315; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5510 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5318; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5513 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5321; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5516 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5324; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5519 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5327; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5522 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5330; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5525 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5333; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5528 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5336; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5531 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5339; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5534 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5342; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5537 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5345; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5540 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5348; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5543 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5351; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5546 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5354; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5549 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5357; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5552 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5360; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5555 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5363; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5558 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5366; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5561 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5369; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5564 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5372; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5567 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5375; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5570 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5378; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5573 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5381; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5576 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5384; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5579 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5387; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5582 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5390; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5585 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5393; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5588 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5396; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5591 = LUT_mem_MPORT_53_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5399; // @[lut_35.scala 1209:74 lut_35.scala 216:26]
  wire  _GEN_5592 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5400; // @[lut_35.scala 1171:74 lut_35.scala 1172:38]
  wire  _GEN_5593 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5401; // @[lut_35.scala 1171:74 lut_35.scala 1173:38]
  wire  _GEN_5594 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5402; // @[lut_35.scala 1171:74 lut_35.scala 1174:38]
  wire  _GEN_5595 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5403; // @[lut_35.scala 1171:74 lut_35.scala 1175:38]
  wire  _GEN_5596 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5404; // @[lut_35.scala 1171:74 lut_35.scala 1176:38]
  wire  _GEN_5597 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5405; // @[lut_35.scala 1171:74 lut_35.scala 1177:38]
  wire  _GEN_5598 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5406; // @[lut_35.scala 1171:74 lut_35.scala 1178:38]
  wire  _GEN_5599 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5407; // @[lut_35.scala 1171:74 lut_35.scala 1179:38]
  wire  _GEN_5600 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5408; // @[lut_35.scala 1171:74 lut_35.scala 1180:38]
  wire  _GEN_5601 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5409; // @[lut_35.scala 1171:74 lut_35.scala 1181:38]
  wire  _GEN_5602 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5410; // @[lut_35.scala 1171:74 lut_35.scala 1182:39]
  wire  _GEN_5603 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5411; // @[lut_35.scala 1171:74 lut_35.scala 1183:39]
  wire  _GEN_5604 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5412; // @[lut_35.scala 1171:74 lut_35.scala 1184:39]
  wire  _GEN_5605 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5413; // @[lut_35.scala 1171:74 lut_35.scala 1185:39]
  wire  _GEN_5606 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5414; // @[lut_35.scala 1171:74 lut_35.scala 1186:39]
  wire  _GEN_5607 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5415; // @[lut_35.scala 1171:74 lut_35.scala 1187:39]
  wire  _GEN_5608 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5416; // @[lut_35.scala 1171:74 lut_35.scala 1188:39]
  wire  _GEN_5609 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid | _GEN_5417; // @[lut_35.scala 1171:74 lut_35.scala 1189:39]
  wire  _GEN_5610 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5418; // @[lut_35.scala 1171:74 lut_35.scala 1190:39]
  wire  _GEN_5611 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5419; // @[lut_35.scala 1171:74 lut_35.scala 1191:39]
  wire  _GEN_5612 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5420; // @[lut_35.scala 1171:74 lut_35.scala 1192:39]
  wire  _GEN_5613 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5421; // @[lut_35.scala 1171:74 lut_35.scala 1193:39]
  wire  _GEN_5614 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5422; // @[lut_35.scala 1171:74 lut_35.scala 1194:39]
  wire  _GEN_5615 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5423; // @[lut_35.scala 1171:74 lut_35.scala 1195:39]
  wire  _GEN_5616 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5424; // @[lut_35.scala 1171:74 lut_35.scala 1196:39]
  wire  _GEN_5617 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5425; // @[lut_35.scala 1171:74 lut_35.scala 1197:39]
  wire  _GEN_5618 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5426; // @[lut_35.scala 1171:74 lut_35.scala 1198:39]
  wire  _GEN_5619 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5427; // @[lut_35.scala 1171:74 lut_35.scala 1199:39]
  wire  _GEN_5620 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5428; // @[lut_35.scala 1171:74 lut_35.scala 1200:39]
  wire  _GEN_5621 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5429; // @[lut_35.scala 1171:74 lut_35.scala 1201:39]
  wire  _GEN_5622 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5430; // @[lut_35.scala 1171:74 lut_35.scala 1202:39]
  wire  _GEN_5623 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5431; // @[lut_35.scala 1171:74 lut_35.scala 1203:39]
  wire  _GEN_5624 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5432; // @[lut_35.scala 1171:74 lut_35.scala 1204:39]
  wire  _GEN_5625 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5433; // @[lut_35.scala 1171:74 lut_35.scala 1205:39]
  wire  _GEN_5626 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5434; // @[lut_35.scala 1171:74 lut_35.scala 1206:39]
  wire  _GEN_5627 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid | _GEN_5435; // @[lut_35.scala 1171:74 lut_35.scala 1207:34]
  wire  _GEN_5631 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1171:74 lut_35.scala 216:26 lut_35.scala 1209:27]
  wire  _GEN_5634 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5439; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5637 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5442; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5640 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5445; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5643 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5448; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5646 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5451; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5649 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5454; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5652 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5457; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5655 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5460; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5658 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5463; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5661 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5466; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5664 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5469; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5667 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5472; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5670 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5475; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5673 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5478; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5676 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5481; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5679 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5484; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5682 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5487; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire [5:0] _GEN_5683 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? push_mem_temp : _GEN_5488; // @[lut_35.scala 1171:74 lut_35.scala 521:39]
  wire [31:0] _GEN_5684 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? push_id_temp : _GEN_5489; // @[lut_35.scala 1171:74 lut_35.scala 522:39]
  wire  _GEN_5687 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5492; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5690 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5495; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5693 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5498; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5696 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5501; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5699 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5504; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5702 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5507; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5705 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5510; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5708 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5513; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5711 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5516; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5714 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5519; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5717 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5522; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5720 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5525; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5723 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5528; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5726 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5531; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5729 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5534; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5732 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5537; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5735 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5540; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5738 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5543; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5741 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5546; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5744 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5549; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5747 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5552; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5750 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5555; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5753 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5558; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5756 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5561; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5759 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5564; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5762 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5567; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5765 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5570; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5768 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5573; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5771 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5576; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5774 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5579; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5777 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5582; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5780 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5585; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5783 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5588; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5786 = LUT_mem_MPORT_52_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5591; // @[lut_35.scala 1171:74 lut_35.scala 216:26]
  wire  _GEN_5787 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5592; // @[lut_35.scala 1133:74 lut_35.scala 1134:38]
  wire  _GEN_5788 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5593; // @[lut_35.scala 1133:74 lut_35.scala 1135:38]
  wire  _GEN_5789 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5594; // @[lut_35.scala 1133:74 lut_35.scala 1136:38]
  wire  _GEN_5790 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5595; // @[lut_35.scala 1133:74 lut_35.scala 1137:38]
  wire  _GEN_5791 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5596; // @[lut_35.scala 1133:74 lut_35.scala 1138:38]
  wire  _GEN_5792 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5597; // @[lut_35.scala 1133:74 lut_35.scala 1139:38]
  wire  _GEN_5793 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5598; // @[lut_35.scala 1133:74 lut_35.scala 1140:38]
  wire  _GEN_5794 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5599; // @[lut_35.scala 1133:74 lut_35.scala 1141:38]
  wire  _GEN_5795 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5600; // @[lut_35.scala 1133:74 lut_35.scala 1142:38]
  wire  _GEN_5796 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5601; // @[lut_35.scala 1133:74 lut_35.scala 1143:38]
  wire  _GEN_5797 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5602; // @[lut_35.scala 1133:74 lut_35.scala 1144:39]
  wire  _GEN_5798 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5603; // @[lut_35.scala 1133:74 lut_35.scala 1145:39]
  wire  _GEN_5799 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5604; // @[lut_35.scala 1133:74 lut_35.scala 1146:39]
  wire  _GEN_5800 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5605; // @[lut_35.scala 1133:74 lut_35.scala 1147:39]
  wire  _GEN_5801 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5606; // @[lut_35.scala 1133:74 lut_35.scala 1148:39]
  wire  _GEN_5802 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5607; // @[lut_35.scala 1133:74 lut_35.scala 1149:39]
  wire  _GEN_5803 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid | _GEN_5608; // @[lut_35.scala 1133:74 lut_35.scala 1150:39]
  wire  _GEN_5804 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5609; // @[lut_35.scala 1133:74 lut_35.scala 1151:39]
  wire  _GEN_5805 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5610; // @[lut_35.scala 1133:74 lut_35.scala 1152:39]
  wire  _GEN_5806 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5611; // @[lut_35.scala 1133:74 lut_35.scala 1153:39]
  wire  _GEN_5807 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5612; // @[lut_35.scala 1133:74 lut_35.scala 1154:39]
  wire  _GEN_5808 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5613; // @[lut_35.scala 1133:74 lut_35.scala 1155:39]
  wire  _GEN_5809 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5614; // @[lut_35.scala 1133:74 lut_35.scala 1156:39]
  wire  _GEN_5810 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5615; // @[lut_35.scala 1133:74 lut_35.scala 1157:39]
  wire  _GEN_5811 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5616; // @[lut_35.scala 1133:74 lut_35.scala 1158:39]
  wire  _GEN_5812 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5617; // @[lut_35.scala 1133:74 lut_35.scala 1159:39]
  wire  _GEN_5813 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5618; // @[lut_35.scala 1133:74 lut_35.scala 1160:39]
  wire  _GEN_5814 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5619; // @[lut_35.scala 1133:74 lut_35.scala 1161:39]
  wire  _GEN_5815 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5620; // @[lut_35.scala 1133:74 lut_35.scala 1162:39]
  wire  _GEN_5816 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5621; // @[lut_35.scala 1133:74 lut_35.scala 1163:39]
  wire  _GEN_5817 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5622; // @[lut_35.scala 1133:74 lut_35.scala 1164:39]
  wire  _GEN_5818 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5623; // @[lut_35.scala 1133:74 lut_35.scala 1165:39]
  wire  _GEN_5819 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5624; // @[lut_35.scala 1133:74 lut_35.scala 1166:39]
  wire  _GEN_5820 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5625; // @[lut_35.scala 1133:74 lut_35.scala 1167:39]
  wire  _GEN_5821 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5626; // @[lut_35.scala 1133:74 lut_35.scala 1168:39]
  wire  _GEN_5822 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid | _GEN_5627; // @[lut_35.scala 1133:74 lut_35.scala 1169:34]
  wire  _GEN_5826 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1133:74 lut_35.scala 216:26 lut_35.scala 1171:27]
  wire  _GEN_5829 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5631; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5832 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5634; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5835 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5637; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5838 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5640; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5841 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5643; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5844 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5646; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5847 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5649; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5850 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5652; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5853 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5655; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5856 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5658; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5859 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5661; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5862 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5664; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5865 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5667; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5868 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5670; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5871 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5673; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5874 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5676; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5877 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5679; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5880 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5682; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire [5:0] _GEN_5881 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? push_mem_temp : _GEN_5683; // @[lut_35.scala 1133:74 lut_35.scala 521:39]
  wire [31:0] _GEN_5882 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? push_id_temp : _GEN_5684; // @[lut_35.scala 1133:74 lut_35.scala 522:39]
  wire  _GEN_5885 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5687; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5888 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5690; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5891 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5693; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5894 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5696; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5897 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5699; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5900 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5702; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5903 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5705; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5906 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5708; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5909 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5711; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5912 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5714; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5915 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5717; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5918 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5720; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5921 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5723; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5924 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5726; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5927 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5729; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5930 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5732; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5933 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5735; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5936 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5738; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5939 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5741; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5942 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5744; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5945 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5747; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5948 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5750; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5951 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5753; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5954 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5756; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5957 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5759; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5960 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5762; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5963 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5765; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5966 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5768; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5969 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5771; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5972 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5774; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5975 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5777; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5978 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5780; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5981 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5783; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5984 = LUT_mem_MPORT_51_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5786; // @[lut_35.scala 1133:74 lut_35.scala 216:26]
  wire  _GEN_5985 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5787; // @[lut_35.scala 1095:74 lut_35.scala 1096:38]
  wire  _GEN_5986 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5788; // @[lut_35.scala 1095:74 lut_35.scala 1097:38]
  wire  _GEN_5987 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5789; // @[lut_35.scala 1095:74 lut_35.scala 1098:38]
  wire  _GEN_5988 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5790; // @[lut_35.scala 1095:74 lut_35.scala 1099:38]
  wire  _GEN_5989 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5791; // @[lut_35.scala 1095:74 lut_35.scala 1100:38]
  wire  _GEN_5990 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5792; // @[lut_35.scala 1095:74 lut_35.scala 1101:38]
  wire  _GEN_5991 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5793; // @[lut_35.scala 1095:74 lut_35.scala 1102:38]
  wire  _GEN_5992 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5794; // @[lut_35.scala 1095:74 lut_35.scala 1103:38]
  wire  _GEN_5993 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5795; // @[lut_35.scala 1095:74 lut_35.scala 1104:38]
  wire  _GEN_5994 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5796; // @[lut_35.scala 1095:74 lut_35.scala 1105:38]
  wire  _GEN_5995 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5797; // @[lut_35.scala 1095:74 lut_35.scala 1106:39]
  wire  _GEN_5996 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5798; // @[lut_35.scala 1095:74 lut_35.scala 1107:39]
  wire  _GEN_5997 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5799; // @[lut_35.scala 1095:74 lut_35.scala 1108:39]
  wire  _GEN_5998 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5800; // @[lut_35.scala 1095:74 lut_35.scala 1109:39]
  wire  _GEN_5999 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5801; // @[lut_35.scala 1095:74 lut_35.scala 1110:39]
  wire  _GEN_6000 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid | _GEN_5802; // @[lut_35.scala 1095:74 lut_35.scala 1111:39]
  wire  _GEN_6001 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5803; // @[lut_35.scala 1095:74 lut_35.scala 1112:39]
  wire  _GEN_6002 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5804; // @[lut_35.scala 1095:74 lut_35.scala 1113:39]
  wire  _GEN_6003 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5805; // @[lut_35.scala 1095:74 lut_35.scala 1114:39]
  wire  _GEN_6004 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5806; // @[lut_35.scala 1095:74 lut_35.scala 1115:39]
  wire  _GEN_6005 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5807; // @[lut_35.scala 1095:74 lut_35.scala 1116:39]
  wire  _GEN_6006 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5808; // @[lut_35.scala 1095:74 lut_35.scala 1117:39]
  wire  _GEN_6007 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5809; // @[lut_35.scala 1095:74 lut_35.scala 1118:39]
  wire  _GEN_6008 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5810; // @[lut_35.scala 1095:74 lut_35.scala 1119:39]
  wire  _GEN_6009 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5811; // @[lut_35.scala 1095:74 lut_35.scala 1120:39]
  wire  _GEN_6010 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5812; // @[lut_35.scala 1095:74 lut_35.scala 1121:39]
  wire  _GEN_6011 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5813; // @[lut_35.scala 1095:74 lut_35.scala 1122:39]
  wire  _GEN_6012 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5814; // @[lut_35.scala 1095:74 lut_35.scala 1123:39]
  wire  _GEN_6013 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5815; // @[lut_35.scala 1095:74 lut_35.scala 1124:39]
  wire  _GEN_6014 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5816; // @[lut_35.scala 1095:74 lut_35.scala 1125:39]
  wire  _GEN_6015 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5817; // @[lut_35.scala 1095:74 lut_35.scala 1126:39]
  wire  _GEN_6016 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5818; // @[lut_35.scala 1095:74 lut_35.scala 1127:39]
  wire  _GEN_6017 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5819; // @[lut_35.scala 1095:74 lut_35.scala 1128:39]
  wire  _GEN_6018 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5820; // @[lut_35.scala 1095:74 lut_35.scala 1129:39]
  wire  _GEN_6019 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5821; // @[lut_35.scala 1095:74 lut_35.scala 1130:39]
  wire  _GEN_6020 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid | _GEN_5822; // @[lut_35.scala 1095:74 lut_35.scala 1131:34]
  wire  _GEN_6024 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1095:74 lut_35.scala 216:26 lut_35.scala 1133:27]
  wire  _GEN_6027 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5826; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6030 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5829; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6033 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5832; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6036 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5835; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6039 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5838; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6042 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5841; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6045 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5844; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6048 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5847; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6051 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5850; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6054 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5853; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6057 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5856; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6060 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5859; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6063 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5862; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6066 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5865; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6069 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5868; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6072 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5871; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6075 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5874; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6078 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5877; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6081 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5880; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire [5:0] _GEN_6082 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? push_mem_temp : _GEN_5881; // @[lut_35.scala 1095:74 lut_35.scala 521:39]
  wire [31:0] _GEN_6083 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? push_id_temp : _GEN_5882; // @[lut_35.scala 1095:74 lut_35.scala 522:39]
  wire  _GEN_6086 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5885; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6089 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5888; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6092 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5891; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6095 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5894; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6098 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5897; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6101 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5900; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6104 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5903; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6107 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5906; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6110 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5909; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6113 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5912; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6116 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5915; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6119 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5918; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6122 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5921; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6125 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5924; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6128 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5927; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6131 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5930; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6134 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5933; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6137 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5936; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6140 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5939; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6143 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5942; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6146 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5945; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6149 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5948; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6152 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5951; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6155 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5954; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6158 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5957; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6161 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5960; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6164 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5963; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6167 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5966; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6170 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5969; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6173 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5972; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6176 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5975; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6179 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5978; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6182 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5981; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6185 = LUT_mem_MPORT_50_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5984; // @[lut_35.scala 1095:74 lut_35.scala 216:26]
  wire  _GEN_6186 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5985; // @[lut_35.scala 1057:74 lut_35.scala 1058:38]
  wire  _GEN_6187 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5986; // @[lut_35.scala 1057:74 lut_35.scala 1059:38]
  wire  _GEN_6188 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5987; // @[lut_35.scala 1057:74 lut_35.scala 1060:38]
  wire  _GEN_6189 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5988; // @[lut_35.scala 1057:74 lut_35.scala 1061:38]
  wire  _GEN_6190 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5989; // @[lut_35.scala 1057:74 lut_35.scala 1062:38]
  wire  _GEN_6191 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5990; // @[lut_35.scala 1057:74 lut_35.scala 1063:38]
  wire  _GEN_6192 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5991; // @[lut_35.scala 1057:74 lut_35.scala 1064:38]
  wire  _GEN_6193 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5992; // @[lut_35.scala 1057:74 lut_35.scala 1065:38]
  wire  _GEN_6194 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5993; // @[lut_35.scala 1057:74 lut_35.scala 1066:38]
  wire  _GEN_6195 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5994; // @[lut_35.scala 1057:74 lut_35.scala 1067:38]
  wire  _GEN_6196 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5995; // @[lut_35.scala 1057:74 lut_35.scala 1068:39]
  wire  _GEN_6197 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5996; // @[lut_35.scala 1057:74 lut_35.scala 1069:39]
  wire  _GEN_6198 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5997; // @[lut_35.scala 1057:74 lut_35.scala 1070:39]
  wire  _GEN_6199 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5998; // @[lut_35.scala 1057:74 lut_35.scala 1071:39]
  wire  _GEN_6200 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid | _GEN_5999; // @[lut_35.scala 1057:74 lut_35.scala 1072:39]
  wire  _GEN_6201 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6000; // @[lut_35.scala 1057:74 lut_35.scala 1073:39]
  wire  _GEN_6202 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6001; // @[lut_35.scala 1057:74 lut_35.scala 1074:39]
  wire  _GEN_6203 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6002; // @[lut_35.scala 1057:74 lut_35.scala 1075:39]
  wire  _GEN_6204 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6003; // @[lut_35.scala 1057:74 lut_35.scala 1076:39]
  wire  _GEN_6205 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6004; // @[lut_35.scala 1057:74 lut_35.scala 1077:39]
  wire  _GEN_6206 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6005; // @[lut_35.scala 1057:74 lut_35.scala 1078:39]
  wire  _GEN_6207 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6006; // @[lut_35.scala 1057:74 lut_35.scala 1079:39]
  wire  _GEN_6208 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6007; // @[lut_35.scala 1057:74 lut_35.scala 1080:39]
  wire  _GEN_6209 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6008; // @[lut_35.scala 1057:74 lut_35.scala 1081:39]
  wire  _GEN_6210 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6009; // @[lut_35.scala 1057:74 lut_35.scala 1082:39]
  wire  _GEN_6211 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6010; // @[lut_35.scala 1057:74 lut_35.scala 1083:39]
  wire  _GEN_6212 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6011; // @[lut_35.scala 1057:74 lut_35.scala 1084:39]
  wire  _GEN_6213 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6012; // @[lut_35.scala 1057:74 lut_35.scala 1085:39]
  wire  _GEN_6214 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6013; // @[lut_35.scala 1057:74 lut_35.scala 1086:39]
  wire  _GEN_6215 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6014; // @[lut_35.scala 1057:74 lut_35.scala 1087:39]
  wire  _GEN_6216 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6015; // @[lut_35.scala 1057:74 lut_35.scala 1088:39]
  wire  _GEN_6217 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6016; // @[lut_35.scala 1057:74 lut_35.scala 1089:39]
  wire  _GEN_6218 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6017; // @[lut_35.scala 1057:74 lut_35.scala 1090:39]
  wire  _GEN_6219 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6018; // @[lut_35.scala 1057:74 lut_35.scala 1091:39]
  wire  _GEN_6220 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6019; // @[lut_35.scala 1057:74 lut_35.scala 1092:39]
  wire  _GEN_6221 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid | _GEN_6020; // @[lut_35.scala 1057:74 lut_35.scala 1093:34]
  wire  _GEN_6225 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1057:74 lut_35.scala 216:26 lut_35.scala 1095:27]
  wire  _GEN_6228 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6024; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6231 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6027; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6234 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6030; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6237 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6033; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6240 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6036; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6243 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6039; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6246 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6042; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6249 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6045; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6252 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6048; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6255 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6051; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6258 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6054; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6261 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6057; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6264 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6060; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6267 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6063; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6270 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6066; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6273 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6069; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6276 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6072; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6279 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6075; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6282 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6078; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6285 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6081; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire [5:0] _GEN_6286 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? push_mem_temp : _GEN_6082; // @[lut_35.scala 1057:74 lut_35.scala 521:39]
  wire [31:0] _GEN_6287 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? push_id_temp : _GEN_6083; // @[lut_35.scala 1057:74 lut_35.scala 522:39]
  wire  _GEN_6290 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6086; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6293 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6089; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6296 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6092; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6299 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6095; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6302 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6098; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6305 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6101; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6308 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6104; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6311 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6107; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6314 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6110; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6317 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6113; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6320 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6116; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6323 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6119; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6326 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6122; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6329 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6125; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6332 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6128; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6335 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6131; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6338 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6134; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6341 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6137; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6344 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6140; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6347 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6143; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6350 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6146; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6353 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6149; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6356 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6152; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6359 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6155; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6362 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6158; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6365 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6161; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6368 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6164; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6371 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6167; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6374 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6170; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6377 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6173; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6380 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6176; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6383 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6179; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6386 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6182; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6389 = LUT_mem_MPORT_49_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6185; // @[lut_35.scala 1057:74 lut_35.scala 216:26]
  wire  _GEN_6390 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6186; // @[lut_35.scala 1019:74 lut_35.scala 1020:38]
  wire  _GEN_6391 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6187; // @[lut_35.scala 1019:74 lut_35.scala 1021:38]
  wire  _GEN_6392 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6188; // @[lut_35.scala 1019:74 lut_35.scala 1022:38]
  wire  _GEN_6393 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6189; // @[lut_35.scala 1019:74 lut_35.scala 1023:38]
  wire  _GEN_6394 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6190; // @[lut_35.scala 1019:74 lut_35.scala 1024:38]
  wire  _GEN_6395 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6191; // @[lut_35.scala 1019:74 lut_35.scala 1025:38]
  wire  _GEN_6396 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6192; // @[lut_35.scala 1019:74 lut_35.scala 1026:38]
  wire  _GEN_6397 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6193; // @[lut_35.scala 1019:74 lut_35.scala 1027:38]
  wire  _GEN_6398 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6194; // @[lut_35.scala 1019:74 lut_35.scala 1028:38]
  wire  _GEN_6399 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6195; // @[lut_35.scala 1019:74 lut_35.scala 1029:38]
  wire  _GEN_6400 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6196; // @[lut_35.scala 1019:74 lut_35.scala 1030:39]
  wire  _GEN_6401 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6197; // @[lut_35.scala 1019:74 lut_35.scala 1031:39]
  wire  _GEN_6402 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6198; // @[lut_35.scala 1019:74 lut_35.scala 1032:39]
  wire  _GEN_6403 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid | _GEN_6199; // @[lut_35.scala 1019:74 lut_35.scala 1033:39]
  wire  _GEN_6404 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6200; // @[lut_35.scala 1019:74 lut_35.scala 1034:39]
  wire  _GEN_6405 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6201; // @[lut_35.scala 1019:74 lut_35.scala 1035:39]
  wire  _GEN_6406 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6202; // @[lut_35.scala 1019:74 lut_35.scala 1036:39]
  wire  _GEN_6407 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6203; // @[lut_35.scala 1019:74 lut_35.scala 1037:39]
  wire  _GEN_6408 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6204; // @[lut_35.scala 1019:74 lut_35.scala 1038:39]
  wire  _GEN_6409 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6205; // @[lut_35.scala 1019:74 lut_35.scala 1039:39]
  wire  _GEN_6410 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6206; // @[lut_35.scala 1019:74 lut_35.scala 1040:39]
  wire  _GEN_6411 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6207; // @[lut_35.scala 1019:74 lut_35.scala 1041:39]
  wire  _GEN_6412 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6208; // @[lut_35.scala 1019:74 lut_35.scala 1042:39]
  wire  _GEN_6413 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6209; // @[lut_35.scala 1019:74 lut_35.scala 1043:39]
  wire  _GEN_6414 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6210; // @[lut_35.scala 1019:74 lut_35.scala 1044:39]
  wire  _GEN_6415 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6211; // @[lut_35.scala 1019:74 lut_35.scala 1045:39]
  wire  _GEN_6416 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6212; // @[lut_35.scala 1019:74 lut_35.scala 1046:39]
  wire  _GEN_6417 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6213; // @[lut_35.scala 1019:74 lut_35.scala 1047:39]
  wire  _GEN_6418 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6214; // @[lut_35.scala 1019:74 lut_35.scala 1048:39]
  wire  _GEN_6419 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6215; // @[lut_35.scala 1019:74 lut_35.scala 1049:39]
  wire  _GEN_6420 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6216; // @[lut_35.scala 1019:74 lut_35.scala 1050:39]
  wire  _GEN_6421 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6217; // @[lut_35.scala 1019:74 lut_35.scala 1051:39]
  wire  _GEN_6422 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6218; // @[lut_35.scala 1019:74 lut_35.scala 1052:39]
  wire  _GEN_6423 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6219; // @[lut_35.scala 1019:74 lut_35.scala 1053:39]
  wire  _GEN_6424 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6220; // @[lut_35.scala 1019:74 lut_35.scala 1054:39]
  wire  _GEN_6425 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid | _GEN_6221; // @[lut_35.scala 1019:74 lut_35.scala 1055:34]
  wire  _GEN_6429 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1019:74 lut_35.scala 216:26 lut_35.scala 1057:27]
  wire  _GEN_6432 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6225; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6435 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6228; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6438 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6231; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6441 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6234; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6444 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6237; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6447 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6240; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6450 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6243; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6453 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6246; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6456 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6249; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6459 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6252; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6462 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6255; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6465 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6258; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6468 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6261; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6471 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6264; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6474 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6267; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6477 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6270; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6480 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6273; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6483 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6276; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6486 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6279; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6489 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6282; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6492 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6285; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire [5:0] _GEN_6493 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? push_mem_temp : _GEN_6286; // @[lut_35.scala 1019:74 lut_35.scala 521:39]
  wire [31:0] _GEN_6494 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? push_id_temp : _GEN_6287; // @[lut_35.scala 1019:74 lut_35.scala 522:39]
  wire  _GEN_6497 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6290; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6500 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6293; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6503 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6296; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6506 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6299; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6509 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6302; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6512 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6305; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6515 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6308; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6518 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6311; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6521 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6314; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6524 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6317; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6527 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6320; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6530 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6323; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6533 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6326; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6536 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6329; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6539 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6332; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6542 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6335; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6545 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6338; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6548 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6341; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6551 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6344; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6554 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6347; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6557 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6350; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6560 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6353; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6563 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6356; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6566 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6359; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6569 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6362; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6572 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6365; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6575 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6368; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6578 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6371; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6581 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6374; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6584 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6377; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6587 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6380; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6590 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6383; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6593 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6386; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6596 = LUT_mem_MPORT_48_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6389; // @[lut_35.scala 1019:74 lut_35.scala 216:26]
  wire  _GEN_6597 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6390; // @[lut_35.scala 981:74 lut_35.scala 982:38]
  wire  _GEN_6598 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6391; // @[lut_35.scala 981:74 lut_35.scala 983:38]
  wire  _GEN_6599 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6392; // @[lut_35.scala 981:74 lut_35.scala 984:38]
  wire  _GEN_6600 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6393; // @[lut_35.scala 981:74 lut_35.scala 985:38]
  wire  _GEN_6601 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6394; // @[lut_35.scala 981:74 lut_35.scala 986:38]
  wire  _GEN_6602 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6395; // @[lut_35.scala 981:74 lut_35.scala 987:38]
  wire  _GEN_6603 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6396; // @[lut_35.scala 981:74 lut_35.scala 988:38]
  wire  _GEN_6604 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6397; // @[lut_35.scala 981:74 lut_35.scala 989:38]
  wire  _GEN_6605 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6398; // @[lut_35.scala 981:74 lut_35.scala 990:38]
  wire  _GEN_6606 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6399; // @[lut_35.scala 981:74 lut_35.scala 991:38]
  wire  _GEN_6607 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6400; // @[lut_35.scala 981:74 lut_35.scala 992:39]
  wire  _GEN_6608 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6401; // @[lut_35.scala 981:74 lut_35.scala 993:39]
  wire  _GEN_6609 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid | _GEN_6402; // @[lut_35.scala 981:74 lut_35.scala 994:39]
  wire  _GEN_6610 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6403; // @[lut_35.scala 981:74 lut_35.scala 995:39]
  wire  _GEN_6611 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6404; // @[lut_35.scala 981:74 lut_35.scala 996:39]
  wire  _GEN_6612 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6405; // @[lut_35.scala 981:74 lut_35.scala 997:39]
  wire  _GEN_6613 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6406; // @[lut_35.scala 981:74 lut_35.scala 998:39]
  wire  _GEN_6614 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6407; // @[lut_35.scala 981:74 lut_35.scala 999:39]
  wire  _GEN_6615 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6408; // @[lut_35.scala 981:74 lut_35.scala 1000:39]
  wire  _GEN_6616 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6409; // @[lut_35.scala 981:74 lut_35.scala 1001:39]
  wire  _GEN_6617 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6410; // @[lut_35.scala 981:74 lut_35.scala 1002:39]
  wire  _GEN_6618 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6411; // @[lut_35.scala 981:74 lut_35.scala 1003:39]
  wire  _GEN_6619 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6412; // @[lut_35.scala 981:74 lut_35.scala 1004:39]
  wire  _GEN_6620 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6413; // @[lut_35.scala 981:74 lut_35.scala 1005:39]
  wire  _GEN_6621 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6414; // @[lut_35.scala 981:74 lut_35.scala 1006:39]
  wire  _GEN_6622 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6415; // @[lut_35.scala 981:74 lut_35.scala 1007:39]
  wire  _GEN_6623 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6416; // @[lut_35.scala 981:74 lut_35.scala 1008:39]
  wire  _GEN_6624 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6417; // @[lut_35.scala 981:74 lut_35.scala 1009:39]
  wire  _GEN_6625 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6418; // @[lut_35.scala 981:74 lut_35.scala 1010:39]
  wire  _GEN_6626 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6419; // @[lut_35.scala 981:74 lut_35.scala 1011:39]
  wire  _GEN_6627 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6420; // @[lut_35.scala 981:74 lut_35.scala 1012:39]
  wire  _GEN_6628 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6421; // @[lut_35.scala 981:74 lut_35.scala 1013:39]
  wire  _GEN_6629 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6422; // @[lut_35.scala 981:74 lut_35.scala 1014:39]
  wire  _GEN_6630 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6423; // @[lut_35.scala 981:74 lut_35.scala 1015:39]
  wire  _GEN_6631 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6424; // @[lut_35.scala 981:74 lut_35.scala 1016:39]
  wire  _GEN_6632 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid | _GEN_6425; // @[lut_35.scala 981:74 lut_35.scala 1017:34]
  wire  _GEN_6636 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 981:74 lut_35.scala 216:26 lut_35.scala 1019:27]
  wire  _GEN_6639 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6429; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6642 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6432; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6645 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6435; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6648 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6438; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6651 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6441; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6654 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6444; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6657 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6447; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6660 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6450; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6663 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6453; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6666 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6456; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6669 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6459; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6672 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6462; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6675 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6465; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6678 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6468; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6681 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6471; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6684 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6474; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6687 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6477; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6690 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6480; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6693 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6483; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6696 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6486; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6699 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6489; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6702 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6492; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire [5:0] _GEN_6703 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? push_mem_temp : _GEN_6493; // @[lut_35.scala 981:74 lut_35.scala 521:39]
  wire [31:0] _GEN_6704 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? push_id_temp : _GEN_6494; // @[lut_35.scala 981:74 lut_35.scala 522:39]
  wire  _GEN_6707 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6497; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6710 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6500; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6713 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6503; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6716 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6506; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6719 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6509; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6722 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6512; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6725 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6515; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6728 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6518; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6731 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6521; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6734 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6524; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6737 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6527; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6740 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6530; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6743 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6533; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6746 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6536; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6749 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6539; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6752 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6542; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6755 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6545; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6758 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6548; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6761 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6551; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6764 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6554; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6767 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6557; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6770 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6560; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6773 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6563; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6776 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6566; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6779 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6569; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6782 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6572; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6785 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6575; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6788 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6578; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6791 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6581; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6794 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6584; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6797 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6587; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6800 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6590; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6803 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6593; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6806 = LUT_mem_MPORT_47_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6596; // @[lut_35.scala 981:74 lut_35.scala 216:26]
  wire  _GEN_6807 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6597; // @[lut_35.scala 943:74 lut_35.scala 944:38]
  wire  _GEN_6808 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6598; // @[lut_35.scala 943:74 lut_35.scala 945:38]
  wire  _GEN_6809 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6599; // @[lut_35.scala 943:74 lut_35.scala 946:38]
  wire  _GEN_6810 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6600; // @[lut_35.scala 943:74 lut_35.scala 947:38]
  wire  _GEN_6811 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6601; // @[lut_35.scala 943:74 lut_35.scala 948:38]
  wire  _GEN_6812 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6602; // @[lut_35.scala 943:74 lut_35.scala 949:38]
  wire  _GEN_6813 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6603; // @[lut_35.scala 943:74 lut_35.scala 950:38]
  wire  _GEN_6814 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6604; // @[lut_35.scala 943:74 lut_35.scala 951:38]
  wire  _GEN_6815 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6605; // @[lut_35.scala 943:74 lut_35.scala 952:38]
  wire  _GEN_6816 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6606; // @[lut_35.scala 943:74 lut_35.scala 953:38]
  wire  _GEN_6817 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6607; // @[lut_35.scala 943:74 lut_35.scala 954:39]
  wire  _GEN_6818 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid | _GEN_6608; // @[lut_35.scala 943:74 lut_35.scala 955:39]
  wire  _GEN_6819 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6609; // @[lut_35.scala 943:74 lut_35.scala 956:39]
  wire  _GEN_6820 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6610; // @[lut_35.scala 943:74 lut_35.scala 957:39]
  wire  _GEN_6821 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6611; // @[lut_35.scala 943:74 lut_35.scala 958:39]
  wire  _GEN_6822 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6612; // @[lut_35.scala 943:74 lut_35.scala 959:39]
  wire  _GEN_6823 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6613; // @[lut_35.scala 943:74 lut_35.scala 960:39]
  wire  _GEN_6824 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6614; // @[lut_35.scala 943:74 lut_35.scala 961:39]
  wire  _GEN_6825 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6615; // @[lut_35.scala 943:74 lut_35.scala 962:39]
  wire  _GEN_6826 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6616; // @[lut_35.scala 943:74 lut_35.scala 963:39]
  wire  _GEN_6827 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6617; // @[lut_35.scala 943:74 lut_35.scala 964:39]
  wire  _GEN_6828 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6618; // @[lut_35.scala 943:74 lut_35.scala 965:39]
  wire  _GEN_6829 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6619; // @[lut_35.scala 943:74 lut_35.scala 966:39]
  wire  _GEN_6830 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6620; // @[lut_35.scala 943:74 lut_35.scala 967:39]
  wire  _GEN_6831 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6621; // @[lut_35.scala 943:74 lut_35.scala 968:39]
  wire  _GEN_6832 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6622; // @[lut_35.scala 943:74 lut_35.scala 969:39]
  wire  _GEN_6833 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6623; // @[lut_35.scala 943:74 lut_35.scala 970:39]
  wire  _GEN_6834 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6624; // @[lut_35.scala 943:74 lut_35.scala 971:39]
  wire  _GEN_6835 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6625; // @[lut_35.scala 943:74 lut_35.scala 972:39]
  wire  _GEN_6836 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6626; // @[lut_35.scala 943:74 lut_35.scala 973:39]
  wire  _GEN_6837 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6627; // @[lut_35.scala 943:74 lut_35.scala 974:39]
  wire  _GEN_6838 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6628; // @[lut_35.scala 943:74 lut_35.scala 975:39]
  wire  _GEN_6839 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6629; // @[lut_35.scala 943:74 lut_35.scala 976:39]
  wire  _GEN_6840 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6630; // @[lut_35.scala 943:74 lut_35.scala 977:39]
  wire  _GEN_6841 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6631; // @[lut_35.scala 943:74 lut_35.scala 978:39]
  wire  _GEN_6842 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid | _GEN_6632; // @[lut_35.scala 943:74 lut_35.scala 979:34]
  wire  _GEN_6846 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 943:74 lut_35.scala 216:26 lut_35.scala 981:27]
  wire  _GEN_6849 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6636; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6852 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6639; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6855 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6642; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6858 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6645; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6861 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6648; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6864 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6651; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6867 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6654; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6870 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6657; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6873 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6660; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6876 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6663; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6879 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6666; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6882 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6669; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6885 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6672; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6888 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6675; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6891 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6678; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6894 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6681; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6897 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6684; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6900 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6687; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6903 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6690; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6906 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6693; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6909 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6696; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6912 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6699; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6915 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6702; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire [5:0] _GEN_6916 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? push_mem_temp : _GEN_6703; // @[lut_35.scala 943:74 lut_35.scala 521:39]
  wire [31:0] _GEN_6917 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? push_id_temp : _GEN_6704; // @[lut_35.scala 943:74 lut_35.scala 522:39]
  wire  _GEN_6920 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6707; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6923 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6710; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6926 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6713; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6929 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6716; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6932 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6719; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6935 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6722; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6938 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6725; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6941 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6728; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6944 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6731; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6947 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6734; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6950 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6737; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6953 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6740; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6956 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6743; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6959 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6746; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6962 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6749; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6965 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6752; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6968 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6755; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6971 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6758; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6974 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6761; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6977 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6764; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6980 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6767; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6983 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6770; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6986 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6773; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6989 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6776; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6992 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6779; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6995 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6782; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_6998 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6785; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_7001 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6788; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_7004 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6791; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_7007 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6794; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_7010 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6797; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_7013 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6800; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_7016 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6803; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_7019 = LUT_mem_MPORT_46_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6806; // @[lut_35.scala 943:74 lut_35.scala 216:26]
  wire  _GEN_7020 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6807; // @[lut_35.scala 905:74 lut_35.scala 906:38]
  wire  _GEN_7021 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6808; // @[lut_35.scala 905:74 lut_35.scala 907:38]
  wire  _GEN_7022 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6809; // @[lut_35.scala 905:74 lut_35.scala 908:38]
  wire  _GEN_7023 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6810; // @[lut_35.scala 905:74 lut_35.scala 909:38]
  wire  _GEN_7024 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6811; // @[lut_35.scala 905:74 lut_35.scala 910:38]
  wire  _GEN_7025 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6812; // @[lut_35.scala 905:74 lut_35.scala 911:38]
  wire  _GEN_7026 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6813; // @[lut_35.scala 905:74 lut_35.scala 912:38]
  wire  _GEN_7027 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6814; // @[lut_35.scala 905:74 lut_35.scala 913:38]
  wire  _GEN_7028 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6815; // @[lut_35.scala 905:74 lut_35.scala 914:38]
  wire  _GEN_7029 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6816; // @[lut_35.scala 905:74 lut_35.scala 915:38]
  wire  _GEN_7030 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid | _GEN_6817; // @[lut_35.scala 905:74 lut_35.scala 916:39]
  wire  _GEN_7031 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6818; // @[lut_35.scala 905:74 lut_35.scala 917:39]
  wire  _GEN_7032 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6819; // @[lut_35.scala 905:74 lut_35.scala 918:39]
  wire  _GEN_7033 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6820; // @[lut_35.scala 905:74 lut_35.scala 919:39]
  wire  _GEN_7034 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6821; // @[lut_35.scala 905:74 lut_35.scala 920:39]
  wire  _GEN_7035 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6822; // @[lut_35.scala 905:74 lut_35.scala 921:39]
  wire  _GEN_7036 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6823; // @[lut_35.scala 905:74 lut_35.scala 922:39]
  wire  _GEN_7037 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6824; // @[lut_35.scala 905:74 lut_35.scala 923:39]
  wire  _GEN_7038 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6825; // @[lut_35.scala 905:74 lut_35.scala 924:39]
  wire  _GEN_7039 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6826; // @[lut_35.scala 905:74 lut_35.scala 925:39]
  wire  _GEN_7040 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6827; // @[lut_35.scala 905:74 lut_35.scala 926:39]
  wire  _GEN_7041 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6828; // @[lut_35.scala 905:74 lut_35.scala 927:39]
  wire  _GEN_7042 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6829; // @[lut_35.scala 905:74 lut_35.scala 928:39]
  wire  _GEN_7043 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6830; // @[lut_35.scala 905:74 lut_35.scala 929:39]
  wire  _GEN_7044 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6831; // @[lut_35.scala 905:74 lut_35.scala 930:39]
  wire  _GEN_7045 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6832; // @[lut_35.scala 905:74 lut_35.scala 931:39]
  wire  _GEN_7046 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6833; // @[lut_35.scala 905:74 lut_35.scala 932:39]
  wire  _GEN_7047 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6834; // @[lut_35.scala 905:74 lut_35.scala 933:39]
  wire  _GEN_7048 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6835; // @[lut_35.scala 905:74 lut_35.scala 934:39]
  wire  _GEN_7049 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6836; // @[lut_35.scala 905:74 lut_35.scala 935:39]
  wire  _GEN_7050 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6837; // @[lut_35.scala 905:74 lut_35.scala 936:39]
  wire  _GEN_7051 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6838; // @[lut_35.scala 905:74 lut_35.scala 937:39]
  wire  _GEN_7052 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6839; // @[lut_35.scala 905:74 lut_35.scala 938:39]
  wire  _GEN_7053 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6840; // @[lut_35.scala 905:74 lut_35.scala 939:39]
  wire  _GEN_7054 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6841; // @[lut_35.scala 905:74 lut_35.scala 940:39]
  wire  _GEN_7055 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid | _GEN_6842; // @[lut_35.scala 905:74 lut_35.scala 941:34]
  wire  _GEN_7059 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 905:74 lut_35.scala 216:26 lut_35.scala 943:27]
  wire  _GEN_7062 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6846; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7065 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6849; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7068 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6852; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7071 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6855; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7074 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6858; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7077 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6861; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7080 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6864; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7083 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6867; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7086 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6870; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7089 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6873; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7092 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6876; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7095 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6879; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7098 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6882; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7101 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6885; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7104 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6888; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7107 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6891; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7110 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6894; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7113 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6897; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7116 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6900; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7119 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6903; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7122 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6906; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7125 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6909; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7128 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6912; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7131 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6915; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire [5:0] _GEN_7132 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? push_mem_temp : _GEN_6916; // @[lut_35.scala 905:74 lut_35.scala 521:39]
  wire [31:0] _GEN_7133 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? push_id_temp : _GEN_6917; // @[lut_35.scala 905:74 lut_35.scala 522:39]
  wire  _GEN_7136 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6920; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7139 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6923; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7142 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6926; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7145 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6929; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7148 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6932; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7151 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6935; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7154 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6938; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7157 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6941; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7160 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6944; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7163 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6947; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7166 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6950; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7169 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6953; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7172 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6956; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7175 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6959; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7178 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6962; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7181 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6965; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7184 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6968; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7187 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6971; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7190 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6974; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7193 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6977; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7196 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6980; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7199 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6983; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7202 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6986; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7205 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6989; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7208 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6992; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7211 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6995; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7214 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6998; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7217 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7001; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7220 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7004; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7223 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7007; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7226 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7010; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7229 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7013; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7232 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7016; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7235 = LUT_mem_MPORT_45_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7019; // @[lut_35.scala 905:74 lut_35.scala 216:26]
  wire  _GEN_7236 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7020; // @[lut_35.scala 867:73 lut_35.scala 868:38]
  wire  _GEN_7237 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7021; // @[lut_35.scala 867:73 lut_35.scala 869:38]
  wire  _GEN_7238 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7022; // @[lut_35.scala 867:73 lut_35.scala 870:38]
  wire  _GEN_7239 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7023; // @[lut_35.scala 867:73 lut_35.scala 871:38]
  wire  _GEN_7240 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7024; // @[lut_35.scala 867:73 lut_35.scala 872:38]
  wire  _GEN_7241 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7025; // @[lut_35.scala 867:73 lut_35.scala 873:38]
  wire  _GEN_7242 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7026; // @[lut_35.scala 867:73 lut_35.scala 874:38]
  wire  _GEN_7243 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7027; // @[lut_35.scala 867:73 lut_35.scala 875:38]
  wire  _GEN_7244 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7028; // @[lut_35.scala 867:73 lut_35.scala 876:38]
  wire  _GEN_7245 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid | _GEN_7029; // @[lut_35.scala 867:73 lut_35.scala 877:38]
  wire  _GEN_7246 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7030; // @[lut_35.scala 867:73 lut_35.scala 878:39]
  wire  _GEN_7247 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7031; // @[lut_35.scala 867:73 lut_35.scala 879:39]
  wire  _GEN_7248 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7032; // @[lut_35.scala 867:73 lut_35.scala 880:39]
  wire  _GEN_7249 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7033; // @[lut_35.scala 867:73 lut_35.scala 881:39]
  wire  _GEN_7250 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7034; // @[lut_35.scala 867:73 lut_35.scala 882:39]
  wire  _GEN_7251 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7035; // @[lut_35.scala 867:73 lut_35.scala 883:39]
  wire  _GEN_7252 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7036; // @[lut_35.scala 867:73 lut_35.scala 884:39]
  wire  _GEN_7253 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7037; // @[lut_35.scala 867:73 lut_35.scala 885:39]
  wire  _GEN_7254 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7038; // @[lut_35.scala 867:73 lut_35.scala 886:39]
  wire  _GEN_7255 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7039; // @[lut_35.scala 867:73 lut_35.scala 887:39]
  wire  _GEN_7256 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7040; // @[lut_35.scala 867:73 lut_35.scala 888:39]
  wire  _GEN_7257 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7041; // @[lut_35.scala 867:73 lut_35.scala 889:39]
  wire  _GEN_7258 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7042; // @[lut_35.scala 867:73 lut_35.scala 890:39]
  wire  _GEN_7259 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7043; // @[lut_35.scala 867:73 lut_35.scala 891:39]
  wire  _GEN_7260 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7044; // @[lut_35.scala 867:73 lut_35.scala 892:39]
  wire  _GEN_7261 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7045; // @[lut_35.scala 867:73 lut_35.scala 893:39]
  wire  _GEN_7262 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7046; // @[lut_35.scala 867:73 lut_35.scala 894:39]
  wire  _GEN_7263 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7047; // @[lut_35.scala 867:73 lut_35.scala 895:39]
  wire  _GEN_7264 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7048; // @[lut_35.scala 867:73 lut_35.scala 896:39]
  wire  _GEN_7265 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7049; // @[lut_35.scala 867:73 lut_35.scala 897:39]
  wire  _GEN_7266 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7050; // @[lut_35.scala 867:73 lut_35.scala 898:39]
  wire  _GEN_7267 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7051; // @[lut_35.scala 867:73 lut_35.scala 899:39]
  wire  _GEN_7268 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7052; // @[lut_35.scala 867:73 lut_35.scala 900:39]
  wire  _GEN_7269 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7053; // @[lut_35.scala 867:73 lut_35.scala 901:39]
  wire  _GEN_7270 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7054; // @[lut_35.scala 867:73 lut_35.scala 902:39]
  wire  _GEN_7271 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid | _GEN_7055; // @[lut_35.scala 867:73 lut_35.scala 903:34]
  wire  _GEN_7275 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 867:73 lut_35.scala 216:26 lut_35.scala 905:27]
  wire  _GEN_7278 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7059; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7281 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7062; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7284 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7065; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7287 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7068; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7290 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7071; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7293 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7074; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7296 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7077; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7299 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7080; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7302 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7083; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7305 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7086; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7308 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7089; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7311 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7092; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7314 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7095; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7317 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7098; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7320 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7101; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7323 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7104; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7326 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7107; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7329 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7110; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7332 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7113; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7335 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7116; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7338 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7119; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7341 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7122; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7344 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7125; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7347 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7128; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7350 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7131; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire [5:0] _GEN_7351 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? push_mem_temp : _GEN_7132; // @[lut_35.scala 867:73 lut_35.scala 521:39]
  wire [31:0] _GEN_7352 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? push_id_temp : _GEN_7133; // @[lut_35.scala 867:73 lut_35.scala 522:39]
  wire  _GEN_7355 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7136; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7358 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7139; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7361 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7142; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7364 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7145; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7367 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7148; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7370 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7151; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7373 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7154; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7376 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7157; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7379 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7160; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7382 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7163; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7385 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7166; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7388 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7169; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7391 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7172; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7394 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7175; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7397 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7178; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7400 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7181; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7403 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7184; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7406 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7187; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7409 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7190; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7412 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7193; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7415 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7196; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7418 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7199; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7421 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7202; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7424 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7205; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7427 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7208; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7430 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7211; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7433 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7214; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7436 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7217; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7439 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7220; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7442 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7223; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7445 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7226; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7448 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7229; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7451 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7232; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7454 = LUT_mem_MPORT_44_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7235; // @[lut_35.scala 867:73 lut_35.scala 216:26]
  wire  _GEN_7455 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7236; // @[lut_35.scala 829:73 lut_35.scala 830:38]
  wire  _GEN_7456 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7237; // @[lut_35.scala 829:73 lut_35.scala 831:38]
  wire  _GEN_7457 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7238; // @[lut_35.scala 829:73 lut_35.scala 832:38]
  wire  _GEN_7458 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7239; // @[lut_35.scala 829:73 lut_35.scala 833:38]
  wire  _GEN_7459 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7240; // @[lut_35.scala 829:73 lut_35.scala 834:38]
  wire  _GEN_7460 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7241; // @[lut_35.scala 829:73 lut_35.scala 835:38]
  wire  _GEN_7461 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7242; // @[lut_35.scala 829:73 lut_35.scala 836:38]
  wire  _GEN_7462 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7243; // @[lut_35.scala 829:73 lut_35.scala 837:38]
  wire  _GEN_7463 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid | _GEN_7244; // @[lut_35.scala 829:73 lut_35.scala 838:38]
  wire  _GEN_7464 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7245; // @[lut_35.scala 829:73 lut_35.scala 839:38]
  wire  _GEN_7465 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7246; // @[lut_35.scala 829:73 lut_35.scala 840:39]
  wire  _GEN_7466 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7247; // @[lut_35.scala 829:73 lut_35.scala 841:39]
  wire  _GEN_7467 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7248; // @[lut_35.scala 829:73 lut_35.scala 842:39]
  wire  _GEN_7468 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7249; // @[lut_35.scala 829:73 lut_35.scala 843:39]
  wire  _GEN_7469 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7250; // @[lut_35.scala 829:73 lut_35.scala 844:39]
  wire  _GEN_7470 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7251; // @[lut_35.scala 829:73 lut_35.scala 845:39]
  wire  _GEN_7471 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7252; // @[lut_35.scala 829:73 lut_35.scala 846:39]
  wire  _GEN_7472 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7253; // @[lut_35.scala 829:73 lut_35.scala 847:39]
  wire  _GEN_7473 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7254; // @[lut_35.scala 829:73 lut_35.scala 848:39]
  wire  _GEN_7474 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7255; // @[lut_35.scala 829:73 lut_35.scala 849:39]
  wire  _GEN_7475 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7256; // @[lut_35.scala 829:73 lut_35.scala 850:39]
  wire  _GEN_7476 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7257; // @[lut_35.scala 829:73 lut_35.scala 851:39]
  wire  _GEN_7477 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7258; // @[lut_35.scala 829:73 lut_35.scala 852:39]
  wire  _GEN_7478 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7259; // @[lut_35.scala 829:73 lut_35.scala 853:39]
  wire  _GEN_7479 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7260; // @[lut_35.scala 829:73 lut_35.scala 854:39]
  wire  _GEN_7480 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7261; // @[lut_35.scala 829:73 lut_35.scala 855:39]
  wire  _GEN_7481 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7262; // @[lut_35.scala 829:73 lut_35.scala 856:39]
  wire  _GEN_7482 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7263; // @[lut_35.scala 829:73 lut_35.scala 857:39]
  wire  _GEN_7483 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7264; // @[lut_35.scala 829:73 lut_35.scala 858:39]
  wire  _GEN_7484 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7265; // @[lut_35.scala 829:73 lut_35.scala 859:39]
  wire  _GEN_7485 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7266; // @[lut_35.scala 829:73 lut_35.scala 860:39]
  wire  _GEN_7486 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7267; // @[lut_35.scala 829:73 lut_35.scala 861:39]
  wire  _GEN_7487 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7268; // @[lut_35.scala 829:73 lut_35.scala 862:39]
  wire  _GEN_7488 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7269; // @[lut_35.scala 829:73 lut_35.scala 863:39]
  wire  _GEN_7489 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7270; // @[lut_35.scala 829:73 lut_35.scala 864:39]
  wire  _GEN_7490 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid | _GEN_7271; // @[lut_35.scala 829:73 lut_35.scala 865:34]
  wire  _GEN_7494 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 829:73 lut_35.scala 216:26 lut_35.scala 867:27]
  wire  _GEN_7497 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7275; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7500 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7278; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7503 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7281; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7506 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7284; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7509 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7287; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7512 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7290; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7515 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7293; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7518 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7296; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7521 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7299; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7524 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7302; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7527 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7305; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7530 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7308; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7533 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7311; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7536 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7314; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7539 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7317; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7542 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7320; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7545 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7323; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7548 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7326; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7551 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7329; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7554 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7332; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7557 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7335; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7560 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7338; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7563 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7341; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7566 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7344; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7569 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7347; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7572 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7350; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire [5:0] _GEN_7573 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? push_mem_temp : _GEN_7351; // @[lut_35.scala 829:73 lut_35.scala 521:39]
  wire [31:0] _GEN_7574 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? push_id_temp : _GEN_7352; // @[lut_35.scala 829:73 lut_35.scala 522:39]
  wire  _GEN_7577 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7355; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7580 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7358; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7583 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7361; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7586 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7364; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7589 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7367; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7592 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7370; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7595 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7373; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7598 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7376; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7601 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7379; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7604 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7382; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7607 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7385; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7610 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7388; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7613 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7391; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7616 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7394; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7619 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7397; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7622 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7400; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7625 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7403; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7628 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7406; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7631 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7409; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7634 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7412; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7637 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7415; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7640 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7418; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7643 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7421; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7646 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7424; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7649 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7427; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7652 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7430; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7655 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7433; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7658 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7436; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7661 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7439; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7664 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7442; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7667 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7445; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7670 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7448; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7673 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7451; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7676 = LUT_mem_MPORT_43_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7454; // @[lut_35.scala 829:73 lut_35.scala 216:26]
  wire  _GEN_7677 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7455; // @[lut_35.scala 791:73 lut_35.scala 792:38]
  wire  _GEN_7678 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7456; // @[lut_35.scala 791:73 lut_35.scala 793:38]
  wire  _GEN_7679 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7457; // @[lut_35.scala 791:73 lut_35.scala 794:38]
  wire  _GEN_7680 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7458; // @[lut_35.scala 791:73 lut_35.scala 795:38]
  wire  _GEN_7681 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7459; // @[lut_35.scala 791:73 lut_35.scala 796:38]
  wire  _GEN_7682 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7460; // @[lut_35.scala 791:73 lut_35.scala 797:38]
  wire  _GEN_7683 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7461; // @[lut_35.scala 791:73 lut_35.scala 798:38]
  wire  _GEN_7684 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid | _GEN_7462; // @[lut_35.scala 791:73 lut_35.scala 799:38]
  wire  _GEN_7685 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7463; // @[lut_35.scala 791:73 lut_35.scala 800:38]
  wire  _GEN_7686 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7464; // @[lut_35.scala 791:73 lut_35.scala 801:38]
  wire  _GEN_7687 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7465; // @[lut_35.scala 791:73 lut_35.scala 802:39]
  wire  _GEN_7688 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7466; // @[lut_35.scala 791:73 lut_35.scala 803:39]
  wire  _GEN_7689 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7467; // @[lut_35.scala 791:73 lut_35.scala 804:39]
  wire  _GEN_7690 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7468; // @[lut_35.scala 791:73 lut_35.scala 805:39]
  wire  _GEN_7691 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7469; // @[lut_35.scala 791:73 lut_35.scala 806:39]
  wire  _GEN_7692 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7470; // @[lut_35.scala 791:73 lut_35.scala 807:39]
  wire  _GEN_7693 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7471; // @[lut_35.scala 791:73 lut_35.scala 808:39]
  wire  _GEN_7694 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7472; // @[lut_35.scala 791:73 lut_35.scala 809:39]
  wire  _GEN_7695 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7473; // @[lut_35.scala 791:73 lut_35.scala 810:39]
  wire  _GEN_7696 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7474; // @[lut_35.scala 791:73 lut_35.scala 811:39]
  wire  _GEN_7697 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7475; // @[lut_35.scala 791:73 lut_35.scala 812:39]
  wire  _GEN_7698 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7476; // @[lut_35.scala 791:73 lut_35.scala 813:39]
  wire  _GEN_7699 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7477; // @[lut_35.scala 791:73 lut_35.scala 814:39]
  wire  _GEN_7700 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7478; // @[lut_35.scala 791:73 lut_35.scala 815:39]
  wire  _GEN_7701 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7479; // @[lut_35.scala 791:73 lut_35.scala 816:39]
  wire  _GEN_7702 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7480; // @[lut_35.scala 791:73 lut_35.scala 817:39]
  wire  _GEN_7703 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7481; // @[lut_35.scala 791:73 lut_35.scala 818:39]
  wire  _GEN_7704 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7482; // @[lut_35.scala 791:73 lut_35.scala 819:39]
  wire  _GEN_7705 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7483; // @[lut_35.scala 791:73 lut_35.scala 820:39]
  wire  _GEN_7706 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7484; // @[lut_35.scala 791:73 lut_35.scala 821:39]
  wire  _GEN_7707 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7485; // @[lut_35.scala 791:73 lut_35.scala 822:39]
  wire  _GEN_7708 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7486; // @[lut_35.scala 791:73 lut_35.scala 823:39]
  wire  _GEN_7709 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7487; // @[lut_35.scala 791:73 lut_35.scala 824:39]
  wire  _GEN_7710 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7488; // @[lut_35.scala 791:73 lut_35.scala 825:39]
  wire  _GEN_7711 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7489; // @[lut_35.scala 791:73 lut_35.scala 826:39]
  wire  _GEN_7712 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid | _GEN_7490; // @[lut_35.scala 791:73 lut_35.scala 827:34]
  wire  _GEN_7716 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 791:73 lut_35.scala 216:26 lut_35.scala 829:27]
  wire  _GEN_7719 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7494; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7722 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7497; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7725 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7500; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7728 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7503; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7731 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7506; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7734 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7509; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7737 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7512; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7740 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7515; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7743 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7518; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7746 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7521; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7749 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7524; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7752 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7527; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7755 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7530; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7758 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7533; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7761 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7536; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7764 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7539; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7767 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7542; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7770 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7545; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7773 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7548; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7776 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7551; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7779 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7554; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7782 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7557; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7785 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7560; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7788 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7563; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7791 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7566; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7794 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7569; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7797 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7572; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire [5:0] _GEN_7798 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? push_mem_temp : _GEN_7573; // @[lut_35.scala 791:73 lut_35.scala 521:39]
  wire [31:0] _GEN_7799 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? push_id_temp : _GEN_7574; // @[lut_35.scala 791:73 lut_35.scala 522:39]
  wire  _GEN_7802 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7577; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7805 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7580; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7808 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7583; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7811 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7586; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7814 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7589; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7817 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7592; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7820 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7595; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7823 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7598; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7826 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7601; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7829 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7604; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7832 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7607; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7835 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7610; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7838 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7613; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7841 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7616; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7844 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7619; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7847 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7622; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7850 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7625; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7853 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7628; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7856 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7631; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7859 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7634; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7862 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7637; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7865 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7640; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7868 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7643; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7871 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7646; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7874 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7649; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7877 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7652; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7880 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7655; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7883 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7658; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7886 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7661; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7889 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7664; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7892 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7667; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7895 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7670; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7898 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7673; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7901 = LUT_mem_MPORT_42_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7676; // @[lut_35.scala 791:73 lut_35.scala 216:26]
  wire  _GEN_7902 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7677; // @[lut_35.scala 753:73 lut_35.scala 754:38]
  wire  _GEN_7903 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7678; // @[lut_35.scala 753:73 lut_35.scala 755:38]
  wire  _GEN_7904 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7679; // @[lut_35.scala 753:73 lut_35.scala 756:38]
  wire  _GEN_7905 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7680; // @[lut_35.scala 753:73 lut_35.scala 757:38]
  wire  _GEN_7906 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7681; // @[lut_35.scala 753:73 lut_35.scala 758:38]
  wire  _GEN_7907 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7682; // @[lut_35.scala 753:73 lut_35.scala 759:38]
  wire  _GEN_7908 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid | _GEN_7683; // @[lut_35.scala 753:73 lut_35.scala 760:38]
  wire  _GEN_7909 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7684; // @[lut_35.scala 753:73 lut_35.scala 761:38]
  wire  _GEN_7910 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7685; // @[lut_35.scala 753:73 lut_35.scala 762:38]
  wire  _GEN_7911 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7686; // @[lut_35.scala 753:73 lut_35.scala 763:38]
  wire  _GEN_7912 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7687; // @[lut_35.scala 753:73 lut_35.scala 764:39]
  wire  _GEN_7913 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7688; // @[lut_35.scala 753:73 lut_35.scala 765:39]
  wire  _GEN_7914 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7689; // @[lut_35.scala 753:73 lut_35.scala 766:39]
  wire  _GEN_7915 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7690; // @[lut_35.scala 753:73 lut_35.scala 767:39]
  wire  _GEN_7916 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7691; // @[lut_35.scala 753:73 lut_35.scala 768:39]
  wire  _GEN_7917 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7692; // @[lut_35.scala 753:73 lut_35.scala 769:39]
  wire  _GEN_7918 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7693; // @[lut_35.scala 753:73 lut_35.scala 770:39]
  wire  _GEN_7919 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7694; // @[lut_35.scala 753:73 lut_35.scala 771:39]
  wire  _GEN_7920 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7695; // @[lut_35.scala 753:73 lut_35.scala 772:39]
  wire  _GEN_7921 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7696; // @[lut_35.scala 753:73 lut_35.scala 773:39]
  wire  _GEN_7922 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7697; // @[lut_35.scala 753:73 lut_35.scala 774:39]
  wire  _GEN_7923 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7698; // @[lut_35.scala 753:73 lut_35.scala 775:39]
  wire  _GEN_7924 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7699; // @[lut_35.scala 753:73 lut_35.scala 776:39]
  wire  _GEN_7925 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7700; // @[lut_35.scala 753:73 lut_35.scala 777:39]
  wire  _GEN_7926 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7701; // @[lut_35.scala 753:73 lut_35.scala 778:39]
  wire  _GEN_7927 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7702; // @[lut_35.scala 753:73 lut_35.scala 779:39]
  wire  _GEN_7928 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7703; // @[lut_35.scala 753:73 lut_35.scala 780:39]
  wire  _GEN_7929 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7704; // @[lut_35.scala 753:73 lut_35.scala 781:39]
  wire  _GEN_7930 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7705; // @[lut_35.scala 753:73 lut_35.scala 782:39]
  wire  _GEN_7931 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7706; // @[lut_35.scala 753:73 lut_35.scala 783:39]
  wire  _GEN_7932 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7707; // @[lut_35.scala 753:73 lut_35.scala 784:39]
  wire  _GEN_7933 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7708; // @[lut_35.scala 753:73 lut_35.scala 785:39]
  wire  _GEN_7934 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7709; // @[lut_35.scala 753:73 lut_35.scala 786:39]
  wire  _GEN_7935 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7710; // @[lut_35.scala 753:73 lut_35.scala 787:39]
  wire  _GEN_7936 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7711; // @[lut_35.scala 753:73 lut_35.scala 788:39]
  wire  _GEN_7937 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid | _GEN_7712; // @[lut_35.scala 753:73 lut_35.scala 789:34]
  wire  _GEN_7941 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 753:73 lut_35.scala 216:26 lut_35.scala 791:27]
  wire  _GEN_7944 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7716; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_7947 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7719; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_7950 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7722; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_7953 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7725; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_7956 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7728; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_7959 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7731; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_7962 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7734; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_7965 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7737; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_7968 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7740; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_7971 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7743; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_7974 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7746; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_7977 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7749; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_7980 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7752; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_7983 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7755; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_7986 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7758; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_7989 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7761; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_7992 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7764; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_7995 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7767; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_7998 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7770; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8001 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7773; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8004 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7776; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8007 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7779; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8010 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7782; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8013 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7785; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8016 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7788; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8019 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7791; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8022 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7794; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8025 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7797; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire [5:0] _GEN_8026 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? push_mem_temp : _GEN_7798; // @[lut_35.scala 753:73 lut_35.scala 521:39]
  wire [31:0] _GEN_8027 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? push_id_temp : _GEN_7799; // @[lut_35.scala 753:73 lut_35.scala 522:39]
  wire  _GEN_8030 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7802; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8033 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7805; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8036 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7808; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8039 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7811; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8042 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7814; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8045 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7817; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8048 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7820; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8051 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7823; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8054 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7826; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8057 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7829; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8060 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7832; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8063 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7835; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8066 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7838; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8069 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7841; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8072 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7844; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8075 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7847; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8078 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7850; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8081 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7853; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8084 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7856; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8087 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7859; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8090 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7862; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8093 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7865; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8096 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7868; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8099 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7871; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8102 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7874; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8105 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7877; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8108 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7880; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8111 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7883; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8114 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7886; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8117 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7889; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8120 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7892; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8123 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7895; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8126 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7898; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8129 = LUT_mem_MPORT_41_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7901; // @[lut_35.scala 753:73 lut_35.scala 216:26]
  wire  _GEN_8130 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7902; // @[lut_35.scala 715:73 lut_35.scala 716:38]
  wire  _GEN_8131 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7903; // @[lut_35.scala 715:73 lut_35.scala 717:38]
  wire  _GEN_8132 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7904; // @[lut_35.scala 715:73 lut_35.scala 718:38]
  wire  _GEN_8133 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7905; // @[lut_35.scala 715:73 lut_35.scala 719:38]
  wire  _GEN_8134 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7906; // @[lut_35.scala 715:73 lut_35.scala 720:38]
  wire  _GEN_8135 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid | _GEN_7907; // @[lut_35.scala 715:73 lut_35.scala 721:38]
  wire  _GEN_8136 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7908; // @[lut_35.scala 715:73 lut_35.scala 722:38]
  wire  _GEN_8137 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7909; // @[lut_35.scala 715:73 lut_35.scala 723:38]
  wire  _GEN_8138 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7910; // @[lut_35.scala 715:73 lut_35.scala 724:38]
  wire  _GEN_8139 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7911; // @[lut_35.scala 715:73 lut_35.scala 725:38]
  wire  _GEN_8140 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7912; // @[lut_35.scala 715:73 lut_35.scala 726:39]
  wire  _GEN_8141 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7913; // @[lut_35.scala 715:73 lut_35.scala 727:39]
  wire  _GEN_8142 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7914; // @[lut_35.scala 715:73 lut_35.scala 728:39]
  wire  _GEN_8143 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7915; // @[lut_35.scala 715:73 lut_35.scala 729:39]
  wire  _GEN_8144 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7916; // @[lut_35.scala 715:73 lut_35.scala 730:39]
  wire  _GEN_8145 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7917; // @[lut_35.scala 715:73 lut_35.scala 731:39]
  wire  _GEN_8146 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7918; // @[lut_35.scala 715:73 lut_35.scala 732:39]
  wire  _GEN_8147 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7919; // @[lut_35.scala 715:73 lut_35.scala 733:39]
  wire  _GEN_8148 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7920; // @[lut_35.scala 715:73 lut_35.scala 734:39]
  wire  _GEN_8149 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7921; // @[lut_35.scala 715:73 lut_35.scala 735:39]
  wire  _GEN_8150 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7922; // @[lut_35.scala 715:73 lut_35.scala 736:39]
  wire  _GEN_8151 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7923; // @[lut_35.scala 715:73 lut_35.scala 737:39]
  wire  _GEN_8152 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7924; // @[lut_35.scala 715:73 lut_35.scala 738:39]
  wire  _GEN_8153 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7925; // @[lut_35.scala 715:73 lut_35.scala 739:39]
  wire  _GEN_8154 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7926; // @[lut_35.scala 715:73 lut_35.scala 740:39]
  wire  _GEN_8155 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7927; // @[lut_35.scala 715:73 lut_35.scala 741:39]
  wire  _GEN_8156 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7928; // @[lut_35.scala 715:73 lut_35.scala 742:39]
  wire  _GEN_8157 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7929; // @[lut_35.scala 715:73 lut_35.scala 743:39]
  wire  _GEN_8158 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7930; // @[lut_35.scala 715:73 lut_35.scala 744:39]
  wire  _GEN_8159 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7931; // @[lut_35.scala 715:73 lut_35.scala 745:39]
  wire  _GEN_8160 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7932; // @[lut_35.scala 715:73 lut_35.scala 746:39]
  wire  _GEN_8161 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7933; // @[lut_35.scala 715:73 lut_35.scala 747:39]
  wire  _GEN_8162 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7934; // @[lut_35.scala 715:73 lut_35.scala 748:39]
  wire  _GEN_8163 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7935; // @[lut_35.scala 715:73 lut_35.scala 749:39]
  wire  _GEN_8164 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7936; // @[lut_35.scala 715:73 lut_35.scala 750:39]
  wire  _GEN_8165 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid | _GEN_7937; // @[lut_35.scala 715:73 lut_35.scala 751:34]
  wire  _GEN_8169 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 715:73 lut_35.scala 216:26 lut_35.scala 753:27]
  wire  _GEN_8172 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7941; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8175 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7944; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8178 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7947; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8181 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7950; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8184 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7953; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8187 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7956; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8190 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7959; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8193 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7962; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8196 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7965; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8199 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7968; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8202 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7971; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8205 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7974; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8208 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7977; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8211 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7980; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8214 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7983; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8217 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7986; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8220 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7989; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8223 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7992; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8226 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7995; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8229 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7998; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8232 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8001; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8235 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8004; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8238 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8007; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8241 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8010; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8244 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8013; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8247 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8016; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8250 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8019; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8253 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8022; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8256 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8025; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire [5:0] _GEN_8257 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? push_mem_temp : _GEN_8026; // @[lut_35.scala 715:73 lut_35.scala 521:39]
  wire [31:0] _GEN_8258 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? push_id_temp : _GEN_8027; // @[lut_35.scala 715:73 lut_35.scala 522:39]
  wire  _GEN_8261 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8030; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8264 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8033; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8267 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8036; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8270 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8039; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8273 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8042; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8276 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8045; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8279 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8048; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8282 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8051; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8285 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8054; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8288 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8057; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8291 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8060; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8294 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8063; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8297 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8066; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8300 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8069; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8303 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8072; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8306 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8075; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8309 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8078; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8312 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8081; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8315 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8084; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8318 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8087; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8321 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8090; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8324 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8093; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8327 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8096; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8330 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8099; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8333 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8102; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8336 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8105; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8339 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8108; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8342 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8111; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8345 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8114; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8348 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8117; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8351 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8120; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8354 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8123; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8357 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8126; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8360 = LUT_mem_MPORT_40_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8129; // @[lut_35.scala 715:73 lut_35.scala 216:26]
  wire  _GEN_8361 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8130; // @[lut_35.scala 677:73 lut_35.scala 678:38]
  wire  _GEN_8362 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8131; // @[lut_35.scala 677:73 lut_35.scala 679:38]
  wire  _GEN_8363 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8132; // @[lut_35.scala 677:73 lut_35.scala 680:38]
  wire  _GEN_8364 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8133; // @[lut_35.scala 677:73 lut_35.scala 681:38]
  wire  _GEN_8365 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid | _GEN_8134; // @[lut_35.scala 677:73 lut_35.scala 682:38]
  wire  _GEN_8366 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8135; // @[lut_35.scala 677:73 lut_35.scala 683:38]
  wire  _GEN_8367 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8136; // @[lut_35.scala 677:73 lut_35.scala 684:38]
  wire  _GEN_8368 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8137; // @[lut_35.scala 677:73 lut_35.scala 685:38]
  wire  _GEN_8369 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8138; // @[lut_35.scala 677:73 lut_35.scala 686:38]
  wire  _GEN_8370 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8139; // @[lut_35.scala 677:73 lut_35.scala 687:38]
  wire  _GEN_8371 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8140; // @[lut_35.scala 677:73 lut_35.scala 688:39]
  wire  _GEN_8372 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8141; // @[lut_35.scala 677:73 lut_35.scala 689:39]
  wire  _GEN_8373 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8142; // @[lut_35.scala 677:73 lut_35.scala 690:39]
  wire  _GEN_8374 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8143; // @[lut_35.scala 677:73 lut_35.scala 691:39]
  wire  _GEN_8375 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8144; // @[lut_35.scala 677:73 lut_35.scala 692:39]
  wire  _GEN_8376 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8145; // @[lut_35.scala 677:73 lut_35.scala 693:39]
  wire  _GEN_8377 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8146; // @[lut_35.scala 677:73 lut_35.scala 694:39]
  wire  _GEN_8378 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8147; // @[lut_35.scala 677:73 lut_35.scala 695:39]
  wire  _GEN_8379 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8148; // @[lut_35.scala 677:73 lut_35.scala 696:39]
  wire  _GEN_8380 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8149; // @[lut_35.scala 677:73 lut_35.scala 697:39]
  wire  _GEN_8381 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8150; // @[lut_35.scala 677:73 lut_35.scala 698:39]
  wire  _GEN_8382 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8151; // @[lut_35.scala 677:73 lut_35.scala 699:39]
  wire  _GEN_8383 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8152; // @[lut_35.scala 677:73 lut_35.scala 700:39]
  wire  _GEN_8384 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8153; // @[lut_35.scala 677:73 lut_35.scala 701:39]
  wire  _GEN_8385 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8154; // @[lut_35.scala 677:73 lut_35.scala 702:39]
  wire  _GEN_8386 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8155; // @[lut_35.scala 677:73 lut_35.scala 703:39]
  wire  _GEN_8387 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8156; // @[lut_35.scala 677:73 lut_35.scala 704:39]
  wire  _GEN_8388 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8157; // @[lut_35.scala 677:73 lut_35.scala 705:39]
  wire  _GEN_8389 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8158; // @[lut_35.scala 677:73 lut_35.scala 706:39]
  wire  _GEN_8390 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8159; // @[lut_35.scala 677:73 lut_35.scala 707:39]
  wire  _GEN_8391 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8160; // @[lut_35.scala 677:73 lut_35.scala 708:39]
  wire  _GEN_8392 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8161; // @[lut_35.scala 677:73 lut_35.scala 709:39]
  wire  _GEN_8393 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8162; // @[lut_35.scala 677:73 lut_35.scala 710:39]
  wire  _GEN_8394 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8163; // @[lut_35.scala 677:73 lut_35.scala 711:39]
  wire  _GEN_8395 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8164; // @[lut_35.scala 677:73 lut_35.scala 712:39]
  wire  _GEN_8396 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid | _GEN_8165; // @[lut_35.scala 677:73 lut_35.scala 713:34]
  wire  _GEN_8400 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 677:73 lut_35.scala 216:26 lut_35.scala 715:27]
  wire  _GEN_8403 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8169; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8406 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8172; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8409 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8175; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8412 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8178; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8415 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8181; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8418 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8184; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8421 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8187; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8424 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8190; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8427 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8193; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8430 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8196; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8433 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8199; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8436 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8202; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8439 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8205; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8442 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8208; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8445 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8211; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8448 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8214; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8451 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8217; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8454 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8220; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8457 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8223; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8460 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8226; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8463 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8229; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8466 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8232; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8469 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8235; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8472 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8238; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8475 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8241; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8478 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8244; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8481 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8247; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8484 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8250; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8487 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8253; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8490 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8256; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire [5:0] _GEN_8491 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? push_mem_temp : _GEN_8257; // @[lut_35.scala 677:73 lut_35.scala 521:39]
  wire [31:0] _GEN_8492 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? push_id_temp : _GEN_8258; // @[lut_35.scala 677:73 lut_35.scala 522:39]
  wire  _GEN_8495 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8261; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8498 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8264; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8501 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8267; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8504 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8270; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8507 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8273; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8510 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8276; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8513 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8279; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8516 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8282; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8519 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8285; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8522 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8288; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8525 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8291; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8528 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8294; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8531 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8297; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8534 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8300; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8537 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8303; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8540 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8306; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8543 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8309; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8546 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8312; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8549 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8315; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8552 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8318; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8555 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8321; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8558 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8324; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8561 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8327; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8564 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8330; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8567 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8333; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8570 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8336; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8573 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8339; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8576 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8342; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8579 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8345; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8582 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8348; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8585 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8351; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8588 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8354; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8591 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8357; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8594 = LUT_mem_MPORT_39_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8360; // @[lut_35.scala 677:73 lut_35.scala 216:26]
  wire  _GEN_8595 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8361; // @[lut_35.scala 639:73 lut_35.scala 640:38]
  wire  _GEN_8596 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8362; // @[lut_35.scala 639:73 lut_35.scala 641:38]
  wire  _GEN_8597 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8363; // @[lut_35.scala 639:73 lut_35.scala 642:38]
  wire  _GEN_8598 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid | _GEN_8364; // @[lut_35.scala 639:73 lut_35.scala 643:38]
  wire  _GEN_8599 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8365; // @[lut_35.scala 639:73 lut_35.scala 644:38]
  wire  _GEN_8600 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8366; // @[lut_35.scala 639:73 lut_35.scala 645:38]
  wire  _GEN_8601 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8367; // @[lut_35.scala 639:73 lut_35.scala 646:38]
  wire  _GEN_8602 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8368; // @[lut_35.scala 639:73 lut_35.scala 647:38]
  wire  _GEN_8603 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8369; // @[lut_35.scala 639:73 lut_35.scala 648:38]
  wire  _GEN_8604 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8370; // @[lut_35.scala 639:73 lut_35.scala 649:38]
  wire  _GEN_8605 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8371; // @[lut_35.scala 639:73 lut_35.scala 650:39]
  wire  _GEN_8606 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8372; // @[lut_35.scala 639:73 lut_35.scala 651:39]
  wire  _GEN_8607 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8373; // @[lut_35.scala 639:73 lut_35.scala 652:39]
  wire  _GEN_8608 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8374; // @[lut_35.scala 639:73 lut_35.scala 653:39]
  wire  _GEN_8609 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8375; // @[lut_35.scala 639:73 lut_35.scala 654:39]
  wire  _GEN_8610 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8376; // @[lut_35.scala 639:73 lut_35.scala 655:39]
  wire  _GEN_8611 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8377; // @[lut_35.scala 639:73 lut_35.scala 656:39]
  wire  _GEN_8612 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8378; // @[lut_35.scala 639:73 lut_35.scala 657:39]
  wire  _GEN_8613 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8379; // @[lut_35.scala 639:73 lut_35.scala 658:39]
  wire  _GEN_8614 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8380; // @[lut_35.scala 639:73 lut_35.scala 659:39]
  wire  _GEN_8615 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8381; // @[lut_35.scala 639:73 lut_35.scala 660:39]
  wire  _GEN_8616 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8382; // @[lut_35.scala 639:73 lut_35.scala 661:39]
  wire  _GEN_8617 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8383; // @[lut_35.scala 639:73 lut_35.scala 662:39]
  wire  _GEN_8618 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8384; // @[lut_35.scala 639:73 lut_35.scala 663:39]
  wire  _GEN_8619 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8385; // @[lut_35.scala 639:73 lut_35.scala 664:39]
  wire  _GEN_8620 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8386; // @[lut_35.scala 639:73 lut_35.scala 665:39]
  wire  _GEN_8621 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8387; // @[lut_35.scala 639:73 lut_35.scala 666:39]
  wire  _GEN_8622 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8388; // @[lut_35.scala 639:73 lut_35.scala 667:39]
  wire  _GEN_8623 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8389; // @[lut_35.scala 639:73 lut_35.scala 668:39]
  wire  _GEN_8624 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8390; // @[lut_35.scala 639:73 lut_35.scala 669:39]
  wire  _GEN_8625 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8391; // @[lut_35.scala 639:73 lut_35.scala 670:39]
  wire  _GEN_8626 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8392; // @[lut_35.scala 639:73 lut_35.scala 671:39]
  wire  _GEN_8627 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8393; // @[lut_35.scala 639:73 lut_35.scala 672:39]
  wire  _GEN_8628 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8394; // @[lut_35.scala 639:73 lut_35.scala 673:39]
  wire  _GEN_8629 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8395; // @[lut_35.scala 639:73 lut_35.scala 674:39]
  wire  _GEN_8630 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid | _GEN_8396; // @[lut_35.scala 639:73 lut_35.scala 675:34]
  wire  _GEN_8634 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 639:73 lut_35.scala 216:26 lut_35.scala 677:27]
  wire  _GEN_8637 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8400; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8640 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8403; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8643 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8406; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8646 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8409; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8649 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8412; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8652 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8415; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8655 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8418; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8658 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8421; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8661 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8424; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8664 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8427; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8667 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8430; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8670 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8433; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8673 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8436; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8676 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8439; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8679 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8442; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8682 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8445; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8685 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8448; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8688 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8451; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8691 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8454; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8694 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8457; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8697 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8460; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8700 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8463; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8703 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8466; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8706 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8469; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8709 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8472; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8712 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8475; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8715 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8478; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8718 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8481; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8721 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8484; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8724 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8487; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8727 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8490; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire [5:0] _GEN_8728 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? push_mem_temp : _GEN_8491; // @[lut_35.scala 639:73 lut_35.scala 521:39]
  wire [31:0] _GEN_8729 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? push_id_temp : _GEN_8492; // @[lut_35.scala 639:73 lut_35.scala 522:39]
  wire  _GEN_8732 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8495; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8735 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8498; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8738 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8501; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8741 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8504; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8744 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8507; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8747 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8510; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8750 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8513; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8753 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8516; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8756 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8519; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8759 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8522; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8762 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8525; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8765 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8528; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8768 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8531; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8771 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8534; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8774 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8537; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8777 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8540; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8780 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8543; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8783 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8546; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8786 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8549; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8789 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8552; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8792 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8555; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8795 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8558; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8798 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8561; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8801 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8564; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8804 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8567; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8807 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8570; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8810 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8573; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8813 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8576; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8816 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8579; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8819 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8582; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8822 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8585; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8825 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8588; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8828 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8591; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8831 = LUT_mem_MPORT_38_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8594; // @[lut_35.scala 639:73 lut_35.scala 216:26]
  wire  _GEN_8832 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8595; // @[lut_35.scala 601:73 lut_35.scala 602:38]
  wire  _GEN_8833 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8596; // @[lut_35.scala 601:73 lut_35.scala 603:38]
  wire  _GEN_8834 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid | _GEN_8597; // @[lut_35.scala 601:73 lut_35.scala 604:38]
  wire  _GEN_8835 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8598; // @[lut_35.scala 601:73 lut_35.scala 605:38]
  wire  _GEN_8836 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8599; // @[lut_35.scala 601:73 lut_35.scala 606:38]
  wire  _GEN_8837 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8600; // @[lut_35.scala 601:73 lut_35.scala 607:38]
  wire  _GEN_8838 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8601; // @[lut_35.scala 601:73 lut_35.scala 608:38]
  wire  _GEN_8839 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8602; // @[lut_35.scala 601:73 lut_35.scala 609:38]
  wire  _GEN_8840 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8603; // @[lut_35.scala 601:73 lut_35.scala 610:38]
  wire  _GEN_8841 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8604; // @[lut_35.scala 601:73 lut_35.scala 611:38]
  wire  _GEN_8842 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8605; // @[lut_35.scala 601:73 lut_35.scala 612:39]
  wire  _GEN_8843 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8606; // @[lut_35.scala 601:73 lut_35.scala 613:39]
  wire  _GEN_8844 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8607; // @[lut_35.scala 601:73 lut_35.scala 614:39]
  wire  _GEN_8845 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8608; // @[lut_35.scala 601:73 lut_35.scala 615:39]
  wire  _GEN_8846 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8609; // @[lut_35.scala 601:73 lut_35.scala 616:39]
  wire  _GEN_8847 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8610; // @[lut_35.scala 601:73 lut_35.scala 617:39]
  wire  _GEN_8848 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8611; // @[lut_35.scala 601:73 lut_35.scala 618:39]
  wire  _GEN_8849 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8612; // @[lut_35.scala 601:73 lut_35.scala 619:39]
  wire  _GEN_8850 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8613; // @[lut_35.scala 601:73 lut_35.scala 620:39]
  wire  _GEN_8851 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8614; // @[lut_35.scala 601:73 lut_35.scala 621:39]
  wire  _GEN_8852 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8615; // @[lut_35.scala 601:73 lut_35.scala 622:39]
  wire  _GEN_8853 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8616; // @[lut_35.scala 601:73 lut_35.scala 623:39]
  wire  _GEN_8854 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8617; // @[lut_35.scala 601:73 lut_35.scala 624:39]
  wire  _GEN_8855 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8618; // @[lut_35.scala 601:73 lut_35.scala 625:39]
  wire  _GEN_8856 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8619; // @[lut_35.scala 601:73 lut_35.scala 626:39]
  wire  _GEN_8857 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8620; // @[lut_35.scala 601:73 lut_35.scala 627:39]
  wire  _GEN_8858 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8621; // @[lut_35.scala 601:73 lut_35.scala 628:39]
  wire  _GEN_8859 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8622; // @[lut_35.scala 601:73 lut_35.scala 629:39]
  wire  _GEN_8860 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8623; // @[lut_35.scala 601:73 lut_35.scala 630:39]
  wire  _GEN_8861 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8624; // @[lut_35.scala 601:73 lut_35.scala 631:39]
  wire  _GEN_8862 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8625; // @[lut_35.scala 601:73 lut_35.scala 632:39]
  wire  _GEN_8863 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8626; // @[lut_35.scala 601:73 lut_35.scala 633:39]
  wire  _GEN_8864 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8627; // @[lut_35.scala 601:73 lut_35.scala 634:39]
  wire  _GEN_8865 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8628; // @[lut_35.scala 601:73 lut_35.scala 635:39]
  wire  _GEN_8866 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8629; // @[lut_35.scala 601:73 lut_35.scala 636:39]
  wire  _GEN_8867 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid | _GEN_8630; // @[lut_35.scala 601:73 lut_35.scala 637:34]
  wire  _GEN_8871 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 601:73 lut_35.scala 216:26 lut_35.scala 639:27]
  wire  _GEN_8874 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8634; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_8877 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8637; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_8880 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8640; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_8883 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8643; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_8886 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8646; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_8889 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8649; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_8892 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8652; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_8895 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8655; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_8898 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8658; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_8901 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8661; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_8904 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8664; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_8907 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8667; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_8910 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8670; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_8913 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8673; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_8916 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8676; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_8919 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8679; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_8922 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8682; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_8925 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8685; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_8928 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8688; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_8931 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8691; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_8934 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8694; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_8937 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8697; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_8940 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8700; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_8943 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8703; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_8946 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8706; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_8949 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8709; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_8952 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8712; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_8955 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8715; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_8958 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8718; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_8961 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8721; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_8964 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8724; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_8967 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8727; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire [5:0] _GEN_8968 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? push_mem_temp : _GEN_8728; // @[lut_35.scala 601:73 lut_35.scala 521:39]
  wire [31:0] _GEN_8969 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? push_id_temp : _GEN_8729; // @[lut_35.scala 601:73 lut_35.scala 522:39]
  wire  _GEN_8972 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8732; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_8975 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8735; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_8978 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8738; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_8981 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8741; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_8984 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8744; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_8987 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8747; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_8990 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8750; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_8993 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8753; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_8996 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8756; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_8999 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8759; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_9002 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8762; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_9005 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8765; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_9008 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8768; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_9011 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8771; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_9014 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8774; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_9017 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8777; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_9020 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8780; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_9023 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8783; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_9026 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8786; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_9029 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8789; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_9032 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8792; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_9035 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8795; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_9038 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8798; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_9041 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8801; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_9044 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8804; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_9047 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8807; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_9050 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8810; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_9053 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8813; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_9056 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8816; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_9059 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8819; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_9062 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8822; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_9065 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8825; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_9068 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8828; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_9071 = LUT_mem_MPORT_37_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8831; // @[lut_35.scala 601:73 lut_35.scala 216:26]
  wire  _GEN_9072 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8832; // @[lut_35.scala 563:74 lut_35.scala 564:38]
  wire  _GEN_9073 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid | _GEN_8833; // @[lut_35.scala 563:74 lut_35.scala 565:38]
  wire  _GEN_9074 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8834; // @[lut_35.scala 563:74 lut_35.scala 566:38]
  wire  _GEN_9075 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8835; // @[lut_35.scala 563:74 lut_35.scala 567:38]
  wire  _GEN_9076 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8836; // @[lut_35.scala 563:74 lut_35.scala 568:38]
  wire  _GEN_9077 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8837; // @[lut_35.scala 563:74 lut_35.scala 569:38]
  wire  _GEN_9078 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8838; // @[lut_35.scala 563:74 lut_35.scala 570:38]
  wire  _GEN_9079 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8839; // @[lut_35.scala 563:74 lut_35.scala 571:38]
  wire  _GEN_9080 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8840; // @[lut_35.scala 563:74 lut_35.scala 572:38]
  wire  _GEN_9081 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8841; // @[lut_35.scala 563:74 lut_35.scala 573:38]
  wire  _GEN_9082 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8842; // @[lut_35.scala 563:74 lut_35.scala 574:39]
  wire  _GEN_9083 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8843; // @[lut_35.scala 563:74 lut_35.scala 575:39]
  wire  _GEN_9084 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8844; // @[lut_35.scala 563:74 lut_35.scala 576:39]
  wire  _GEN_9085 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8845; // @[lut_35.scala 563:74 lut_35.scala 577:39]
  wire  _GEN_9086 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8846; // @[lut_35.scala 563:74 lut_35.scala 578:39]
  wire  _GEN_9087 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8847; // @[lut_35.scala 563:74 lut_35.scala 579:39]
  wire  _GEN_9088 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8848; // @[lut_35.scala 563:74 lut_35.scala 580:39]
  wire  _GEN_9089 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8849; // @[lut_35.scala 563:74 lut_35.scala 581:39]
  wire  _GEN_9090 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8850; // @[lut_35.scala 563:74 lut_35.scala 582:39]
  wire  _GEN_9091 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8851; // @[lut_35.scala 563:74 lut_35.scala 583:39]
  wire  _GEN_9092 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8852; // @[lut_35.scala 563:74 lut_35.scala 584:39]
  wire  _GEN_9093 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8853; // @[lut_35.scala 563:74 lut_35.scala 585:39]
  wire  _GEN_9094 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8854; // @[lut_35.scala 563:74 lut_35.scala 586:39]
  wire  _GEN_9095 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8855; // @[lut_35.scala 563:74 lut_35.scala 587:39]
  wire  _GEN_9096 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8856; // @[lut_35.scala 563:74 lut_35.scala 588:39]
  wire  _GEN_9097 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8857; // @[lut_35.scala 563:74 lut_35.scala 589:39]
  wire  _GEN_9098 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8858; // @[lut_35.scala 563:74 lut_35.scala 590:39]
  wire  _GEN_9099 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8859; // @[lut_35.scala 563:74 lut_35.scala 591:39]
  wire  _GEN_9100 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8860; // @[lut_35.scala 563:74 lut_35.scala 592:39]
  wire  _GEN_9101 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8861; // @[lut_35.scala 563:74 lut_35.scala 593:39]
  wire  _GEN_9102 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8862; // @[lut_35.scala 563:74 lut_35.scala 594:39]
  wire  _GEN_9103 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8863; // @[lut_35.scala 563:74 lut_35.scala 595:39]
  wire  _GEN_9104 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8864; // @[lut_35.scala 563:74 lut_35.scala 596:39]
  wire  _GEN_9105 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8865; // @[lut_35.scala 563:74 lut_35.scala 597:39]
  wire  _GEN_9106 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8866; // @[lut_35.scala 563:74 lut_35.scala 598:39]
  wire  _GEN_9107 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid | _GEN_8867; // @[lut_35.scala 563:74 lut_35.scala 599:34]
  wire  _GEN_9111 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 563:74 lut_35.scala 216:26 lut_35.scala 601:27]
  wire  _GEN_9114 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8871; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9117 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8874; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9120 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8877; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9123 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8880; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9126 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8883; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9129 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8886; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9132 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8889; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9135 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8892; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9138 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8895; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9141 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8898; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9144 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8901; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9147 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8904; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9150 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8907; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9153 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8910; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9156 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8913; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9159 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8916; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9162 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8919; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9165 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8922; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9168 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8925; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9171 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8928; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9174 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8931; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9177 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8934; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9180 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8937; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9183 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8940; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9186 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8943; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9189 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8946; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9192 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8949; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9195 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8952; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9198 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8955; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9201 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8958; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9204 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8961; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9207 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8964; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9210 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8967; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9215 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8972; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9218 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8975; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9221 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8978; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9224 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8981; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9227 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8984; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9230 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8987; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9233 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8990; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9236 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8993; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9239 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8996; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9242 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8999; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9245 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9002; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9248 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9005; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9251 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9008; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9254 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9011; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9257 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9014; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9260 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9017; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9263 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9020; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9266 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9023; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9269 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9026; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9272 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9029; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9275 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9032; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9278 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9035; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9281 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9038; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9284 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9041; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9287 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9044; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9290 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9047; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9293 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9050; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9296 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9053; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9299 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9056; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9302 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9059; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9305 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9062; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9308 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9065; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9311 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9068; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9314 = LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9071; // @[lut_35.scala 563:74 lut_35.scala 216:26]
  wire  _GEN_9315 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid | _GEN_9072; // @[lut_35.scala 525:68 lut_35.scala 526:38]
  wire  _GEN_9316 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9073; // @[lut_35.scala 525:68 lut_35.scala 527:38]
  wire  _GEN_9317 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9074; // @[lut_35.scala 525:68 lut_35.scala 528:38]
  wire  _GEN_9318 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9075; // @[lut_35.scala 525:68 lut_35.scala 529:38]
  wire  _GEN_9319 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9076; // @[lut_35.scala 525:68 lut_35.scala 530:38]
  wire  _GEN_9320 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9077; // @[lut_35.scala 525:68 lut_35.scala 531:38]
  wire  _GEN_9321 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9078; // @[lut_35.scala 525:68 lut_35.scala 532:38]
  wire  _GEN_9322 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9079; // @[lut_35.scala 525:68 lut_35.scala 533:38]
  wire  _GEN_9323 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9080; // @[lut_35.scala 525:68 lut_35.scala 534:38]
  wire  _GEN_9324 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9081; // @[lut_35.scala 525:68 lut_35.scala 535:38]
  wire  _GEN_9325 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9082; // @[lut_35.scala 525:68 lut_35.scala 536:39]
  wire  _GEN_9326 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9083; // @[lut_35.scala 525:68 lut_35.scala 537:39]
  wire  _GEN_9327 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9084; // @[lut_35.scala 525:68 lut_35.scala 538:39]
  wire  _GEN_9328 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9085; // @[lut_35.scala 525:68 lut_35.scala 539:39]
  wire  _GEN_9329 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9086; // @[lut_35.scala 525:68 lut_35.scala 540:39]
  wire  _GEN_9330 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9087; // @[lut_35.scala 525:68 lut_35.scala 541:39]
  wire  _GEN_9331 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9088; // @[lut_35.scala 525:68 lut_35.scala 542:39]
  wire  _GEN_9332 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9089; // @[lut_35.scala 525:68 lut_35.scala 543:39]
  wire  _GEN_9333 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9090; // @[lut_35.scala 525:68 lut_35.scala 544:39]
  wire  _GEN_9334 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9091; // @[lut_35.scala 525:68 lut_35.scala 545:39]
  wire  _GEN_9335 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9092; // @[lut_35.scala 525:68 lut_35.scala 546:39]
  wire  _GEN_9336 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9093; // @[lut_35.scala 525:68 lut_35.scala 547:39]
  wire  _GEN_9337 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9094; // @[lut_35.scala 525:68 lut_35.scala 548:39]
  wire  _GEN_9338 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9095; // @[lut_35.scala 525:68 lut_35.scala 549:39]
  wire  _GEN_9339 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9096; // @[lut_35.scala 525:68 lut_35.scala 550:39]
  wire  _GEN_9340 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9097; // @[lut_35.scala 525:68 lut_35.scala 551:39]
  wire  _GEN_9341 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9098; // @[lut_35.scala 525:68 lut_35.scala 552:39]
  wire  _GEN_9342 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9099; // @[lut_35.scala 525:68 lut_35.scala 553:39]
  wire  _GEN_9343 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9100; // @[lut_35.scala 525:68 lut_35.scala 554:39]
  wire  _GEN_9344 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9101; // @[lut_35.scala 525:68 lut_35.scala 555:39]
  wire  _GEN_9345 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9102; // @[lut_35.scala 525:68 lut_35.scala 556:39]
  wire  _GEN_9346 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9103; // @[lut_35.scala 525:68 lut_35.scala 557:39]
  wire  _GEN_9347 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9104; // @[lut_35.scala 525:68 lut_35.scala 558:39]
  wire  _GEN_9348 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9105; // @[lut_35.scala 525:68 lut_35.scala 559:39]
  wire  _GEN_9349 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9106; // @[lut_35.scala 525:68 lut_35.scala 560:39]
  wire  _GEN_9350 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid | _GEN_9107; // @[lut_35.scala 525:68 lut_35.scala 561:34]
  wire  _GEN_9354 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 525:68 lut_35.scala 216:26 lut_35.scala 563:27]
  wire  _GEN_9357 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9111; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9360 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9114; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9363 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9117; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9366 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9120; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9369 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9123; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9372 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9126; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9375 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9129; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9378 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9132; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9381 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9135; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9384 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9138; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9387 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9141; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9390 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9144; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9393 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9147; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9396 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9150; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9399 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9153; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9402 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9156; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9405 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9159; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9408 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9162; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9411 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9165; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9414 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9168; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9417 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9171; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9420 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9174; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9423 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9177; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9426 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9180; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9429 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9183; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9432 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9186; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9435 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9189; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9438 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9192; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9441 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9195; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9444 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9198; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9447 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9201; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9450 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9204; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9453 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9207; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9456 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9210; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9461 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9215; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9464 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9218; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9467 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9221; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9470 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9224; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9473 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9227; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9476 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9230; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9479 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9233; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9482 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9236; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9485 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9239; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9488 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9242; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9491 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9245; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9494 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9248; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9497 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9251; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9500 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9254; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9503 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9257; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9506 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9260; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9509 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9263; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9512 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9266; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9515 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9269; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9518 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9272; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9521 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9275; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9524 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9278; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9527 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9281; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9530 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9284; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9533 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9287; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9536 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9290; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9539 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9293; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9542 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9296; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9545 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9299; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9548 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9302; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9551 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9305; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9554 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9308; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9557 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9311; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9560 = LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9314; // @[lut_35.scala 525:68 lut_35.scala 216:26]
  wire  _GEN_9564 = push_1 & push_valid & _GEN_9315; // @[lut_35.scala 524:46 lut_35.scala 3415:32]
  wire  _GEN_9565 = push_1 & push_valid & _GEN_9316; // @[lut_35.scala 524:46 lut_35.scala 3416:32]
  wire  _GEN_9566 = push_1 & push_valid & _GEN_9317; // @[lut_35.scala 524:46 lut_35.scala 3417:32]
  wire  _GEN_9567 = push_1 & push_valid & _GEN_9318; // @[lut_35.scala 524:46 lut_35.scala 3418:32]
  wire  _GEN_9568 = push_1 & push_valid & _GEN_9319; // @[lut_35.scala 524:46 lut_35.scala 3419:32]
  wire  _GEN_9569 = push_1 & push_valid & _GEN_9320; // @[lut_35.scala 524:46 lut_35.scala 3420:32]
  wire  _GEN_9570 = push_1 & push_valid & _GEN_9321; // @[lut_35.scala 524:46 lut_35.scala 3421:32]
  wire  _GEN_9571 = push_1 & push_valid & _GEN_9322; // @[lut_35.scala 524:46 lut_35.scala 3422:32]
  wire  _GEN_9572 = push_1 & push_valid & _GEN_9323; // @[lut_35.scala 524:46 lut_35.scala 3423:42]
  wire  _GEN_9573 = push_1 & push_valid & _GEN_9324; // @[lut_35.scala 524:46 lut_35.scala 3424:42]
  wire  _GEN_9574 = push_1 & push_valid & _GEN_9325; // @[lut_35.scala 524:46 lut_35.scala 3425:43]
  wire  _GEN_9575 = push_1 & push_valid & _GEN_9326; // @[lut_35.scala 524:46 lut_35.scala 3426:43]
  wire  _GEN_9576 = push_1 & push_valid & _GEN_9327; // @[lut_35.scala 524:46 lut_35.scala 3427:43]
  wire  _GEN_9577 = push_1 & push_valid & _GEN_9328; // @[lut_35.scala 524:46 lut_35.scala 3428:43]
  wire  _GEN_9578 = push_1 & push_valid & _GEN_9329; // @[lut_35.scala 524:46 lut_35.scala 3429:43]
  wire  _GEN_9579 = push_1 & push_valid & _GEN_9330; // @[lut_35.scala 524:46 lut_35.scala 3430:43]
  wire  _GEN_9580 = push_1 & push_valid & _GEN_9331; // @[lut_35.scala 524:46 lut_35.scala 3431:43]
  wire  _GEN_9581 = push_1 & push_valid & _GEN_9332; // @[lut_35.scala 524:46 lut_35.scala 3432:43]
  wire  _GEN_9582 = push_1 & push_valid & _GEN_9333; // @[lut_35.scala 524:46 lut_35.scala 3433:43]
  wire  _GEN_9583 = push_1 & push_valid & _GEN_9334; // @[lut_35.scala 524:46 lut_35.scala 3434:43]
  wire  _GEN_9584 = push_1 & push_valid & _GEN_9335; // @[lut_35.scala 524:46 lut_35.scala 3435:43]
  wire  _GEN_9585 = push_1 & push_valid & _GEN_9336; // @[lut_35.scala 524:46 lut_35.scala 3436:43]
  wire  _GEN_9586 = push_1 & push_valid & _GEN_9337; // @[lut_35.scala 524:46 lut_35.scala 3437:43]
  wire  _GEN_9587 = push_1 & push_valid & _GEN_9338; // @[lut_35.scala 524:46 lut_35.scala 3438:43]
  wire  _GEN_9588 = push_1 & push_valid & _GEN_9339; // @[lut_35.scala 524:46 lut_35.scala 3439:43]
  wire  _GEN_9589 = push_1 & push_valid & _GEN_9340; // @[lut_35.scala 524:46 lut_35.scala 3440:43]
  wire  _GEN_9590 = push_1 & push_valid & _GEN_9341; // @[lut_35.scala 524:46 lut_35.scala 3441:43]
  wire  _GEN_9591 = push_1 & push_valid & _GEN_9342; // @[lut_35.scala 524:46 lut_35.scala 3442:43]
  wire  _GEN_9592 = push_1 & push_valid & _GEN_9343; // @[lut_35.scala 524:46 lut_35.scala 3443:43]
  wire  _GEN_9593 = push_1 & push_valid & _GEN_9344; // @[lut_35.scala 524:46 lut_35.scala 3444:43]
  wire  _GEN_9594 = push_1 & push_valid & _GEN_9345; // @[lut_35.scala 524:46 lut_35.scala 3445:43]
  wire  _GEN_9595 = push_1 & push_valid & _GEN_9346; // @[lut_35.scala 524:46 lut_35.scala 3446:43]
  wire  _GEN_9596 = push_1 & push_valid & _GEN_9347; // @[lut_35.scala 524:46 lut_35.scala 3447:43]
  wire  _GEN_9597 = push_1 & push_valid & _GEN_9348; // @[lut_35.scala 524:46 lut_35.scala 3448:43]
  wire  _GEN_9598 = push_1 & push_valid & _GEN_9349; // @[lut_35.scala 524:46 lut_35.scala 3449:43]
  wire  _GEN_9599 = push_1 & push_valid & _GEN_9350; // @[lut_35.scala 524:46 lut_35.scala 3450:30]
  reg  pop_1; // @[lut_35.scala 3494:50]
  reg [31:0] read_stack0_pop; // @[lut_35.scala 3495:38]
  reg [31:0] read_stack1_pop; // @[lut_35.scala 3496:38]
  reg [31:0] read_stack2_pop; // @[lut_35.scala 3497:38]
  reg [31:0] read_stack3_pop; // @[lut_35.scala 3498:38]
  reg [31:0] read_stack4_pop; // @[lut_35.scala 3499:38]
  reg [31:0] read_stack5_pop; // @[lut_35.scala 3500:38]
  reg [31:0] read_stack6_pop; // @[lut_35.scala 3501:38]
  reg [31:0] read_stack7_pop; // @[lut_35.scala 3502:38]
  reg [31:0] read_stack8_pop; // @[lut_35.scala 3503:38]
  reg [31:0] read_stack9_pop; // @[lut_35.scala 3504:38]
  reg [31:0] read_stack10_pop; // @[lut_35.scala 3505:39]
  reg [31:0] read_stack11_pop; // @[lut_35.scala 3506:39]
  reg [31:0] read_stack12_pop; // @[lut_35.scala 3507:39]
  reg [31:0] read_stack13_pop; // @[lut_35.scala 3508:39]
  reg [31:0] read_stack14_pop; // @[lut_35.scala 3509:39]
  reg [31:0] read_stack15_pop; // @[lut_35.scala 3510:39]
  reg [31:0] read_stack16_pop; // @[lut_35.scala 3511:39]
  reg [31:0] read_stack17_pop; // @[lut_35.scala 3512:39]
  reg [31:0] read_stack18_pop; // @[lut_35.scala 3513:39]
  reg [31:0] read_stack19_pop; // @[lut_35.scala 3514:39]
  reg [31:0] read_stack20_pop; // @[lut_35.scala 3515:39]
  reg [31:0] read_stack21_pop; // @[lut_35.scala 3516:39]
  reg [31:0] read_stack22_pop; // @[lut_35.scala 3517:39]
  reg [31:0] read_stack23_pop; // @[lut_35.scala 3518:39]
  reg [31:0] read_stack24_pop; // @[lut_35.scala 3519:39]
  reg [31:0] read_stack25_pop; // @[lut_35.scala 3520:39]
  reg [31:0] read_stack26_pop; // @[lut_35.scala 3521:39]
  reg [31:0] read_stack27_pop; // @[lut_35.scala 3522:39]
  reg [31:0] read_stack28_pop; // @[lut_35.scala 3523:39]
  reg [31:0] read_stack29_pop; // @[lut_35.scala 3524:39]
  reg [31:0] read_stack30_pop; // @[lut_35.scala 3525:39]
  reg [31:0] read_stack31_pop; // @[lut_35.scala 3526:39]
  reg [31:0] read_stack32_pop; // @[lut_35.scala 3527:39]
  reg [31:0] read_stack33_pop; // @[lut_35.scala 3528:39]
  reg [31:0] read_stack34_pop; // @[lut_35.scala 3529:39]
  reg [31:0] pop_ray_id; // @[lut_35.scala 3532:37]
  reg [31:0] pop_hitT_1; // @[lut_35.scala 3533:37]
  reg  pop_valid; // @[lut_35.scala 3534:36]
  reg  pop_0_1; // @[lut_35.scala 3537:46]
  reg  pop_1_1; // @[lut_35.scala 3538:46]
  reg  pop_2_1; // @[lut_35.scala 3539:46]
  reg  pop_3_1; // @[lut_35.scala 3540:46]
  reg  pop_4_1; // @[lut_35.scala 3541:46]
  reg  pop_5_1; // @[lut_35.scala 3542:46]
  reg  pop_6_1; // @[lut_35.scala 3543:46]
  reg  pop_7_1; // @[lut_35.scala 3544:46]
  reg  pop_8_1; // @[lut_35.scala 3545:46]
  reg  pop_9_1; // @[lut_35.scala 3546:46]
  reg  pop_10_1; // @[lut_35.scala 3547:47]
  reg  pop_11_1; // @[lut_35.scala 3548:47]
  reg  pop_12_1; // @[lut_35.scala 3549:47]
  reg  pop_13_1; // @[lut_35.scala 3550:47]
  reg  pop_14_1; // @[lut_35.scala 3551:47]
  reg  pop_15_1; // @[lut_35.scala 3552:47]
  reg  pop_16_1; // @[lut_35.scala 3553:47]
  reg  pop_17_1; // @[lut_35.scala 3554:47]
  reg  pop_18_1; // @[lut_35.scala 3555:47]
  reg  pop_19_1; // @[lut_35.scala 3556:47]
  reg  pop_20_1; // @[lut_35.scala 3557:47]
  reg  pop_21_1; // @[lut_35.scala 3558:47]
  reg  pop_22_1; // @[lut_35.scala 3559:47]
  reg  pop_23_1; // @[lut_35.scala 3560:47]
  reg  pop_24_1; // @[lut_35.scala 3561:47]
  reg  pop_25_1; // @[lut_35.scala 3562:47]
  reg  pop_26_1; // @[lut_35.scala 3563:47]
  reg  pop_27_1; // @[lut_35.scala 3564:47]
  reg  pop_28_1; // @[lut_35.scala 3565:47]
  reg  pop_29_1; // @[lut_35.scala 3566:47]
  reg  pop_30_1; // @[lut_35.scala 3567:47]
  reg  pop_31_1; // @[lut_35.scala 3568:47]
  reg  pop_32_1; // @[lut_35.scala 3569:47]
  reg  pop_33_1; // @[lut_35.scala 3570:47]
  reg  pop_34_1; // @[lut_35.scala 3571:47]
  reg  pop_valid_2; // @[lut_35.scala 3573:47]
  reg [31:0] pop_ray_id_2; // @[lut_35.scala 3575:47]
  reg [31:0] pop_hitT_2; // @[lut_35.scala 3576:47]
  reg  no_match; // @[lut_35.scala 3578:47]
  wire  _T_567 = io_pop & io_pop_valid; // @[lut_35.scala 3619:28]
  wire  _T_576 = pop_1 & pop_ray_id != read_stack0_pop & pop_ray_id != read_stack1_pop & pop_ray_id != read_stack2_pop
     & pop_ray_id != read_stack3_pop; // @[lut_35.scala 3631:124]
  wire  _T_584 = _T_576 & pop_ray_id != read_stack4_pop & pop_ray_id != read_stack5_pop & pop_ray_id != read_stack6_pop
     & pop_ray_id != read_stack7_pop; // @[lut_35.scala 3632:108]
  wire  _T_592 = _T_584 & pop_ray_id != read_stack8_pop & pop_ray_id != read_stack9_pop & pop_ray_id != read_stack10_pop
     & pop_ray_id != read_stack11_pop; // @[lut_35.scala 3633:109]
  wire  _T_600 = _T_592 & pop_ray_id != read_stack12_pop & pop_ray_id != read_stack13_pop & pop_ray_id !=
    read_stack14_pop & pop_ray_id != read_stack15_pop; // @[lut_35.scala 3634:111]
  wire  _T_608 = _T_600 & pop_ray_id != read_stack16_pop & pop_ray_id != read_stack17_pop & pop_ray_id !=
    read_stack18_pop & pop_ray_id != read_stack19_pop; // @[lut_35.scala 3635:111]
  wire  _T_616 = _T_608 & pop_ray_id != read_stack20_pop & pop_ray_id != read_stack21_pop & pop_ray_id !=
    read_stack22_pop & pop_ray_id != read_stack23_pop; // @[lut_35.scala 3636:111]
  wire  _T_624 = _T_616 & pop_ray_id != read_stack24_pop & pop_ray_id != read_stack25_pop & pop_ray_id !=
    read_stack26_pop & pop_ray_id != read_stack27_pop; // @[lut_35.scala 3637:111]
  wire  _T_631 = pop_ray_id != read_stack31_pop; // @[lut_35.scala 3638:125]
  wire  _T_632 = _T_624 & pop_ray_id != read_stack28_pop & pop_ray_id != read_stack29_pop & pop_ray_id !=
    read_stack30_pop & pop_ray_id != read_stack31_pop; // @[lut_35.scala 3638:111]
  wire  _T_640 = _T_632 & _T_631 & pop_ray_id != read_stack32_pop & pop_ray_id != read_stack33_pop & pop_ray_id !=
    read_stack34_pop; // @[lut_35.scala 3639:111]
  reg  no_match_1; // @[lut_35.scala 3644:51]
  reg  no_match_2; // @[lut_35.scala 3645:51]
  wire  _T_646 = read_stack0_pop == pop_ray_id & pop_valid; // @[lut_35.scala 3650:45]
  wire  _T_649 = read_stack1_pop == pop_ray_id & pop_valid; // @[lut_35.scala 3690:55]
  wire  _T_652 = read_stack2_pop == pop_ray_id & pop_valid; // @[lut_35.scala 3730:55]
  wire  _T_655 = read_stack3_pop == pop_ray_id & pop_valid; // @[lut_35.scala 3770:55]
  wire  _T_658 = read_stack4_pop == pop_ray_id & pop_valid; // @[lut_35.scala 3810:55]
  wire  _T_661 = read_stack5_pop == pop_ray_id & pop_valid; // @[lut_35.scala 3850:55]
  wire  _T_664 = read_stack6_pop == pop_ray_id & pop_valid; // @[lut_35.scala 3890:55]
  wire  _T_667 = read_stack7_pop == pop_ray_id & pop_valid; // @[lut_35.scala 3930:55]
  wire  _T_670 = read_stack8_pop == pop_ray_id & pop_valid; // @[lut_35.scala 3970:55]
  wire  _T_673 = read_stack9_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4011:55]
  wire  _T_676 = read_stack10_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4051:56]
  wire  _T_679 = read_stack11_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4091:56]
  wire  _T_682 = read_stack12_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4131:56]
  wire  _T_685 = read_stack13_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4171:56]
  wire  _T_688 = read_stack14_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4211:56]
  wire  _T_691 = read_stack15_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4251:56]
  wire  _T_694 = read_stack16_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4291:56]
  wire  _T_697 = read_stack17_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4331:56]
  wire  _T_700 = read_stack18_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4371:56]
  wire  _T_703 = read_stack19_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4411:56]
  wire  _T_706 = read_stack20_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4451:56]
  wire  _T_709 = read_stack21_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4491:56]
  wire  _T_712 = read_stack22_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4531:56]
  wire  _T_715 = read_stack23_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4571:56]
  wire  _T_718 = read_stack24_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4611:56]
  wire  _T_721 = read_stack25_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4651:56]
  wire  _T_724 = read_stack26_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4691:56]
  wire  _T_727 = read_stack27_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4731:56]
  wire  _T_730 = read_stack28_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4771:56]
  wire  _T_733 = read_stack29_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4811:56]
  wire  _T_736 = read_stack30_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4851:56]
  wire  _T_739 = read_stack31_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4891:56]
  wire  _T_742 = read_stack32_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4931:56]
  wire  _T_745 = read_stack33_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4971:56]
  wire  _T_748 = read_stack34_pop == pop_ray_id & pop_valid; // @[lut_35.scala 5011:56]
  wire [31:0] _GEN_9818 = read_stack34_pop == pop_ray_id & pop_valid ? pop_ray_id : pop_ray_id_2; // @[lut_35.scala 5011:78 lut_35.scala 5049:38 lut_35.scala 3575:47]
  wire [31:0] _GEN_9819 = read_stack34_pop == pop_ray_id & pop_valid ? pop_hitT_1 : pop_hitT_2; // @[lut_35.scala 5011:78 lut_35.scala 5050:41 lut_35.scala 3576:47]
  wire  _GEN_9822 = read_stack33_pop == pop_ray_id & pop_valid ? 1'h0 : _T_748; // @[lut_35.scala 4971:78 lut_35.scala 5006:45]
  wire  _GEN_9823 = read_stack33_pop == pop_ray_id & pop_valid | _T_748; // @[lut_35.scala 4971:78 lut_35.scala 5007:40]
  wire [31:0] _GEN_9825 = read_stack33_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_9818; // @[lut_35.scala 4971:78 lut_35.scala 5009:38]
  wire [31:0] _GEN_9826 = read_stack33_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_9819; // @[lut_35.scala 4971:78 lut_35.scala 5010:41]
  wire  _GEN_9829 = read_stack32_pop == pop_ray_id & pop_valid ? 1'h0 : _T_745; // @[lut_35.scala 4931:78 lut_35.scala 4965:45]
  wire  _GEN_9830 = read_stack32_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9822; // @[lut_35.scala 4931:78 lut_35.scala 4966:45]
  wire  _GEN_9831 = read_stack32_pop == pop_ray_id & pop_valid | _GEN_9823; // @[lut_35.scala 4931:78 lut_35.scala 4967:40]
  wire [31:0] _GEN_9833 = read_stack32_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_9825; // @[lut_35.scala 4931:78 lut_35.scala 4969:38]
  wire [31:0] _GEN_9834 = read_stack32_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_9826; // @[lut_35.scala 4931:78 lut_35.scala 4970:41]
  wire  _GEN_9837 = read_stack31_pop == pop_ray_id & pop_valid ? 1'h0 : _T_742; // @[lut_35.scala 4891:78 lut_35.scala 4924:45]
  wire  _GEN_9838 = read_stack31_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9829; // @[lut_35.scala 4891:78 lut_35.scala 4925:45]
  wire  _GEN_9839 = read_stack31_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9830; // @[lut_35.scala 4891:78 lut_35.scala 4926:45]
  wire  _GEN_9840 = read_stack31_pop == pop_ray_id & pop_valid | _GEN_9831; // @[lut_35.scala 4891:78 lut_35.scala 4927:40]
  wire [31:0] _GEN_9842 = read_stack31_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_9833; // @[lut_35.scala 4891:78 lut_35.scala 4929:38]
  wire [31:0] _GEN_9843 = read_stack31_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_9834; // @[lut_35.scala 4891:78 lut_35.scala 4930:41]
  wire  _GEN_9846 = read_stack30_pop == pop_ray_id & pop_valid ? 1'h0 : _T_739; // @[lut_35.scala 4851:78 lut_35.scala 4883:45]
  wire  _GEN_9847 = read_stack30_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9837; // @[lut_35.scala 4851:78 lut_35.scala 4884:45]
  wire  _GEN_9848 = read_stack30_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9838; // @[lut_35.scala 4851:78 lut_35.scala 4885:45]
  wire  _GEN_9849 = read_stack30_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9839; // @[lut_35.scala 4851:78 lut_35.scala 4886:45]
  wire  _GEN_9850 = read_stack30_pop == pop_ray_id & pop_valid | _GEN_9840; // @[lut_35.scala 4851:78 lut_35.scala 4887:40]
  wire [31:0] _GEN_9852 = read_stack30_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_9842; // @[lut_35.scala 4851:78 lut_35.scala 4889:38]
  wire [31:0] _GEN_9853 = read_stack30_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_9843; // @[lut_35.scala 4851:78 lut_35.scala 4890:41]
  wire  _GEN_9856 = read_stack29_pop == pop_ray_id & pop_valid ? 1'h0 : _T_736; // @[lut_35.scala 4811:78 lut_35.scala 4842:45]
  wire  _GEN_9857 = read_stack29_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9846; // @[lut_35.scala 4811:78 lut_35.scala 4843:45]
  wire  _GEN_9858 = read_stack29_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9847; // @[lut_35.scala 4811:78 lut_35.scala 4844:45]
  wire  _GEN_9859 = read_stack29_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9848; // @[lut_35.scala 4811:78 lut_35.scala 4845:45]
  wire  _GEN_9860 = read_stack29_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9849; // @[lut_35.scala 4811:78 lut_35.scala 4846:45]
  wire  _GEN_9861 = read_stack29_pop == pop_ray_id & pop_valid | _GEN_9850; // @[lut_35.scala 4811:78 lut_35.scala 4847:40]
  wire [31:0] _GEN_9863 = read_stack29_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_9852; // @[lut_35.scala 4811:78 lut_35.scala 4849:38]
  wire [31:0] _GEN_9864 = read_stack29_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_9853; // @[lut_35.scala 4811:78 lut_35.scala 4850:41]
  wire  _GEN_9867 = read_stack28_pop == pop_ray_id & pop_valid ? 1'h0 : _T_733; // @[lut_35.scala 4771:78 lut_35.scala 4801:45]
  wire  _GEN_9868 = read_stack28_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9856; // @[lut_35.scala 4771:78 lut_35.scala 4802:45]
  wire  _GEN_9869 = read_stack28_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9857; // @[lut_35.scala 4771:78 lut_35.scala 4803:45]
  wire  _GEN_9870 = read_stack28_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9858; // @[lut_35.scala 4771:78 lut_35.scala 4804:45]
  wire  _GEN_9871 = read_stack28_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9859; // @[lut_35.scala 4771:78 lut_35.scala 4805:45]
  wire  _GEN_9872 = read_stack28_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9860; // @[lut_35.scala 4771:78 lut_35.scala 4806:45]
  wire  _GEN_9873 = read_stack28_pop == pop_ray_id & pop_valid | _GEN_9861; // @[lut_35.scala 4771:78 lut_35.scala 4807:40]
  wire [31:0] _GEN_9875 = read_stack28_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_9863; // @[lut_35.scala 4771:78 lut_35.scala 4809:38]
  wire [31:0] _GEN_9876 = read_stack28_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_9864; // @[lut_35.scala 4771:78 lut_35.scala 4810:41]
  wire  _GEN_9879 = read_stack27_pop == pop_ray_id & pop_valid ? 1'h0 : _T_730; // @[lut_35.scala 4731:78 lut_35.scala 4760:45]
  wire  _GEN_9880 = read_stack27_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9867; // @[lut_35.scala 4731:78 lut_35.scala 4761:45]
  wire  _GEN_9881 = read_stack27_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9868; // @[lut_35.scala 4731:78 lut_35.scala 4762:45]
  wire  _GEN_9882 = read_stack27_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9869; // @[lut_35.scala 4731:78 lut_35.scala 4763:45]
  wire  _GEN_9883 = read_stack27_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9870; // @[lut_35.scala 4731:78 lut_35.scala 4764:45]
  wire  _GEN_9884 = read_stack27_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9871; // @[lut_35.scala 4731:78 lut_35.scala 4765:45]
  wire  _GEN_9885 = read_stack27_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9872; // @[lut_35.scala 4731:78 lut_35.scala 4766:45]
  wire  _GEN_9886 = read_stack27_pop == pop_ray_id & pop_valid | _GEN_9873; // @[lut_35.scala 4731:78 lut_35.scala 4767:40]
  wire [31:0] _GEN_9888 = read_stack27_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_9875; // @[lut_35.scala 4731:78 lut_35.scala 4769:38]
  wire [31:0] _GEN_9889 = read_stack27_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_9876; // @[lut_35.scala 4731:78 lut_35.scala 4770:41]
  wire  _GEN_9892 = read_stack26_pop == pop_ray_id & pop_valid ? 1'h0 : _T_727; // @[lut_35.scala 4691:78 lut_35.scala 4719:45]
  wire  _GEN_9893 = read_stack26_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9879; // @[lut_35.scala 4691:78 lut_35.scala 4720:45]
  wire  _GEN_9894 = read_stack26_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9880; // @[lut_35.scala 4691:78 lut_35.scala 4721:45]
  wire  _GEN_9895 = read_stack26_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9881; // @[lut_35.scala 4691:78 lut_35.scala 4722:45]
  wire  _GEN_9896 = read_stack26_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9882; // @[lut_35.scala 4691:78 lut_35.scala 4723:45]
  wire  _GEN_9897 = read_stack26_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9883; // @[lut_35.scala 4691:78 lut_35.scala 4724:45]
  wire  _GEN_9898 = read_stack26_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9884; // @[lut_35.scala 4691:78 lut_35.scala 4725:45]
  wire  _GEN_9899 = read_stack26_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9885; // @[lut_35.scala 4691:78 lut_35.scala 4726:45]
  wire  _GEN_9900 = read_stack26_pop == pop_ray_id & pop_valid | _GEN_9886; // @[lut_35.scala 4691:78 lut_35.scala 4727:40]
  wire [31:0] _GEN_9902 = read_stack26_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_9888; // @[lut_35.scala 4691:78 lut_35.scala 4729:38]
  wire [31:0] _GEN_9903 = read_stack26_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_9889; // @[lut_35.scala 4691:78 lut_35.scala 4730:41]
  wire  _GEN_9906 = read_stack25_pop == pop_ray_id & pop_valid ? 1'h0 : _T_724; // @[lut_35.scala 4651:78 lut_35.scala 4678:45]
  wire  _GEN_9907 = read_stack25_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9892; // @[lut_35.scala 4651:78 lut_35.scala 4679:45]
  wire  _GEN_9908 = read_stack25_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9893; // @[lut_35.scala 4651:78 lut_35.scala 4680:45]
  wire  _GEN_9909 = read_stack25_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9894; // @[lut_35.scala 4651:78 lut_35.scala 4681:45]
  wire  _GEN_9910 = read_stack25_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9895; // @[lut_35.scala 4651:78 lut_35.scala 4682:45]
  wire  _GEN_9911 = read_stack25_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9896; // @[lut_35.scala 4651:78 lut_35.scala 4683:45]
  wire  _GEN_9912 = read_stack25_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9897; // @[lut_35.scala 4651:78 lut_35.scala 4684:45]
  wire  _GEN_9913 = read_stack25_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9898; // @[lut_35.scala 4651:78 lut_35.scala 4685:45]
  wire  _GEN_9914 = read_stack25_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9899; // @[lut_35.scala 4651:78 lut_35.scala 4686:45]
  wire  _GEN_9915 = read_stack25_pop == pop_ray_id & pop_valid | _GEN_9900; // @[lut_35.scala 4651:78 lut_35.scala 4687:40]
  wire [31:0] _GEN_9917 = read_stack25_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_9902; // @[lut_35.scala 4651:78 lut_35.scala 4689:38]
  wire [31:0] _GEN_9918 = read_stack25_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_9903; // @[lut_35.scala 4651:78 lut_35.scala 4690:41]
  wire  _GEN_9921 = read_stack24_pop == pop_ray_id & pop_valid ? 1'h0 : _T_721; // @[lut_35.scala 4611:78 lut_35.scala 4637:45]
  wire  _GEN_9922 = read_stack24_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9906; // @[lut_35.scala 4611:78 lut_35.scala 4638:45]
  wire  _GEN_9923 = read_stack24_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9907; // @[lut_35.scala 4611:78 lut_35.scala 4639:45]
  wire  _GEN_9924 = read_stack24_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9908; // @[lut_35.scala 4611:78 lut_35.scala 4640:45]
  wire  _GEN_9925 = read_stack24_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9909; // @[lut_35.scala 4611:78 lut_35.scala 4641:45]
  wire  _GEN_9926 = read_stack24_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9910; // @[lut_35.scala 4611:78 lut_35.scala 4642:45]
  wire  _GEN_9927 = read_stack24_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9911; // @[lut_35.scala 4611:78 lut_35.scala 4643:45]
  wire  _GEN_9928 = read_stack24_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9912; // @[lut_35.scala 4611:78 lut_35.scala 4644:45]
  wire  _GEN_9929 = read_stack24_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9913; // @[lut_35.scala 4611:78 lut_35.scala 4645:45]
  wire  _GEN_9930 = read_stack24_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9914; // @[lut_35.scala 4611:78 lut_35.scala 4646:45]
  wire  _GEN_9931 = read_stack24_pop == pop_ray_id & pop_valid | _GEN_9915; // @[lut_35.scala 4611:78 lut_35.scala 4647:40]
  wire [31:0] _GEN_9933 = read_stack24_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_9917; // @[lut_35.scala 4611:78 lut_35.scala 4649:38]
  wire [31:0] _GEN_9934 = read_stack24_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_9918; // @[lut_35.scala 4611:78 lut_35.scala 4650:41]
  wire  _GEN_9937 = read_stack23_pop == pop_ray_id & pop_valid ? 1'h0 : _T_718; // @[lut_35.scala 4571:78 lut_35.scala 4596:45]
  wire  _GEN_9938 = read_stack23_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9921; // @[lut_35.scala 4571:78 lut_35.scala 4597:45]
  wire  _GEN_9939 = read_stack23_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9922; // @[lut_35.scala 4571:78 lut_35.scala 4598:45]
  wire  _GEN_9940 = read_stack23_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9923; // @[lut_35.scala 4571:78 lut_35.scala 4599:45]
  wire  _GEN_9941 = read_stack23_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9924; // @[lut_35.scala 4571:78 lut_35.scala 4600:45]
  wire  _GEN_9942 = read_stack23_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9925; // @[lut_35.scala 4571:78 lut_35.scala 4601:45]
  wire  _GEN_9943 = read_stack23_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9926; // @[lut_35.scala 4571:78 lut_35.scala 4602:45]
  wire  _GEN_9944 = read_stack23_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9927; // @[lut_35.scala 4571:78 lut_35.scala 4603:45]
  wire  _GEN_9945 = read_stack23_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9928; // @[lut_35.scala 4571:78 lut_35.scala 4604:45]
  wire  _GEN_9946 = read_stack23_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9929; // @[lut_35.scala 4571:78 lut_35.scala 4605:45]
  wire  _GEN_9947 = read_stack23_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9930; // @[lut_35.scala 4571:78 lut_35.scala 4606:45]
  wire  _GEN_9948 = read_stack23_pop == pop_ray_id & pop_valid | _GEN_9931; // @[lut_35.scala 4571:78 lut_35.scala 4607:40]
  wire [31:0] _GEN_9950 = read_stack23_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_9933; // @[lut_35.scala 4571:78 lut_35.scala 4609:38]
  wire [31:0] _GEN_9951 = read_stack23_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_9934; // @[lut_35.scala 4571:78 lut_35.scala 4610:41]
  wire  _GEN_9954 = read_stack22_pop == pop_ray_id & pop_valid ? 1'h0 : _T_715; // @[lut_35.scala 4531:78 lut_35.scala 4555:45]
  wire  _GEN_9955 = read_stack22_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9937; // @[lut_35.scala 4531:78 lut_35.scala 4556:45]
  wire  _GEN_9956 = read_stack22_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9938; // @[lut_35.scala 4531:78 lut_35.scala 4557:45]
  wire  _GEN_9957 = read_stack22_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9939; // @[lut_35.scala 4531:78 lut_35.scala 4558:45]
  wire  _GEN_9958 = read_stack22_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9940; // @[lut_35.scala 4531:78 lut_35.scala 4559:45]
  wire  _GEN_9959 = read_stack22_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9941; // @[lut_35.scala 4531:78 lut_35.scala 4560:45]
  wire  _GEN_9960 = read_stack22_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9942; // @[lut_35.scala 4531:78 lut_35.scala 4561:45]
  wire  _GEN_9961 = read_stack22_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9943; // @[lut_35.scala 4531:78 lut_35.scala 4562:45]
  wire  _GEN_9962 = read_stack22_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9944; // @[lut_35.scala 4531:78 lut_35.scala 4563:45]
  wire  _GEN_9963 = read_stack22_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9945; // @[lut_35.scala 4531:78 lut_35.scala 4564:45]
  wire  _GEN_9964 = read_stack22_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9946; // @[lut_35.scala 4531:78 lut_35.scala 4565:45]
  wire  _GEN_9965 = read_stack22_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9947; // @[lut_35.scala 4531:78 lut_35.scala 4566:45]
  wire  _GEN_9966 = read_stack22_pop == pop_ray_id & pop_valid | _GEN_9948; // @[lut_35.scala 4531:78 lut_35.scala 4567:40]
  wire [31:0] _GEN_9968 = read_stack22_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_9950; // @[lut_35.scala 4531:78 lut_35.scala 4569:38]
  wire [31:0] _GEN_9969 = read_stack22_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_9951; // @[lut_35.scala 4531:78 lut_35.scala 4570:41]
  wire  _GEN_9972 = read_stack21_pop == pop_ray_id & pop_valid ? 1'h0 : _T_712; // @[lut_35.scala 4491:78 lut_35.scala 4514:45]
  wire  _GEN_9973 = read_stack21_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9954; // @[lut_35.scala 4491:78 lut_35.scala 4515:45]
  wire  _GEN_9974 = read_stack21_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9955; // @[lut_35.scala 4491:78 lut_35.scala 4516:45]
  wire  _GEN_9975 = read_stack21_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9956; // @[lut_35.scala 4491:78 lut_35.scala 4517:45]
  wire  _GEN_9976 = read_stack21_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9957; // @[lut_35.scala 4491:78 lut_35.scala 4518:45]
  wire  _GEN_9977 = read_stack21_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9958; // @[lut_35.scala 4491:78 lut_35.scala 4519:45]
  wire  _GEN_9978 = read_stack21_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9959; // @[lut_35.scala 4491:78 lut_35.scala 4520:45]
  wire  _GEN_9979 = read_stack21_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9960; // @[lut_35.scala 4491:78 lut_35.scala 4521:45]
  wire  _GEN_9980 = read_stack21_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9961; // @[lut_35.scala 4491:78 lut_35.scala 4522:45]
  wire  _GEN_9981 = read_stack21_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9962; // @[lut_35.scala 4491:78 lut_35.scala 4523:45]
  wire  _GEN_9982 = read_stack21_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9963; // @[lut_35.scala 4491:78 lut_35.scala 4524:45]
  wire  _GEN_9983 = read_stack21_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9964; // @[lut_35.scala 4491:78 lut_35.scala 4525:45]
  wire  _GEN_9984 = read_stack21_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9965; // @[lut_35.scala 4491:78 lut_35.scala 4526:45]
  wire  _GEN_9985 = read_stack21_pop == pop_ray_id & pop_valid | _GEN_9966; // @[lut_35.scala 4491:78 lut_35.scala 4527:40]
  wire [31:0] _GEN_9987 = read_stack21_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_9968; // @[lut_35.scala 4491:78 lut_35.scala 4529:38]
  wire [31:0] _GEN_9988 = read_stack21_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_9969; // @[lut_35.scala 4491:78 lut_35.scala 4530:41]
  wire  _GEN_9991 = read_stack20_pop == pop_ray_id & pop_valid ? 1'h0 : _T_709; // @[lut_35.scala 4451:78 lut_35.scala 4473:45]
  wire  _GEN_9992 = read_stack20_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9972; // @[lut_35.scala 4451:78 lut_35.scala 4474:45]
  wire  _GEN_9993 = read_stack20_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9973; // @[lut_35.scala 4451:78 lut_35.scala 4475:45]
  wire  _GEN_9994 = read_stack20_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9974; // @[lut_35.scala 4451:78 lut_35.scala 4476:45]
  wire  _GEN_9995 = read_stack20_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9975; // @[lut_35.scala 4451:78 lut_35.scala 4477:45]
  wire  _GEN_9996 = read_stack20_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9976; // @[lut_35.scala 4451:78 lut_35.scala 4478:45]
  wire  _GEN_9997 = read_stack20_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9977; // @[lut_35.scala 4451:78 lut_35.scala 4479:45]
  wire  _GEN_9998 = read_stack20_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9978; // @[lut_35.scala 4451:78 lut_35.scala 4480:45]
  wire  _GEN_9999 = read_stack20_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9979; // @[lut_35.scala 4451:78 lut_35.scala 4481:45]
  wire  _GEN_10000 = read_stack20_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9980; // @[lut_35.scala 4451:78 lut_35.scala 4482:45]
  wire  _GEN_10001 = read_stack20_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9981; // @[lut_35.scala 4451:78 lut_35.scala 4483:45]
  wire  _GEN_10002 = read_stack20_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9982; // @[lut_35.scala 4451:78 lut_35.scala 4484:45]
  wire  _GEN_10003 = read_stack20_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9983; // @[lut_35.scala 4451:78 lut_35.scala 4485:45]
  wire  _GEN_10004 = read_stack20_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9984; // @[lut_35.scala 4451:78 lut_35.scala 4486:45]
  wire  _GEN_10005 = read_stack20_pop == pop_ray_id & pop_valid | _GEN_9985; // @[lut_35.scala 4451:78 lut_35.scala 4487:40]
  wire [31:0] _GEN_10007 = read_stack20_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_9987; // @[lut_35.scala 4451:78 lut_35.scala 4489:38]
  wire [31:0] _GEN_10008 = read_stack20_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_9988; // @[lut_35.scala 4451:78 lut_35.scala 4490:41]
  wire  _GEN_10011 = read_stack19_pop == pop_ray_id & pop_valid ? 1'h0 : _T_706; // @[lut_35.scala 4411:78 lut_35.scala 4432:45]
  wire  _GEN_10012 = read_stack19_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9991; // @[lut_35.scala 4411:78 lut_35.scala 4433:45]
  wire  _GEN_10013 = read_stack19_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9992; // @[lut_35.scala 4411:78 lut_35.scala 4434:45]
  wire  _GEN_10014 = read_stack19_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9993; // @[lut_35.scala 4411:78 lut_35.scala 4435:45]
  wire  _GEN_10015 = read_stack19_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9994; // @[lut_35.scala 4411:78 lut_35.scala 4436:45]
  wire  _GEN_10016 = read_stack19_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9995; // @[lut_35.scala 4411:78 lut_35.scala 4437:45]
  wire  _GEN_10017 = read_stack19_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9996; // @[lut_35.scala 4411:78 lut_35.scala 4438:45]
  wire  _GEN_10018 = read_stack19_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9997; // @[lut_35.scala 4411:78 lut_35.scala 4439:45]
  wire  _GEN_10019 = read_stack19_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9998; // @[lut_35.scala 4411:78 lut_35.scala 4440:45]
  wire  _GEN_10020 = read_stack19_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_9999; // @[lut_35.scala 4411:78 lut_35.scala 4441:45]
  wire  _GEN_10021 = read_stack19_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10000; // @[lut_35.scala 4411:78 lut_35.scala 4442:45]
  wire  _GEN_10022 = read_stack19_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10001; // @[lut_35.scala 4411:78 lut_35.scala 4443:45]
  wire  _GEN_10023 = read_stack19_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10002; // @[lut_35.scala 4411:78 lut_35.scala 4444:45]
  wire  _GEN_10024 = read_stack19_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10003; // @[lut_35.scala 4411:78 lut_35.scala 4445:45]
  wire  _GEN_10025 = read_stack19_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10004; // @[lut_35.scala 4411:78 lut_35.scala 4446:45]
  wire  _GEN_10026 = read_stack19_pop == pop_ray_id & pop_valid | _GEN_10005; // @[lut_35.scala 4411:78 lut_35.scala 4447:40]
  wire [31:0] _GEN_10028 = read_stack19_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_10007; // @[lut_35.scala 4411:78 lut_35.scala 4449:38]
  wire [31:0] _GEN_10029 = read_stack19_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_10008; // @[lut_35.scala 4411:78 lut_35.scala 4450:41]
  wire  _GEN_10032 = read_stack18_pop == pop_ray_id & pop_valid ? 1'h0 : _T_703; // @[lut_35.scala 4371:78 lut_35.scala 4391:45]
  wire  _GEN_10033 = read_stack18_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10011; // @[lut_35.scala 4371:78 lut_35.scala 4392:45]
  wire  _GEN_10034 = read_stack18_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10012; // @[lut_35.scala 4371:78 lut_35.scala 4393:45]
  wire  _GEN_10035 = read_stack18_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10013; // @[lut_35.scala 4371:78 lut_35.scala 4394:45]
  wire  _GEN_10036 = read_stack18_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10014; // @[lut_35.scala 4371:78 lut_35.scala 4395:45]
  wire  _GEN_10037 = read_stack18_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10015; // @[lut_35.scala 4371:78 lut_35.scala 4396:45]
  wire  _GEN_10038 = read_stack18_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10016; // @[lut_35.scala 4371:78 lut_35.scala 4397:45]
  wire  _GEN_10039 = read_stack18_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10017; // @[lut_35.scala 4371:78 lut_35.scala 4398:45]
  wire  _GEN_10040 = read_stack18_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10018; // @[lut_35.scala 4371:78 lut_35.scala 4399:45]
  wire  _GEN_10041 = read_stack18_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10019; // @[lut_35.scala 4371:78 lut_35.scala 4400:45]
  wire  _GEN_10042 = read_stack18_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10020; // @[lut_35.scala 4371:78 lut_35.scala 4401:45]
  wire  _GEN_10043 = read_stack18_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10021; // @[lut_35.scala 4371:78 lut_35.scala 4402:45]
  wire  _GEN_10044 = read_stack18_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10022; // @[lut_35.scala 4371:78 lut_35.scala 4403:45]
  wire  _GEN_10045 = read_stack18_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10023; // @[lut_35.scala 4371:78 lut_35.scala 4404:45]
  wire  _GEN_10046 = read_stack18_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10024; // @[lut_35.scala 4371:78 lut_35.scala 4405:45]
  wire  _GEN_10047 = read_stack18_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10025; // @[lut_35.scala 4371:78 lut_35.scala 4406:45]
  wire  _GEN_10048 = read_stack18_pop == pop_ray_id & pop_valid | _GEN_10026; // @[lut_35.scala 4371:78 lut_35.scala 4407:40]
  wire [31:0] _GEN_10050 = read_stack18_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_10028; // @[lut_35.scala 4371:78 lut_35.scala 4409:38]
  wire [31:0] _GEN_10051 = read_stack18_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_10029; // @[lut_35.scala 4371:78 lut_35.scala 4410:41]
  wire  _GEN_10054 = read_stack17_pop == pop_ray_id & pop_valid ? 1'h0 : _T_700; // @[lut_35.scala 4331:78 lut_35.scala 4350:45]
  wire  _GEN_10055 = read_stack17_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10032; // @[lut_35.scala 4331:78 lut_35.scala 4351:45]
  wire  _GEN_10056 = read_stack17_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10033; // @[lut_35.scala 4331:78 lut_35.scala 4352:45]
  wire  _GEN_10057 = read_stack17_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10034; // @[lut_35.scala 4331:78 lut_35.scala 4353:45]
  wire  _GEN_10058 = read_stack17_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10035; // @[lut_35.scala 4331:78 lut_35.scala 4354:45]
  wire  _GEN_10059 = read_stack17_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10036; // @[lut_35.scala 4331:78 lut_35.scala 4355:45]
  wire  _GEN_10060 = read_stack17_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10037; // @[lut_35.scala 4331:78 lut_35.scala 4356:45]
  wire  _GEN_10061 = read_stack17_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10038; // @[lut_35.scala 4331:78 lut_35.scala 4357:45]
  wire  _GEN_10062 = read_stack17_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10039; // @[lut_35.scala 4331:78 lut_35.scala 4358:45]
  wire  _GEN_10063 = read_stack17_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10040; // @[lut_35.scala 4331:78 lut_35.scala 4359:45]
  wire  _GEN_10064 = read_stack17_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10041; // @[lut_35.scala 4331:78 lut_35.scala 4360:45]
  wire  _GEN_10065 = read_stack17_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10042; // @[lut_35.scala 4331:78 lut_35.scala 4361:45]
  wire  _GEN_10066 = read_stack17_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10043; // @[lut_35.scala 4331:78 lut_35.scala 4362:45]
  wire  _GEN_10067 = read_stack17_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10044; // @[lut_35.scala 4331:78 lut_35.scala 4363:45]
  wire  _GEN_10068 = read_stack17_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10045; // @[lut_35.scala 4331:78 lut_35.scala 4364:45]
  wire  _GEN_10069 = read_stack17_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10046; // @[lut_35.scala 4331:78 lut_35.scala 4365:45]
  wire  _GEN_10070 = read_stack17_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10047; // @[lut_35.scala 4331:78 lut_35.scala 4366:45]
  wire  _GEN_10071 = read_stack17_pop == pop_ray_id & pop_valid | _GEN_10048; // @[lut_35.scala 4331:78 lut_35.scala 4367:40]
  wire [31:0] _GEN_10073 = read_stack17_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_10050; // @[lut_35.scala 4331:78 lut_35.scala 4369:38]
  wire [31:0] _GEN_10074 = read_stack17_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_10051; // @[lut_35.scala 4331:78 lut_35.scala 4370:41]
  wire  _GEN_10077 = read_stack16_pop == pop_ray_id & pop_valid ? 1'h0 : _T_697; // @[lut_35.scala 4291:78 lut_35.scala 4309:45]
  wire  _GEN_10078 = read_stack16_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10054; // @[lut_35.scala 4291:78 lut_35.scala 4310:45]
  wire  _GEN_10079 = read_stack16_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10055; // @[lut_35.scala 4291:78 lut_35.scala 4311:45]
  wire  _GEN_10080 = read_stack16_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10056; // @[lut_35.scala 4291:78 lut_35.scala 4312:45]
  wire  _GEN_10081 = read_stack16_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10057; // @[lut_35.scala 4291:78 lut_35.scala 4313:45]
  wire  _GEN_10082 = read_stack16_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10058; // @[lut_35.scala 4291:78 lut_35.scala 4314:45]
  wire  _GEN_10083 = read_stack16_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10059; // @[lut_35.scala 4291:78 lut_35.scala 4315:45]
  wire  _GEN_10084 = read_stack16_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10060; // @[lut_35.scala 4291:78 lut_35.scala 4316:45]
  wire  _GEN_10085 = read_stack16_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10061; // @[lut_35.scala 4291:78 lut_35.scala 4317:45]
  wire  _GEN_10086 = read_stack16_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10062; // @[lut_35.scala 4291:78 lut_35.scala 4318:45]
  wire  _GEN_10087 = read_stack16_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10063; // @[lut_35.scala 4291:78 lut_35.scala 4319:45]
  wire  _GEN_10088 = read_stack16_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10064; // @[lut_35.scala 4291:78 lut_35.scala 4320:45]
  wire  _GEN_10089 = read_stack16_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10065; // @[lut_35.scala 4291:78 lut_35.scala 4321:45]
  wire  _GEN_10090 = read_stack16_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10066; // @[lut_35.scala 4291:78 lut_35.scala 4322:45]
  wire  _GEN_10091 = read_stack16_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10067; // @[lut_35.scala 4291:78 lut_35.scala 4323:45]
  wire  _GEN_10092 = read_stack16_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10068; // @[lut_35.scala 4291:78 lut_35.scala 4324:45]
  wire  _GEN_10093 = read_stack16_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10069; // @[lut_35.scala 4291:78 lut_35.scala 4325:45]
  wire  _GEN_10094 = read_stack16_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10070; // @[lut_35.scala 4291:78 lut_35.scala 4326:45]
  wire  _GEN_10095 = read_stack16_pop == pop_ray_id & pop_valid | _GEN_10071; // @[lut_35.scala 4291:78 lut_35.scala 4327:40]
  wire [31:0] _GEN_10097 = read_stack16_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_10073; // @[lut_35.scala 4291:78 lut_35.scala 4329:38]
  wire [31:0] _GEN_10098 = read_stack16_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_10074; // @[lut_35.scala 4291:78 lut_35.scala 4330:41]
  wire  _GEN_10101 = read_stack15_pop == pop_ray_id & pop_valid ? 1'h0 : _T_694; // @[lut_35.scala 4251:78 lut_35.scala 4268:45]
  wire  _GEN_10102 = read_stack15_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10077; // @[lut_35.scala 4251:78 lut_35.scala 4269:45]
  wire  _GEN_10103 = read_stack15_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10078; // @[lut_35.scala 4251:78 lut_35.scala 4270:45]
  wire  _GEN_10104 = read_stack15_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10079; // @[lut_35.scala 4251:78 lut_35.scala 4271:45]
  wire  _GEN_10105 = read_stack15_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10080; // @[lut_35.scala 4251:78 lut_35.scala 4272:45]
  wire  _GEN_10106 = read_stack15_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10081; // @[lut_35.scala 4251:78 lut_35.scala 4273:45]
  wire  _GEN_10107 = read_stack15_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10082; // @[lut_35.scala 4251:78 lut_35.scala 4274:45]
  wire  _GEN_10108 = read_stack15_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10083; // @[lut_35.scala 4251:78 lut_35.scala 4275:45]
  wire  _GEN_10109 = read_stack15_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10084; // @[lut_35.scala 4251:78 lut_35.scala 4276:45]
  wire  _GEN_10110 = read_stack15_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10085; // @[lut_35.scala 4251:78 lut_35.scala 4277:45]
  wire  _GEN_10111 = read_stack15_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10086; // @[lut_35.scala 4251:78 lut_35.scala 4278:45]
  wire  _GEN_10112 = read_stack15_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10087; // @[lut_35.scala 4251:78 lut_35.scala 4279:45]
  wire  _GEN_10113 = read_stack15_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10088; // @[lut_35.scala 4251:78 lut_35.scala 4280:45]
  wire  _GEN_10114 = read_stack15_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10089; // @[lut_35.scala 4251:78 lut_35.scala 4281:45]
  wire  _GEN_10115 = read_stack15_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10090; // @[lut_35.scala 4251:78 lut_35.scala 4282:45]
  wire  _GEN_10116 = read_stack15_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10091; // @[lut_35.scala 4251:78 lut_35.scala 4283:45]
  wire  _GEN_10117 = read_stack15_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10092; // @[lut_35.scala 4251:78 lut_35.scala 4284:45]
  wire  _GEN_10118 = read_stack15_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10093; // @[lut_35.scala 4251:78 lut_35.scala 4285:45]
  wire  _GEN_10119 = read_stack15_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10094; // @[lut_35.scala 4251:78 lut_35.scala 4286:45]
  wire  _GEN_10120 = read_stack15_pop == pop_ray_id & pop_valid | _GEN_10095; // @[lut_35.scala 4251:78 lut_35.scala 4287:40]
  wire [31:0] _GEN_10122 = read_stack15_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_10097; // @[lut_35.scala 4251:78 lut_35.scala 4289:38]
  wire [31:0] _GEN_10123 = read_stack15_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_10098; // @[lut_35.scala 4251:78 lut_35.scala 4290:41]
  wire  _GEN_10126 = read_stack14_pop == pop_ray_id & pop_valid ? 1'h0 : _T_691; // @[lut_35.scala 4211:78 lut_35.scala 4227:45]
  wire  _GEN_10127 = read_stack14_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10101; // @[lut_35.scala 4211:78 lut_35.scala 4228:45]
  wire  _GEN_10128 = read_stack14_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10102; // @[lut_35.scala 4211:78 lut_35.scala 4229:45]
  wire  _GEN_10129 = read_stack14_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10103; // @[lut_35.scala 4211:78 lut_35.scala 4230:45]
  wire  _GEN_10130 = read_stack14_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10104; // @[lut_35.scala 4211:78 lut_35.scala 4231:45]
  wire  _GEN_10131 = read_stack14_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10105; // @[lut_35.scala 4211:78 lut_35.scala 4232:45]
  wire  _GEN_10132 = read_stack14_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10106; // @[lut_35.scala 4211:78 lut_35.scala 4233:45]
  wire  _GEN_10133 = read_stack14_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10107; // @[lut_35.scala 4211:78 lut_35.scala 4234:45]
  wire  _GEN_10134 = read_stack14_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10108; // @[lut_35.scala 4211:78 lut_35.scala 4235:45]
  wire  _GEN_10135 = read_stack14_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10109; // @[lut_35.scala 4211:78 lut_35.scala 4236:45]
  wire  _GEN_10136 = read_stack14_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10110; // @[lut_35.scala 4211:78 lut_35.scala 4237:45]
  wire  _GEN_10137 = read_stack14_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10111; // @[lut_35.scala 4211:78 lut_35.scala 4238:45]
  wire  _GEN_10138 = read_stack14_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10112; // @[lut_35.scala 4211:78 lut_35.scala 4239:45]
  wire  _GEN_10139 = read_stack14_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10113; // @[lut_35.scala 4211:78 lut_35.scala 4240:45]
  wire  _GEN_10140 = read_stack14_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10114; // @[lut_35.scala 4211:78 lut_35.scala 4241:45]
  wire  _GEN_10141 = read_stack14_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10115; // @[lut_35.scala 4211:78 lut_35.scala 4242:45]
  wire  _GEN_10142 = read_stack14_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10116; // @[lut_35.scala 4211:78 lut_35.scala 4243:45]
  wire  _GEN_10143 = read_stack14_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10117; // @[lut_35.scala 4211:78 lut_35.scala 4244:45]
  wire  _GEN_10144 = read_stack14_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10118; // @[lut_35.scala 4211:78 lut_35.scala 4245:45]
  wire  _GEN_10145 = read_stack14_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10119; // @[lut_35.scala 4211:78 lut_35.scala 4246:45]
  wire  _GEN_10146 = read_stack14_pop == pop_ray_id & pop_valid | _GEN_10120; // @[lut_35.scala 4211:78 lut_35.scala 4247:40]
  wire [31:0] _GEN_10148 = read_stack14_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_10122; // @[lut_35.scala 4211:78 lut_35.scala 4249:38]
  wire [31:0] _GEN_10149 = read_stack14_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_10123; // @[lut_35.scala 4211:78 lut_35.scala 4250:41]
  wire  _GEN_10152 = read_stack13_pop == pop_ray_id & pop_valid ? 1'h0 : _T_688; // @[lut_35.scala 4171:78 lut_35.scala 4186:45]
  wire  _GEN_10153 = read_stack13_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10126; // @[lut_35.scala 4171:78 lut_35.scala 4187:45]
  wire  _GEN_10154 = read_stack13_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10127; // @[lut_35.scala 4171:78 lut_35.scala 4188:45]
  wire  _GEN_10155 = read_stack13_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10128; // @[lut_35.scala 4171:78 lut_35.scala 4189:45]
  wire  _GEN_10156 = read_stack13_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10129; // @[lut_35.scala 4171:78 lut_35.scala 4190:45]
  wire  _GEN_10157 = read_stack13_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10130; // @[lut_35.scala 4171:78 lut_35.scala 4191:45]
  wire  _GEN_10158 = read_stack13_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10131; // @[lut_35.scala 4171:78 lut_35.scala 4192:45]
  wire  _GEN_10159 = read_stack13_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10132; // @[lut_35.scala 4171:78 lut_35.scala 4193:45]
  wire  _GEN_10160 = read_stack13_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10133; // @[lut_35.scala 4171:78 lut_35.scala 4194:45]
  wire  _GEN_10161 = read_stack13_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10134; // @[lut_35.scala 4171:78 lut_35.scala 4195:45]
  wire  _GEN_10162 = read_stack13_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10135; // @[lut_35.scala 4171:78 lut_35.scala 4196:45]
  wire  _GEN_10163 = read_stack13_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10136; // @[lut_35.scala 4171:78 lut_35.scala 4197:45]
  wire  _GEN_10164 = read_stack13_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10137; // @[lut_35.scala 4171:78 lut_35.scala 4198:45]
  wire  _GEN_10165 = read_stack13_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10138; // @[lut_35.scala 4171:78 lut_35.scala 4199:45]
  wire  _GEN_10166 = read_stack13_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10139; // @[lut_35.scala 4171:78 lut_35.scala 4200:45]
  wire  _GEN_10167 = read_stack13_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10140; // @[lut_35.scala 4171:78 lut_35.scala 4201:45]
  wire  _GEN_10168 = read_stack13_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10141; // @[lut_35.scala 4171:78 lut_35.scala 4202:45]
  wire  _GEN_10169 = read_stack13_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10142; // @[lut_35.scala 4171:78 lut_35.scala 4203:45]
  wire  _GEN_10170 = read_stack13_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10143; // @[lut_35.scala 4171:78 lut_35.scala 4204:45]
  wire  _GEN_10171 = read_stack13_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10144; // @[lut_35.scala 4171:78 lut_35.scala 4205:45]
  wire  _GEN_10172 = read_stack13_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10145; // @[lut_35.scala 4171:78 lut_35.scala 4206:45]
  wire  _GEN_10173 = read_stack13_pop == pop_ray_id & pop_valid | _GEN_10146; // @[lut_35.scala 4171:78 lut_35.scala 4207:40]
  wire [31:0] _GEN_10175 = read_stack13_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_10148; // @[lut_35.scala 4171:78 lut_35.scala 4209:38]
  wire [31:0] _GEN_10176 = read_stack13_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_10149; // @[lut_35.scala 4171:78 lut_35.scala 4210:41]
  wire  _GEN_10179 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _T_685; // @[lut_35.scala 4131:78 lut_35.scala 4145:45]
  wire  _GEN_10180 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10152; // @[lut_35.scala 4131:78 lut_35.scala 4146:45]
  wire  _GEN_10181 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10153; // @[lut_35.scala 4131:78 lut_35.scala 4147:45]
  wire  _GEN_10182 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10154; // @[lut_35.scala 4131:78 lut_35.scala 4148:45]
  wire  _GEN_10183 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10155; // @[lut_35.scala 4131:78 lut_35.scala 4149:45]
  wire  _GEN_10184 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10156; // @[lut_35.scala 4131:78 lut_35.scala 4150:45]
  wire  _GEN_10185 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10157; // @[lut_35.scala 4131:78 lut_35.scala 4151:45]
  wire  _GEN_10186 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10158; // @[lut_35.scala 4131:78 lut_35.scala 4152:45]
  wire  _GEN_10187 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10159; // @[lut_35.scala 4131:78 lut_35.scala 4153:45]
  wire  _GEN_10188 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10160; // @[lut_35.scala 4131:78 lut_35.scala 4154:45]
  wire  _GEN_10189 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10161; // @[lut_35.scala 4131:78 lut_35.scala 4155:45]
  wire  _GEN_10190 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10162; // @[lut_35.scala 4131:78 lut_35.scala 4156:45]
  wire  _GEN_10191 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10163; // @[lut_35.scala 4131:78 lut_35.scala 4157:45]
  wire  _GEN_10192 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10164; // @[lut_35.scala 4131:78 lut_35.scala 4158:45]
  wire  _GEN_10193 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10165; // @[lut_35.scala 4131:78 lut_35.scala 4159:45]
  wire  _GEN_10194 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10166; // @[lut_35.scala 4131:78 lut_35.scala 4160:45]
  wire  _GEN_10195 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10167; // @[lut_35.scala 4131:78 lut_35.scala 4161:45]
  wire  _GEN_10196 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10168; // @[lut_35.scala 4131:78 lut_35.scala 4162:45]
  wire  _GEN_10197 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10169; // @[lut_35.scala 4131:78 lut_35.scala 4163:45]
  wire  _GEN_10198 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10170; // @[lut_35.scala 4131:78 lut_35.scala 4164:45]
  wire  _GEN_10199 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10171; // @[lut_35.scala 4131:78 lut_35.scala 4165:45]
  wire  _GEN_10200 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10172; // @[lut_35.scala 4131:78 lut_35.scala 4166:45]
  wire  _GEN_10201 = read_stack12_pop == pop_ray_id & pop_valid | _GEN_10173; // @[lut_35.scala 4131:78 lut_35.scala 4167:40]
  wire [31:0] _GEN_10203 = read_stack12_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_10175; // @[lut_35.scala 4131:78 lut_35.scala 4169:38]
  wire [31:0] _GEN_10204 = read_stack12_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_10176; // @[lut_35.scala 4131:78 lut_35.scala 4170:41]
  wire  _GEN_10207 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _T_682; // @[lut_35.scala 4091:78 lut_35.scala 4104:45]
  wire  _GEN_10208 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10179; // @[lut_35.scala 4091:78 lut_35.scala 4105:45]
  wire  _GEN_10209 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10180; // @[lut_35.scala 4091:78 lut_35.scala 4106:45]
  wire  _GEN_10210 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10181; // @[lut_35.scala 4091:78 lut_35.scala 4107:45]
  wire  _GEN_10211 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10182; // @[lut_35.scala 4091:78 lut_35.scala 4108:45]
  wire  _GEN_10212 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10183; // @[lut_35.scala 4091:78 lut_35.scala 4109:45]
  wire  _GEN_10213 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10184; // @[lut_35.scala 4091:78 lut_35.scala 4110:45]
  wire  _GEN_10214 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10185; // @[lut_35.scala 4091:78 lut_35.scala 4111:45]
  wire  _GEN_10215 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10186; // @[lut_35.scala 4091:78 lut_35.scala 4112:45]
  wire  _GEN_10216 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10187; // @[lut_35.scala 4091:78 lut_35.scala 4113:45]
  wire  _GEN_10217 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10188; // @[lut_35.scala 4091:78 lut_35.scala 4114:45]
  wire  _GEN_10218 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10189; // @[lut_35.scala 4091:78 lut_35.scala 4115:45]
  wire  _GEN_10219 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10190; // @[lut_35.scala 4091:78 lut_35.scala 4116:45]
  wire  _GEN_10220 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10191; // @[lut_35.scala 4091:78 lut_35.scala 4117:45]
  wire  _GEN_10221 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10192; // @[lut_35.scala 4091:78 lut_35.scala 4118:45]
  wire  _GEN_10222 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10193; // @[lut_35.scala 4091:78 lut_35.scala 4119:45]
  wire  _GEN_10223 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10194; // @[lut_35.scala 4091:78 lut_35.scala 4120:45]
  wire  _GEN_10224 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10195; // @[lut_35.scala 4091:78 lut_35.scala 4121:45]
  wire  _GEN_10225 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10196; // @[lut_35.scala 4091:78 lut_35.scala 4122:45]
  wire  _GEN_10226 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10197; // @[lut_35.scala 4091:78 lut_35.scala 4123:45]
  wire  _GEN_10227 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10198; // @[lut_35.scala 4091:78 lut_35.scala 4124:45]
  wire  _GEN_10228 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10199; // @[lut_35.scala 4091:78 lut_35.scala 4125:45]
  wire  _GEN_10229 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10200; // @[lut_35.scala 4091:78 lut_35.scala 4126:45]
  wire  _GEN_10230 = read_stack11_pop == pop_ray_id & pop_valid | _GEN_10201; // @[lut_35.scala 4091:78 lut_35.scala 4127:40]
  wire [31:0] _GEN_10232 = read_stack11_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_10203; // @[lut_35.scala 4091:78 lut_35.scala 4129:38]
  wire [31:0] _GEN_10233 = read_stack11_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_10204; // @[lut_35.scala 4091:78 lut_35.scala 4130:41]
  wire  _GEN_10236 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _T_679; // @[lut_35.scala 4051:78 lut_35.scala 4063:45]
  wire  _GEN_10237 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10207; // @[lut_35.scala 4051:78 lut_35.scala 4064:45]
  wire  _GEN_10238 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10208; // @[lut_35.scala 4051:78 lut_35.scala 4065:45]
  wire  _GEN_10239 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10209; // @[lut_35.scala 4051:78 lut_35.scala 4066:45]
  wire  _GEN_10240 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10210; // @[lut_35.scala 4051:78 lut_35.scala 4067:45]
  wire  _GEN_10241 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10211; // @[lut_35.scala 4051:78 lut_35.scala 4068:45]
  wire  _GEN_10242 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10212; // @[lut_35.scala 4051:78 lut_35.scala 4069:45]
  wire  _GEN_10243 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10213; // @[lut_35.scala 4051:78 lut_35.scala 4070:45]
  wire  _GEN_10244 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10214; // @[lut_35.scala 4051:78 lut_35.scala 4071:45]
  wire  _GEN_10245 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10215; // @[lut_35.scala 4051:78 lut_35.scala 4072:45]
  wire  _GEN_10246 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10216; // @[lut_35.scala 4051:78 lut_35.scala 4073:45]
  wire  _GEN_10247 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10217; // @[lut_35.scala 4051:78 lut_35.scala 4074:45]
  wire  _GEN_10248 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10218; // @[lut_35.scala 4051:78 lut_35.scala 4075:45]
  wire  _GEN_10249 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10219; // @[lut_35.scala 4051:78 lut_35.scala 4076:45]
  wire  _GEN_10250 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10220; // @[lut_35.scala 4051:78 lut_35.scala 4077:45]
  wire  _GEN_10251 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10221; // @[lut_35.scala 4051:78 lut_35.scala 4078:45]
  wire  _GEN_10252 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10222; // @[lut_35.scala 4051:78 lut_35.scala 4079:45]
  wire  _GEN_10253 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10223; // @[lut_35.scala 4051:78 lut_35.scala 4080:45]
  wire  _GEN_10254 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10224; // @[lut_35.scala 4051:78 lut_35.scala 4081:45]
  wire  _GEN_10255 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10225; // @[lut_35.scala 4051:78 lut_35.scala 4082:45]
  wire  _GEN_10256 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10226; // @[lut_35.scala 4051:78 lut_35.scala 4083:45]
  wire  _GEN_10257 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10227; // @[lut_35.scala 4051:78 lut_35.scala 4084:45]
  wire  _GEN_10258 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10228; // @[lut_35.scala 4051:78 lut_35.scala 4085:45]
  wire  _GEN_10259 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10229; // @[lut_35.scala 4051:78 lut_35.scala 4086:45]
  wire  _GEN_10260 = read_stack10_pop == pop_ray_id & pop_valid | _GEN_10230; // @[lut_35.scala 4051:78 lut_35.scala 4087:40]
  wire [31:0] _GEN_10262 = read_stack10_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_10232; // @[lut_35.scala 4051:78 lut_35.scala 4089:38]
  wire [31:0] _GEN_10263 = read_stack10_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_10233; // @[lut_35.scala 4051:78 lut_35.scala 4090:41]
  wire  _GEN_10266 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _T_676; // @[lut_35.scala 4011:77 lut_35.scala 4022:45]
  wire  _GEN_10267 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10236; // @[lut_35.scala 4011:77 lut_35.scala 4023:45]
  wire  _GEN_10268 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10237; // @[lut_35.scala 4011:77 lut_35.scala 4024:45]
  wire  _GEN_10269 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10238; // @[lut_35.scala 4011:77 lut_35.scala 4025:45]
  wire  _GEN_10270 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10239; // @[lut_35.scala 4011:77 lut_35.scala 4026:45]
  wire  _GEN_10271 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10240; // @[lut_35.scala 4011:77 lut_35.scala 4027:45]
  wire  _GEN_10272 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10241; // @[lut_35.scala 4011:77 lut_35.scala 4028:45]
  wire  _GEN_10273 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10242; // @[lut_35.scala 4011:77 lut_35.scala 4029:45]
  wire  _GEN_10274 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10243; // @[lut_35.scala 4011:77 lut_35.scala 4030:45]
  wire  _GEN_10275 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10244; // @[lut_35.scala 4011:77 lut_35.scala 4031:45]
  wire  _GEN_10276 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10245; // @[lut_35.scala 4011:77 lut_35.scala 4032:45]
  wire  _GEN_10277 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10246; // @[lut_35.scala 4011:77 lut_35.scala 4033:45]
  wire  _GEN_10278 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10247; // @[lut_35.scala 4011:77 lut_35.scala 4034:45]
  wire  _GEN_10279 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10248; // @[lut_35.scala 4011:77 lut_35.scala 4035:45]
  wire  _GEN_10280 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10249; // @[lut_35.scala 4011:77 lut_35.scala 4036:45]
  wire  _GEN_10281 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10250; // @[lut_35.scala 4011:77 lut_35.scala 4037:45]
  wire  _GEN_10282 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10251; // @[lut_35.scala 4011:77 lut_35.scala 4038:45]
  wire  _GEN_10283 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10252; // @[lut_35.scala 4011:77 lut_35.scala 4039:45]
  wire  _GEN_10284 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10253; // @[lut_35.scala 4011:77 lut_35.scala 4040:45]
  wire  _GEN_10285 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10254; // @[lut_35.scala 4011:77 lut_35.scala 4041:45]
  wire  _GEN_10286 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10255; // @[lut_35.scala 4011:77 lut_35.scala 4042:45]
  wire  _GEN_10287 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10256; // @[lut_35.scala 4011:77 lut_35.scala 4043:45]
  wire  _GEN_10288 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10257; // @[lut_35.scala 4011:77 lut_35.scala 4044:45]
  wire  _GEN_10289 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10258; // @[lut_35.scala 4011:77 lut_35.scala 4045:45]
  wire  _GEN_10290 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10259; // @[lut_35.scala 4011:77 lut_35.scala 4046:45]
  wire  _GEN_10291 = read_stack9_pop == pop_ray_id & pop_valid | _GEN_10260; // @[lut_35.scala 4011:77 lut_35.scala 4047:40]
  wire [31:0] _GEN_10293 = read_stack9_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_10262; // @[lut_35.scala 4011:77 lut_35.scala 4049:38]
  wire [31:0] _GEN_10294 = read_stack9_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_10263; // @[lut_35.scala 4011:77 lut_35.scala 4050:41]
  wire  _GEN_10297 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _T_673; // @[lut_35.scala 3970:77 lut_35.scala 3980:44]
  wire  _GEN_10298 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10266; // @[lut_35.scala 3970:77 lut_35.scala 3981:45]
  wire  _GEN_10299 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10267; // @[lut_35.scala 3970:77 lut_35.scala 3982:45]
  wire  _GEN_10300 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10268; // @[lut_35.scala 3970:77 lut_35.scala 3983:45]
  wire  _GEN_10301 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10269; // @[lut_35.scala 3970:77 lut_35.scala 3984:45]
  wire  _GEN_10302 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10270; // @[lut_35.scala 3970:77 lut_35.scala 3985:45]
  wire  _GEN_10303 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10271; // @[lut_35.scala 3970:77 lut_35.scala 3986:45]
  wire  _GEN_10304 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10272; // @[lut_35.scala 3970:77 lut_35.scala 3987:45]
  wire  _GEN_10305 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10273; // @[lut_35.scala 3970:77 lut_35.scala 3988:45]
  wire  _GEN_10306 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10274; // @[lut_35.scala 3970:77 lut_35.scala 3989:45]
  wire  _GEN_10307 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10275; // @[lut_35.scala 3970:77 lut_35.scala 3990:45]
  wire  _GEN_10308 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10276; // @[lut_35.scala 3970:77 lut_35.scala 3991:45]
  wire  _GEN_10309 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10277; // @[lut_35.scala 3970:77 lut_35.scala 3992:45]
  wire  _GEN_10310 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10278; // @[lut_35.scala 3970:77 lut_35.scala 3993:45]
  wire  _GEN_10311 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10279; // @[lut_35.scala 3970:77 lut_35.scala 3994:45]
  wire  _GEN_10312 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10280; // @[lut_35.scala 3970:77 lut_35.scala 3995:45]
  wire  _GEN_10313 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10281; // @[lut_35.scala 3970:77 lut_35.scala 3996:45]
  wire  _GEN_10314 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10282; // @[lut_35.scala 3970:77 lut_35.scala 3997:45]
  wire  _GEN_10315 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10283; // @[lut_35.scala 3970:77 lut_35.scala 3998:45]
  wire  _GEN_10316 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10284; // @[lut_35.scala 3970:77 lut_35.scala 3999:45]
  wire  _GEN_10317 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10285; // @[lut_35.scala 3970:77 lut_35.scala 4000:45]
  wire  _GEN_10318 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10286; // @[lut_35.scala 3970:77 lut_35.scala 4001:45]
  wire  _GEN_10319 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10287; // @[lut_35.scala 3970:77 lut_35.scala 4002:45]
  wire  _GEN_10320 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10288; // @[lut_35.scala 3970:77 lut_35.scala 4003:45]
  wire  _GEN_10321 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10289; // @[lut_35.scala 3970:77 lut_35.scala 4004:45]
  wire  _GEN_10322 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10290; // @[lut_35.scala 3970:77 lut_35.scala 4005:45]
  wire  _GEN_10323 = read_stack8_pop == pop_ray_id & pop_valid | _GEN_10291; // @[lut_35.scala 3970:77 lut_35.scala 4006:40]
  wire [31:0] _GEN_10325 = read_stack8_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_10293; // @[lut_35.scala 3970:77 lut_35.scala 4008:38]
  wire [31:0] _GEN_10326 = read_stack8_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_10294; // @[lut_35.scala 3970:77 lut_35.scala 4009:41]
  wire  _GEN_10329 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _T_670; // @[lut_35.scala 3930:77 lut_35.scala 3939:44]
  wire  _GEN_10330 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10297; // @[lut_35.scala 3930:77 lut_35.scala 3940:44]
  wire  _GEN_10331 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10298; // @[lut_35.scala 3930:77 lut_35.scala 3941:45]
  wire  _GEN_10332 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10299; // @[lut_35.scala 3930:77 lut_35.scala 3942:45]
  wire  _GEN_10333 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10300; // @[lut_35.scala 3930:77 lut_35.scala 3943:45]
  wire  _GEN_10334 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10301; // @[lut_35.scala 3930:77 lut_35.scala 3944:45]
  wire  _GEN_10335 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10302; // @[lut_35.scala 3930:77 lut_35.scala 3945:45]
  wire  _GEN_10336 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10303; // @[lut_35.scala 3930:77 lut_35.scala 3946:45]
  wire  _GEN_10337 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10304; // @[lut_35.scala 3930:77 lut_35.scala 3947:45]
  wire  _GEN_10338 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10305; // @[lut_35.scala 3930:77 lut_35.scala 3948:45]
  wire  _GEN_10339 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10306; // @[lut_35.scala 3930:77 lut_35.scala 3949:45]
  wire  _GEN_10340 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10307; // @[lut_35.scala 3930:77 lut_35.scala 3950:45]
  wire  _GEN_10341 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10308; // @[lut_35.scala 3930:77 lut_35.scala 3951:45]
  wire  _GEN_10342 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10309; // @[lut_35.scala 3930:77 lut_35.scala 3952:45]
  wire  _GEN_10343 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10310; // @[lut_35.scala 3930:77 lut_35.scala 3953:45]
  wire  _GEN_10344 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10311; // @[lut_35.scala 3930:77 lut_35.scala 3954:45]
  wire  _GEN_10345 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10312; // @[lut_35.scala 3930:77 lut_35.scala 3955:45]
  wire  _GEN_10346 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10313; // @[lut_35.scala 3930:77 lut_35.scala 3956:45]
  wire  _GEN_10347 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10314; // @[lut_35.scala 3930:77 lut_35.scala 3957:45]
  wire  _GEN_10348 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10315; // @[lut_35.scala 3930:77 lut_35.scala 3958:45]
  wire  _GEN_10349 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10316; // @[lut_35.scala 3930:77 lut_35.scala 3959:45]
  wire  _GEN_10350 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10317; // @[lut_35.scala 3930:77 lut_35.scala 3960:45]
  wire  _GEN_10351 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10318; // @[lut_35.scala 3930:77 lut_35.scala 3961:45]
  wire  _GEN_10352 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10319; // @[lut_35.scala 3930:77 lut_35.scala 3962:45]
  wire  _GEN_10353 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10320; // @[lut_35.scala 3930:77 lut_35.scala 3963:45]
  wire  _GEN_10354 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10321; // @[lut_35.scala 3930:77 lut_35.scala 3964:45]
  wire  _GEN_10355 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10322; // @[lut_35.scala 3930:77 lut_35.scala 3965:45]
  wire  _GEN_10356 = read_stack7_pop == pop_ray_id & pop_valid | _GEN_10323; // @[lut_35.scala 3930:77 lut_35.scala 3966:40]
  wire [31:0] _GEN_10358 = read_stack7_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_10325; // @[lut_35.scala 3930:77 lut_35.scala 3968:38]
  wire [31:0] _GEN_10359 = read_stack7_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_10326; // @[lut_35.scala 3930:77 lut_35.scala 3969:41]
  wire  _GEN_10362 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _T_667; // @[lut_35.scala 3890:77 lut_35.scala 3898:44]
  wire  _GEN_10363 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10329; // @[lut_35.scala 3890:77 lut_35.scala 3899:44]
  wire  _GEN_10364 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10330; // @[lut_35.scala 3890:77 lut_35.scala 3900:44]
  wire  _GEN_10365 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10331; // @[lut_35.scala 3890:77 lut_35.scala 3901:45]
  wire  _GEN_10366 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10332; // @[lut_35.scala 3890:77 lut_35.scala 3902:45]
  wire  _GEN_10367 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10333; // @[lut_35.scala 3890:77 lut_35.scala 3903:45]
  wire  _GEN_10368 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10334; // @[lut_35.scala 3890:77 lut_35.scala 3904:45]
  wire  _GEN_10369 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10335; // @[lut_35.scala 3890:77 lut_35.scala 3905:45]
  wire  _GEN_10370 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10336; // @[lut_35.scala 3890:77 lut_35.scala 3906:45]
  wire  _GEN_10371 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10337; // @[lut_35.scala 3890:77 lut_35.scala 3907:45]
  wire  _GEN_10372 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10338; // @[lut_35.scala 3890:77 lut_35.scala 3908:45]
  wire  _GEN_10373 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10339; // @[lut_35.scala 3890:77 lut_35.scala 3909:45]
  wire  _GEN_10374 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10340; // @[lut_35.scala 3890:77 lut_35.scala 3910:45]
  wire  _GEN_10375 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10341; // @[lut_35.scala 3890:77 lut_35.scala 3911:45]
  wire  _GEN_10376 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10342; // @[lut_35.scala 3890:77 lut_35.scala 3912:45]
  wire  _GEN_10377 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10343; // @[lut_35.scala 3890:77 lut_35.scala 3913:45]
  wire  _GEN_10378 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10344; // @[lut_35.scala 3890:77 lut_35.scala 3914:45]
  wire  _GEN_10379 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10345; // @[lut_35.scala 3890:77 lut_35.scala 3915:45]
  wire  _GEN_10380 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10346; // @[lut_35.scala 3890:77 lut_35.scala 3916:45]
  wire  _GEN_10381 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10347; // @[lut_35.scala 3890:77 lut_35.scala 3917:45]
  wire  _GEN_10382 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10348; // @[lut_35.scala 3890:77 lut_35.scala 3918:45]
  wire  _GEN_10383 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10349; // @[lut_35.scala 3890:77 lut_35.scala 3919:45]
  wire  _GEN_10384 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10350; // @[lut_35.scala 3890:77 lut_35.scala 3920:45]
  wire  _GEN_10385 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10351; // @[lut_35.scala 3890:77 lut_35.scala 3921:45]
  wire  _GEN_10386 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10352; // @[lut_35.scala 3890:77 lut_35.scala 3922:45]
  wire  _GEN_10387 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10353; // @[lut_35.scala 3890:77 lut_35.scala 3923:45]
  wire  _GEN_10388 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10354; // @[lut_35.scala 3890:77 lut_35.scala 3924:45]
  wire  _GEN_10389 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10355; // @[lut_35.scala 3890:77 lut_35.scala 3925:45]
  wire  _GEN_10390 = read_stack6_pop == pop_ray_id & pop_valid | _GEN_10356; // @[lut_35.scala 3890:77 lut_35.scala 3926:40]
  wire [31:0] _GEN_10392 = read_stack6_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_10358; // @[lut_35.scala 3890:77 lut_35.scala 3928:38]
  wire [31:0] _GEN_10393 = read_stack6_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_10359; // @[lut_35.scala 3890:77 lut_35.scala 3929:41]
  wire  _GEN_10396 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _T_664; // @[lut_35.scala 3850:77 lut_35.scala 3857:44]
  wire  _GEN_10397 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10362; // @[lut_35.scala 3850:77 lut_35.scala 3858:44]
  wire  _GEN_10398 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10363; // @[lut_35.scala 3850:77 lut_35.scala 3859:44]
  wire  _GEN_10399 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10364; // @[lut_35.scala 3850:77 lut_35.scala 3860:44]
  wire  _GEN_10400 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10365; // @[lut_35.scala 3850:77 lut_35.scala 3861:45]
  wire  _GEN_10401 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10366; // @[lut_35.scala 3850:77 lut_35.scala 3862:45]
  wire  _GEN_10402 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10367; // @[lut_35.scala 3850:77 lut_35.scala 3863:45]
  wire  _GEN_10403 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10368; // @[lut_35.scala 3850:77 lut_35.scala 3864:45]
  wire  _GEN_10404 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10369; // @[lut_35.scala 3850:77 lut_35.scala 3865:45]
  wire  _GEN_10405 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10370; // @[lut_35.scala 3850:77 lut_35.scala 3866:45]
  wire  _GEN_10406 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10371; // @[lut_35.scala 3850:77 lut_35.scala 3867:45]
  wire  _GEN_10407 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10372; // @[lut_35.scala 3850:77 lut_35.scala 3868:45]
  wire  _GEN_10408 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10373; // @[lut_35.scala 3850:77 lut_35.scala 3869:45]
  wire  _GEN_10409 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10374; // @[lut_35.scala 3850:77 lut_35.scala 3870:45]
  wire  _GEN_10410 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10375; // @[lut_35.scala 3850:77 lut_35.scala 3871:45]
  wire  _GEN_10411 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10376; // @[lut_35.scala 3850:77 lut_35.scala 3872:45]
  wire  _GEN_10412 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10377; // @[lut_35.scala 3850:77 lut_35.scala 3873:45]
  wire  _GEN_10413 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10378; // @[lut_35.scala 3850:77 lut_35.scala 3874:45]
  wire  _GEN_10414 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10379; // @[lut_35.scala 3850:77 lut_35.scala 3875:45]
  wire  _GEN_10415 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10380; // @[lut_35.scala 3850:77 lut_35.scala 3876:45]
  wire  _GEN_10416 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10381; // @[lut_35.scala 3850:77 lut_35.scala 3877:45]
  wire  _GEN_10417 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10382; // @[lut_35.scala 3850:77 lut_35.scala 3878:45]
  wire  _GEN_10418 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10383; // @[lut_35.scala 3850:77 lut_35.scala 3879:45]
  wire  _GEN_10419 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10384; // @[lut_35.scala 3850:77 lut_35.scala 3880:45]
  wire  _GEN_10420 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10385; // @[lut_35.scala 3850:77 lut_35.scala 3881:45]
  wire  _GEN_10421 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10386; // @[lut_35.scala 3850:77 lut_35.scala 3882:45]
  wire  _GEN_10422 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10387; // @[lut_35.scala 3850:77 lut_35.scala 3883:45]
  wire  _GEN_10423 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10388; // @[lut_35.scala 3850:77 lut_35.scala 3884:45]
  wire  _GEN_10424 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10389; // @[lut_35.scala 3850:77 lut_35.scala 3885:45]
  wire  _GEN_10425 = read_stack5_pop == pop_ray_id & pop_valid | _GEN_10390; // @[lut_35.scala 3850:77 lut_35.scala 3886:40]
  wire [31:0] _GEN_10427 = read_stack5_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_10392; // @[lut_35.scala 3850:77 lut_35.scala 3888:38]
  wire [31:0] _GEN_10428 = read_stack5_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_10393; // @[lut_35.scala 3850:77 lut_35.scala 3889:41]
  wire  _GEN_10431 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _T_661; // @[lut_35.scala 3810:77 lut_35.scala 3816:44]
  wire  _GEN_10432 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10396; // @[lut_35.scala 3810:77 lut_35.scala 3817:44]
  wire  _GEN_10433 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10397; // @[lut_35.scala 3810:77 lut_35.scala 3818:44]
  wire  _GEN_10434 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10398; // @[lut_35.scala 3810:77 lut_35.scala 3819:44]
  wire  _GEN_10435 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10399; // @[lut_35.scala 3810:77 lut_35.scala 3820:44]
  wire  _GEN_10436 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10400; // @[lut_35.scala 3810:77 lut_35.scala 3821:45]
  wire  _GEN_10437 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10401; // @[lut_35.scala 3810:77 lut_35.scala 3822:45]
  wire  _GEN_10438 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10402; // @[lut_35.scala 3810:77 lut_35.scala 3823:45]
  wire  _GEN_10439 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10403; // @[lut_35.scala 3810:77 lut_35.scala 3824:45]
  wire  _GEN_10440 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10404; // @[lut_35.scala 3810:77 lut_35.scala 3825:45]
  wire  _GEN_10441 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10405; // @[lut_35.scala 3810:77 lut_35.scala 3826:45]
  wire  _GEN_10442 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10406; // @[lut_35.scala 3810:77 lut_35.scala 3827:45]
  wire  _GEN_10443 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10407; // @[lut_35.scala 3810:77 lut_35.scala 3828:45]
  wire  _GEN_10444 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10408; // @[lut_35.scala 3810:77 lut_35.scala 3829:45]
  wire  _GEN_10445 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10409; // @[lut_35.scala 3810:77 lut_35.scala 3830:45]
  wire  _GEN_10446 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10410; // @[lut_35.scala 3810:77 lut_35.scala 3831:45]
  wire  _GEN_10447 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10411; // @[lut_35.scala 3810:77 lut_35.scala 3832:45]
  wire  _GEN_10448 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10412; // @[lut_35.scala 3810:77 lut_35.scala 3833:45]
  wire  _GEN_10449 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10413; // @[lut_35.scala 3810:77 lut_35.scala 3834:45]
  wire  _GEN_10450 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10414; // @[lut_35.scala 3810:77 lut_35.scala 3835:45]
  wire  _GEN_10451 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10415; // @[lut_35.scala 3810:77 lut_35.scala 3836:45]
  wire  _GEN_10452 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10416; // @[lut_35.scala 3810:77 lut_35.scala 3837:45]
  wire  _GEN_10453 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10417; // @[lut_35.scala 3810:77 lut_35.scala 3838:45]
  wire  _GEN_10454 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10418; // @[lut_35.scala 3810:77 lut_35.scala 3839:45]
  wire  _GEN_10455 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10419; // @[lut_35.scala 3810:77 lut_35.scala 3840:45]
  wire  _GEN_10456 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10420; // @[lut_35.scala 3810:77 lut_35.scala 3841:45]
  wire  _GEN_10457 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10421; // @[lut_35.scala 3810:77 lut_35.scala 3842:45]
  wire  _GEN_10458 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10422; // @[lut_35.scala 3810:77 lut_35.scala 3843:45]
  wire  _GEN_10459 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10423; // @[lut_35.scala 3810:77 lut_35.scala 3844:45]
  wire  _GEN_10460 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10424; // @[lut_35.scala 3810:77 lut_35.scala 3845:45]
  wire  _GEN_10461 = read_stack4_pop == pop_ray_id & pop_valid | _GEN_10425; // @[lut_35.scala 3810:77 lut_35.scala 3846:40]
  wire [31:0] _GEN_10463 = read_stack4_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_10427; // @[lut_35.scala 3810:77 lut_35.scala 3848:38]
  wire [31:0] _GEN_10464 = read_stack4_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_10428; // @[lut_35.scala 3810:77 lut_35.scala 3849:41]
  wire  _GEN_10467 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _T_658; // @[lut_35.scala 3770:77 lut_35.scala 3775:44]
  wire  _GEN_10468 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10431; // @[lut_35.scala 3770:77 lut_35.scala 3776:44]
  wire  _GEN_10469 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10432; // @[lut_35.scala 3770:77 lut_35.scala 3777:44]
  wire  _GEN_10470 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10433; // @[lut_35.scala 3770:77 lut_35.scala 3778:44]
  wire  _GEN_10471 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10434; // @[lut_35.scala 3770:77 lut_35.scala 3779:44]
  wire  _GEN_10472 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10435; // @[lut_35.scala 3770:77 lut_35.scala 3780:44]
  wire  _GEN_10473 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10436; // @[lut_35.scala 3770:77 lut_35.scala 3781:45]
  wire  _GEN_10474 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10437; // @[lut_35.scala 3770:77 lut_35.scala 3782:45]
  wire  _GEN_10475 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10438; // @[lut_35.scala 3770:77 lut_35.scala 3783:45]
  wire  _GEN_10476 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10439; // @[lut_35.scala 3770:77 lut_35.scala 3784:45]
  wire  _GEN_10477 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10440; // @[lut_35.scala 3770:77 lut_35.scala 3785:45]
  wire  _GEN_10478 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10441; // @[lut_35.scala 3770:77 lut_35.scala 3786:45]
  wire  _GEN_10479 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10442; // @[lut_35.scala 3770:77 lut_35.scala 3787:45]
  wire  _GEN_10480 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10443; // @[lut_35.scala 3770:77 lut_35.scala 3788:45]
  wire  _GEN_10481 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10444; // @[lut_35.scala 3770:77 lut_35.scala 3789:45]
  wire  _GEN_10482 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10445; // @[lut_35.scala 3770:77 lut_35.scala 3790:45]
  wire  _GEN_10483 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10446; // @[lut_35.scala 3770:77 lut_35.scala 3791:45]
  wire  _GEN_10484 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10447; // @[lut_35.scala 3770:77 lut_35.scala 3792:45]
  wire  _GEN_10485 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10448; // @[lut_35.scala 3770:77 lut_35.scala 3793:45]
  wire  _GEN_10486 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10449; // @[lut_35.scala 3770:77 lut_35.scala 3794:45]
  wire  _GEN_10487 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10450; // @[lut_35.scala 3770:77 lut_35.scala 3795:45]
  wire  _GEN_10488 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10451; // @[lut_35.scala 3770:77 lut_35.scala 3796:45]
  wire  _GEN_10489 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10452; // @[lut_35.scala 3770:77 lut_35.scala 3797:45]
  wire  _GEN_10490 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10453; // @[lut_35.scala 3770:77 lut_35.scala 3798:45]
  wire  _GEN_10491 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10454; // @[lut_35.scala 3770:77 lut_35.scala 3799:45]
  wire  _GEN_10492 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10455; // @[lut_35.scala 3770:77 lut_35.scala 3800:45]
  wire  _GEN_10493 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10456; // @[lut_35.scala 3770:77 lut_35.scala 3801:45]
  wire  _GEN_10494 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10457; // @[lut_35.scala 3770:77 lut_35.scala 3802:45]
  wire  _GEN_10495 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10458; // @[lut_35.scala 3770:77 lut_35.scala 3803:45]
  wire  _GEN_10496 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10459; // @[lut_35.scala 3770:77 lut_35.scala 3804:45]
  wire  _GEN_10497 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10460; // @[lut_35.scala 3770:77 lut_35.scala 3805:45]
  wire  _GEN_10498 = read_stack3_pop == pop_ray_id & pop_valid | _GEN_10461; // @[lut_35.scala 3770:77 lut_35.scala 3806:40]
  wire [31:0] _GEN_10500 = read_stack3_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_10463; // @[lut_35.scala 3770:77 lut_35.scala 3808:38]
  wire [31:0] _GEN_10501 = read_stack3_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_10464; // @[lut_35.scala 3770:77 lut_35.scala 3809:41]
  wire  _GEN_10504 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _T_655; // @[lut_35.scala 3730:77 lut_35.scala 3734:44]
  wire  _GEN_10505 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10467; // @[lut_35.scala 3730:77 lut_35.scala 3735:44]
  wire  _GEN_10506 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10468; // @[lut_35.scala 3730:77 lut_35.scala 3736:44]
  wire  _GEN_10507 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10469; // @[lut_35.scala 3730:77 lut_35.scala 3737:44]
  wire  _GEN_10508 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10470; // @[lut_35.scala 3730:77 lut_35.scala 3738:44]
  wire  _GEN_10509 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10471; // @[lut_35.scala 3730:77 lut_35.scala 3739:44]
  wire  _GEN_10510 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10472; // @[lut_35.scala 3730:77 lut_35.scala 3740:44]
  wire  _GEN_10511 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10473; // @[lut_35.scala 3730:77 lut_35.scala 3741:45]
  wire  _GEN_10512 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10474; // @[lut_35.scala 3730:77 lut_35.scala 3742:45]
  wire  _GEN_10513 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10475; // @[lut_35.scala 3730:77 lut_35.scala 3743:45]
  wire  _GEN_10514 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10476; // @[lut_35.scala 3730:77 lut_35.scala 3744:45]
  wire  _GEN_10515 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10477; // @[lut_35.scala 3730:77 lut_35.scala 3745:45]
  wire  _GEN_10516 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10478; // @[lut_35.scala 3730:77 lut_35.scala 3746:45]
  wire  _GEN_10517 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10479; // @[lut_35.scala 3730:77 lut_35.scala 3747:45]
  wire  _GEN_10518 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10480; // @[lut_35.scala 3730:77 lut_35.scala 3748:45]
  wire  _GEN_10519 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10481; // @[lut_35.scala 3730:77 lut_35.scala 3749:45]
  wire  _GEN_10520 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10482; // @[lut_35.scala 3730:77 lut_35.scala 3750:45]
  wire  _GEN_10521 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10483; // @[lut_35.scala 3730:77 lut_35.scala 3751:45]
  wire  _GEN_10522 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10484; // @[lut_35.scala 3730:77 lut_35.scala 3752:45]
  wire  _GEN_10523 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10485; // @[lut_35.scala 3730:77 lut_35.scala 3753:45]
  wire  _GEN_10524 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10486; // @[lut_35.scala 3730:77 lut_35.scala 3754:45]
  wire  _GEN_10525 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10487; // @[lut_35.scala 3730:77 lut_35.scala 3755:45]
  wire  _GEN_10526 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10488; // @[lut_35.scala 3730:77 lut_35.scala 3756:45]
  wire  _GEN_10527 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10489; // @[lut_35.scala 3730:77 lut_35.scala 3757:45]
  wire  _GEN_10528 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10490; // @[lut_35.scala 3730:77 lut_35.scala 3758:45]
  wire  _GEN_10529 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10491; // @[lut_35.scala 3730:77 lut_35.scala 3759:45]
  wire  _GEN_10530 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10492; // @[lut_35.scala 3730:77 lut_35.scala 3760:45]
  wire  _GEN_10531 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10493; // @[lut_35.scala 3730:77 lut_35.scala 3761:45]
  wire  _GEN_10532 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10494; // @[lut_35.scala 3730:77 lut_35.scala 3762:45]
  wire  _GEN_10533 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10495; // @[lut_35.scala 3730:77 lut_35.scala 3763:45]
  wire  _GEN_10534 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10496; // @[lut_35.scala 3730:77 lut_35.scala 3764:45]
  wire  _GEN_10535 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10497; // @[lut_35.scala 3730:77 lut_35.scala 3765:45]
  wire  _GEN_10536 = read_stack2_pop == pop_ray_id & pop_valid | _GEN_10498; // @[lut_35.scala 3730:77 lut_35.scala 3766:40]
  wire [31:0] _GEN_10538 = read_stack2_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_10500; // @[lut_35.scala 3730:77 lut_35.scala 3768:38]
  wire [31:0] _GEN_10539 = read_stack2_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_10501; // @[lut_35.scala 3730:77 lut_35.scala 3769:41]
  wire  _GEN_10542 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _T_652; // @[lut_35.scala 3690:77 lut_35.scala 3693:44]
  wire  _GEN_10543 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10504; // @[lut_35.scala 3690:77 lut_35.scala 3694:44]
  wire  _GEN_10544 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10505; // @[lut_35.scala 3690:77 lut_35.scala 3695:44]
  wire  _GEN_10545 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10506; // @[lut_35.scala 3690:77 lut_35.scala 3696:44]
  wire  _GEN_10546 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10507; // @[lut_35.scala 3690:77 lut_35.scala 3697:44]
  wire  _GEN_10547 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10508; // @[lut_35.scala 3690:77 lut_35.scala 3698:44]
  wire  _GEN_10548 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10509; // @[lut_35.scala 3690:77 lut_35.scala 3699:44]
  wire  _GEN_10549 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10510; // @[lut_35.scala 3690:77 lut_35.scala 3700:44]
  wire  _GEN_10550 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10511; // @[lut_35.scala 3690:77 lut_35.scala 3701:45]
  wire  _GEN_10551 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10512; // @[lut_35.scala 3690:77 lut_35.scala 3702:45]
  wire  _GEN_10552 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10513; // @[lut_35.scala 3690:77 lut_35.scala 3703:45]
  wire  _GEN_10553 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10514; // @[lut_35.scala 3690:77 lut_35.scala 3704:45]
  wire  _GEN_10554 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10515; // @[lut_35.scala 3690:77 lut_35.scala 3705:45]
  wire  _GEN_10555 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10516; // @[lut_35.scala 3690:77 lut_35.scala 3706:45]
  wire  _GEN_10556 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10517; // @[lut_35.scala 3690:77 lut_35.scala 3707:45]
  wire  _GEN_10557 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10518; // @[lut_35.scala 3690:77 lut_35.scala 3708:45]
  wire  _GEN_10558 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10519; // @[lut_35.scala 3690:77 lut_35.scala 3709:45]
  wire  _GEN_10559 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10520; // @[lut_35.scala 3690:77 lut_35.scala 3710:45]
  wire  _GEN_10560 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10521; // @[lut_35.scala 3690:77 lut_35.scala 3711:45]
  wire  _GEN_10561 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10522; // @[lut_35.scala 3690:77 lut_35.scala 3712:45]
  wire  _GEN_10562 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10523; // @[lut_35.scala 3690:77 lut_35.scala 3713:45]
  wire  _GEN_10563 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10524; // @[lut_35.scala 3690:77 lut_35.scala 3714:45]
  wire  _GEN_10564 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10525; // @[lut_35.scala 3690:77 lut_35.scala 3715:45]
  wire  _GEN_10565 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10526; // @[lut_35.scala 3690:77 lut_35.scala 3716:45]
  wire  _GEN_10566 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10527; // @[lut_35.scala 3690:77 lut_35.scala 3717:45]
  wire  _GEN_10567 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10528; // @[lut_35.scala 3690:77 lut_35.scala 3718:45]
  wire  _GEN_10568 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10529; // @[lut_35.scala 3690:77 lut_35.scala 3719:45]
  wire  _GEN_10569 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10530; // @[lut_35.scala 3690:77 lut_35.scala 3720:45]
  wire  _GEN_10570 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10531; // @[lut_35.scala 3690:77 lut_35.scala 3721:45]
  wire  _GEN_10571 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10532; // @[lut_35.scala 3690:77 lut_35.scala 3722:45]
  wire  _GEN_10572 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10533; // @[lut_35.scala 3690:77 lut_35.scala 3723:45]
  wire  _GEN_10573 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10534; // @[lut_35.scala 3690:77 lut_35.scala 3724:45]
  wire  _GEN_10574 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10535; // @[lut_35.scala 3690:77 lut_35.scala 3725:45]
  wire  _GEN_10575 = read_stack1_pop == pop_ray_id & pop_valid | _GEN_10536; // @[lut_35.scala 3690:77 lut_35.scala 3726:40]
  wire  _GEN_10580 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _T_649; // @[lut_35.scala 3650:67 lut_35.scala 3652:40]
  wire  _GEN_10581 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10542; // @[lut_35.scala 3650:67 lut_35.scala 3653:40]
  wire  _GEN_10582 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10543; // @[lut_35.scala 3650:67 lut_35.scala 3654:40]
  wire  _GEN_10583 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10544; // @[lut_35.scala 3650:67 lut_35.scala 3655:40]
  wire  _GEN_10584 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10545; // @[lut_35.scala 3650:67 lut_35.scala 3656:40]
  wire  _GEN_10585 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10546; // @[lut_35.scala 3650:67 lut_35.scala 3657:40]
  wire  _GEN_10586 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10547; // @[lut_35.scala 3650:67 lut_35.scala 3658:40]
  wire  _GEN_10587 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10548; // @[lut_35.scala 3650:67 lut_35.scala 3659:40]
  wire  _GEN_10588 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10549; // @[lut_35.scala 3650:67 lut_35.scala 3660:40]
  wire  _GEN_10589 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10550; // @[lut_35.scala 3650:67 lut_35.scala 3661:41]
  wire  _GEN_10590 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10551; // @[lut_35.scala 3650:67 lut_35.scala 3662:41]
  wire  _GEN_10591 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10552; // @[lut_35.scala 3650:67 lut_35.scala 3663:41]
  wire  _GEN_10592 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10553; // @[lut_35.scala 3650:67 lut_35.scala 3664:41]
  wire  _GEN_10593 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10554; // @[lut_35.scala 3650:67 lut_35.scala 3665:41]
  wire  _GEN_10594 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10555; // @[lut_35.scala 3650:67 lut_35.scala 3666:41]
  wire  _GEN_10595 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10556; // @[lut_35.scala 3650:67 lut_35.scala 3667:41]
  wire  _GEN_10596 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10557; // @[lut_35.scala 3650:67 lut_35.scala 3668:41]
  wire  _GEN_10597 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10558; // @[lut_35.scala 3650:67 lut_35.scala 3669:41]
  wire  _GEN_10598 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10559; // @[lut_35.scala 3650:67 lut_35.scala 3670:41]
  wire  _GEN_10599 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10560; // @[lut_35.scala 3650:67 lut_35.scala 3671:41]
  wire  _GEN_10600 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10561; // @[lut_35.scala 3650:67 lut_35.scala 3672:41]
  wire  _GEN_10601 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10562; // @[lut_35.scala 3650:67 lut_35.scala 3673:41]
  wire  _GEN_10602 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10563; // @[lut_35.scala 3650:67 lut_35.scala 3674:41]
  wire  _GEN_10603 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10564; // @[lut_35.scala 3650:67 lut_35.scala 3675:41]
  wire  _GEN_10604 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10565; // @[lut_35.scala 3650:67 lut_35.scala 3676:41]
  wire  _GEN_10605 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10566; // @[lut_35.scala 3650:67 lut_35.scala 3677:41]
  wire  _GEN_10606 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10567; // @[lut_35.scala 3650:67 lut_35.scala 3678:41]
  wire  _GEN_10607 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10568; // @[lut_35.scala 3650:67 lut_35.scala 3679:41]
  wire  _GEN_10608 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10569; // @[lut_35.scala 3650:67 lut_35.scala 3680:41]
  wire  _GEN_10609 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10570; // @[lut_35.scala 3650:67 lut_35.scala 3681:41]
  wire  _GEN_10610 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10571; // @[lut_35.scala 3650:67 lut_35.scala 3682:41]
  wire  _GEN_10611 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10572; // @[lut_35.scala 3650:67 lut_35.scala 3683:41]
  wire  _GEN_10612 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10573; // @[lut_35.scala 3650:67 lut_35.scala 3684:41]
  wire  _GEN_10613 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_10574; // @[lut_35.scala 3650:67 lut_35.scala 3685:41]
  wire  _GEN_10614 = read_stack0_pop == pop_ray_id & pop_valid | _GEN_10575; // @[lut_35.scala 3650:67 lut_35.scala 3686:36]
  wire  _GEN_10618 = pop_1 & pop_valid & _T_646; // @[lut_35.scala 3649:46 lut_35.scala 5090:40]
  wire  _GEN_10619 = pop_1 & pop_valid & _GEN_10580; // @[lut_35.scala 3649:46 lut_35.scala 5091:40]
  wire  _GEN_10620 = pop_1 & pop_valid & _GEN_10581; // @[lut_35.scala 3649:46 lut_35.scala 5092:40]
  wire  _GEN_10621 = pop_1 & pop_valid & _GEN_10582; // @[lut_35.scala 3649:46 lut_35.scala 5093:40]
  wire  _GEN_10622 = pop_1 & pop_valid & _GEN_10583; // @[lut_35.scala 3649:46 lut_35.scala 5094:40]
  wire  _GEN_10623 = pop_1 & pop_valid & _GEN_10584; // @[lut_35.scala 3649:46 lut_35.scala 5095:40]
  wire  _GEN_10624 = pop_1 & pop_valid & _GEN_10585; // @[lut_35.scala 3649:46 lut_35.scala 5096:40]
  wire  _GEN_10625 = pop_1 & pop_valid & _GEN_10586; // @[lut_35.scala 3649:46 lut_35.scala 5097:40]
  wire  _GEN_10626 = pop_1 & pop_valid & _GEN_10587; // @[lut_35.scala 3649:46 lut_35.scala 5098:40]
  wire  _GEN_10627 = pop_1 & pop_valid & _GEN_10588; // @[lut_35.scala 3649:46 lut_35.scala 5099:40]
  wire  _GEN_10628 = pop_1 & pop_valid & _GEN_10589; // @[lut_35.scala 3649:46 lut_35.scala 5100:41]
  wire  _GEN_10629 = pop_1 & pop_valid & _GEN_10590; // @[lut_35.scala 3649:46 lut_35.scala 5101:41]
  wire  _GEN_10630 = pop_1 & pop_valid & _GEN_10591; // @[lut_35.scala 3649:46 lut_35.scala 5102:41]
  wire  _GEN_10631 = pop_1 & pop_valid & _GEN_10592; // @[lut_35.scala 3649:46 lut_35.scala 5103:41]
  wire  _GEN_10632 = pop_1 & pop_valid & _GEN_10593; // @[lut_35.scala 3649:46 lut_35.scala 5104:41]
  wire  _GEN_10633 = pop_1 & pop_valid & _GEN_10594; // @[lut_35.scala 3649:46 lut_35.scala 5105:41]
  wire  _GEN_10634 = pop_1 & pop_valid & _GEN_10595; // @[lut_35.scala 3649:46 lut_35.scala 5106:41]
  wire  _GEN_10635 = pop_1 & pop_valid & _GEN_10596; // @[lut_35.scala 3649:46 lut_35.scala 5107:41]
  wire  _GEN_10636 = pop_1 & pop_valid & _GEN_10597; // @[lut_35.scala 3649:46 lut_35.scala 5108:41]
  wire  _GEN_10637 = pop_1 & pop_valid & _GEN_10598; // @[lut_35.scala 3649:46 lut_35.scala 5109:41]
  wire  _GEN_10638 = pop_1 & pop_valid & _GEN_10599; // @[lut_35.scala 3649:46 lut_35.scala 5110:41]
  wire  _GEN_10639 = pop_1 & pop_valid & _GEN_10600; // @[lut_35.scala 3649:46 lut_35.scala 5111:41]
  wire  _GEN_10640 = pop_1 & pop_valid & _GEN_10601; // @[lut_35.scala 3649:46 lut_35.scala 5112:41]
  wire  _GEN_10641 = pop_1 & pop_valid & _GEN_10602; // @[lut_35.scala 3649:46 lut_35.scala 5113:41]
  wire  _GEN_10642 = pop_1 & pop_valid & _GEN_10603; // @[lut_35.scala 3649:46 lut_35.scala 5114:41]
  wire  _GEN_10643 = pop_1 & pop_valid & _GEN_10604; // @[lut_35.scala 3649:46 lut_35.scala 5115:41]
  wire  _GEN_10644 = pop_1 & pop_valid & _GEN_10605; // @[lut_35.scala 3649:46 lut_35.scala 5116:41]
  wire  _GEN_10645 = pop_1 & pop_valid & _GEN_10606; // @[lut_35.scala 3649:46 lut_35.scala 5117:41]
  wire  _GEN_10646 = pop_1 & pop_valid & _GEN_10607; // @[lut_35.scala 3649:46 lut_35.scala 5118:41]
  wire  _GEN_10647 = pop_1 & pop_valid & _GEN_10608; // @[lut_35.scala 3649:46 lut_35.scala 5119:41]
  wire  _GEN_10648 = pop_1 & pop_valid & _GEN_10609; // @[lut_35.scala 3649:46 lut_35.scala 5120:41]
  wire  _GEN_10649 = pop_1 & pop_valid & _GEN_10610; // @[lut_35.scala 3649:46 lut_35.scala 5121:41]
  wire  _GEN_10650 = pop_1 & pop_valid & _GEN_10611; // @[lut_35.scala 3649:46 lut_35.scala 5122:41]
  wire  _GEN_10651 = pop_1 & pop_valid & _GEN_10612; // @[lut_35.scala 3649:46 lut_35.scala 5123:41]
  wire  _GEN_10652 = pop_1 & pop_valid & _GEN_10613; // @[lut_35.scala 3649:46 lut_35.scala 5124:41]
  wire  _GEN_10653 = pop_1 & pop_valid & _GEN_10614; // @[lut_35.scala 3649:46 lut_35.scala 5125:37]
  reg  clear_1; // @[lut_35.scala 5175:38]
  reg [31:0] read_stack0_clear; // @[lut_35.scala 5176:40]
  reg [31:0] read_stack1_clear; // @[lut_35.scala 5177:40]
  reg [31:0] read_stack3_clear; // @[lut_35.scala 5179:40]
  reg [31:0] read_stack4_clear; // @[lut_35.scala 5180:40]
  reg [31:0] read_stack5_clear; // @[lut_35.scala 5181:40]
  reg [31:0] read_stack6_clear; // @[lut_35.scala 5182:40]
  reg [31:0] read_stack7_clear; // @[lut_35.scala 5183:40]
  reg [31:0] read_stack8_clear; // @[lut_35.scala 5184:40]
  reg [31:0] read_stack9_clear; // @[lut_35.scala 5185:40]
  reg [31:0] read_stack10_clear; // @[lut_35.scala 5186:41]
  reg [31:0] read_stack11_clear; // @[lut_35.scala 5187:41]
  reg [31:0] read_stack12_clear; // @[lut_35.scala 5188:41]
  reg [31:0] read_stack13_clear; // @[lut_35.scala 5189:41]
  reg [31:0] read_stack14_clear; // @[lut_35.scala 5190:41]
  reg [31:0] read_stack15_clear; // @[lut_35.scala 5191:41]
  reg [31:0] read_stack16_clear; // @[lut_35.scala 5192:41]
  reg [31:0] read_stack17_clear; // @[lut_35.scala 5193:41]
  reg [31:0] read_stack18_clear; // @[lut_35.scala 5194:41]
  reg [31:0] read_stack19_clear; // @[lut_35.scala 5195:41]
  reg [31:0] read_stack20_clear; // @[lut_35.scala 5196:41]
  reg [31:0] read_stack21_clear; // @[lut_35.scala 5197:41]
  reg [31:0] read_stack22_clear; // @[lut_35.scala 5198:41]
  reg [31:0] read_stack23_clear; // @[lut_35.scala 5199:41]
  reg [31:0] read_stack24_clear; // @[lut_35.scala 5200:41]
  reg [31:0] read_stack25_clear; // @[lut_35.scala 5201:41]
  reg [31:0] read_stack26_clear; // @[lut_35.scala 5202:41]
  reg [31:0] read_stack27_clear; // @[lut_35.scala 5203:41]
  reg [31:0] read_stack28_clear; // @[lut_35.scala 5204:41]
  reg [31:0] read_stack29_clear; // @[lut_35.scala 5205:41]
  reg [31:0] read_stack30_clear; // @[lut_35.scala 5206:41]
  reg [31:0] read_stack31_clear; // @[lut_35.scala 5207:41]
  reg [31:0] read_stack32_clear; // @[lut_35.scala 5208:41]
  reg [31:0] read_stack33_clear; // @[lut_35.scala 5209:41]
  reg [31:0] read_stack34_clear; // @[lut_35.scala 5210:41]
  reg [31:0] clear_ray_id; // @[lut_35.scala 5212:39]
  reg  clear_valid; // @[lut_35.scala 5213:38]
  reg  clear_0_1; // @[lut_35.scala 5216:48]
  reg  clear_1_1; // @[lut_35.scala 5217:48]
  reg  clear_2_1; // @[lut_35.scala 5218:48]
  reg  clear_3_1; // @[lut_35.scala 5219:48]
  reg  clear_4_1; // @[lut_35.scala 5220:48]
  reg  clear_5_1; // @[lut_35.scala 5221:48]
  reg  clear_6_1; // @[lut_35.scala 5222:48]
  reg  clear_7_1; // @[lut_35.scala 5223:48]
  reg  clear_8_1; // @[lut_35.scala 5224:48]
  reg  clear_9_1; // @[lut_35.scala 5225:48]
  reg  clear_10_1; // @[lut_35.scala 5226:49]
  reg  clear_11_1; // @[lut_35.scala 5227:49]
  reg  clear_12_1; // @[lut_35.scala 5228:49]
  reg  clear_13_1; // @[lut_35.scala 5229:49]
  reg  clear_14_1; // @[lut_35.scala 5230:49]
  reg  clear_15_1; // @[lut_35.scala 5231:49]
  reg  clear_16_1; // @[lut_35.scala 5232:49]
  reg  clear_17_1; // @[lut_35.scala 5233:49]
  reg  clear_18_1; // @[lut_35.scala 5234:49]
  reg  clear_19_1; // @[lut_35.scala 5235:49]
  reg  clear_20_1; // @[lut_35.scala 5236:49]
  reg  clear_21_1; // @[lut_35.scala 5237:49]
  reg  clear_22_1; // @[lut_35.scala 5238:49]
  reg  clear_23_1; // @[lut_35.scala 5239:49]
  reg  clear_24_1; // @[lut_35.scala 5240:49]
  reg  clear_25_1; // @[lut_35.scala 5241:49]
  reg  clear_26_1; // @[lut_35.scala 5242:49]
  reg  clear_27_1; // @[lut_35.scala 5243:49]
  reg  clear_28_1; // @[lut_35.scala 5244:49]
  reg  clear_29_1; // @[lut_35.scala 5245:49]
  reg  clear_30_1; // @[lut_35.scala 5246:49]
  reg  clear_31_1; // @[lut_35.scala 5247:49]
  reg  clear_32_1; // @[lut_35.scala 5248:49]
  reg  clear_33_1; // @[lut_35.scala 5249:49]
  reg  clear_34_1; // @[lut_35.scala 5250:49]
  wire  _T_790 = read_stack0_clear == clear_ray_id & clear_valid; // @[lut_35.scala 5307:49]
  wire  _T_793 = read_stack1_clear == clear_ray_id & clear_valid; // @[lut_35.scala 5345:59]
  wire  _T_796 = read_stack3_clear == clear_ray_id & clear_valid; // @[lut_35.scala 5383:59]
  wire  _T_802 = read_stack4_clear == clear_ray_id & clear_valid; // @[lut_35.scala 5459:59]
  wire  _T_805 = read_stack5_clear == clear_ray_id & clear_valid; // @[lut_35.scala 5497:59]
  wire  _T_808 = read_stack6_clear == clear_ray_id & clear_valid; // @[lut_35.scala 5535:59]
  wire  _T_811 = read_stack7_clear == clear_ray_id & clear_valid; // @[lut_35.scala 5573:59]
  wire  _T_814 = read_stack8_clear == clear_ray_id & clear_valid; // @[lut_35.scala 5611:59]
  wire  _T_817 = read_stack9_clear == clear_ray_id & clear_valid; // @[lut_35.scala 5649:59]
  wire  _T_820 = read_stack10_clear == clear_ray_id & clear_valid; // @[lut_35.scala 5687:60]
  wire  _T_823 = read_stack11_clear == clear_ray_id & clear_valid; // @[lut_35.scala 5725:60]
  wire  _T_826 = read_stack12_clear == clear_ray_id & clear_valid; // @[lut_35.scala 5763:60]
  wire  _T_829 = read_stack13_clear == clear_ray_id & clear_valid; // @[lut_35.scala 5801:60]
  wire  _T_832 = read_stack14_clear == clear_ray_id & clear_valid; // @[lut_35.scala 5839:60]
  wire  _T_835 = read_stack15_clear == clear_ray_id & clear_valid; // @[lut_35.scala 5877:60]
  wire  _T_838 = read_stack16_clear == clear_ray_id & clear_valid; // @[lut_35.scala 5915:60]
  wire  _T_841 = read_stack17_clear == clear_ray_id & clear_valid; // @[lut_35.scala 5953:60]
  wire  _T_844 = read_stack18_clear == clear_ray_id & clear_valid; // @[lut_35.scala 5991:60]
  wire  _T_847 = read_stack19_clear == clear_ray_id & clear_valid; // @[lut_35.scala 6029:60]
  wire  _T_850 = read_stack20_clear == clear_ray_id & clear_valid; // @[lut_35.scala 6067:60]
  wire  _T_853 = read_stack21_clear == clear_ray_id & clear_valid; // @[lut_35.scala 6105:60]
  wire  _T_856 = read_stack22_clear == clear_ray_id & clear_valid; // @[lut_35.scala 6143:60]
  wire  _T_859 = read_stack23_clear == clear_ray_id & clear_valid; // @[lut_35.scala 6181:60]
  wire  _T_862 = read_stack24_clear == clear_ray_id & clear_valid; // @[lut_35.scala 6219:60]
  wire  _T_865 = read_stack25_clear == clear_ray_id & clear_valid; // @[lut_35.scala 6257:60]
  wire  _T_868 = read_stack26_clear == clear_ray_id & clear_valid; // @[lut_35.scala 6295:60]
  wire  _T_871 = read_stack27_clear == clear_ray_id & clear_valid; // @[lut_35.scala 6333:60]
  wire  _T_874 = read_stack28_clear == clear_ray_id & clear_valid; // @[lut_35.scala 6371:60]
  wire  _T_877 = read_stack29_clear == clear_ray_id & clear_valid; // @[lut_35.scala 6409:60]
  wire  _T_880 = read_stack30_clear == clear_ray_id & clear_valid; // @[lut_35.scala 6447:60]
  wire  _T_883 = read_stack31_clear == clear_ray_id & clear_valid; // @[lut_35.scala 6485:60]
  wire  _T_886 = read_stack32_clear == clear_ray_id & clear_valid; // @[lut_35.scala 6523:60]
  wire  _T_889 = read_stack33_clear == clear_ray_id & clear_valid; // @[lut_35.scala 6561:60]
  wire  _T_892 = read_stack34_clear == clear_ray_id & clear_valid; // @[lut_35.scala 6599:60]
  wire  _GEN_10664 = read_stack33_clear == clear_ray_id & clear_valid ? 1'h0 : _T_892; // @[lut_35.scala 6561:84 lut_35.scala 6596:47]
  wire  _GEN_10669 = read_stack32_clear == clear_ray_id & clear_valid ? 1'h0 : _T_889; // @[lut_35.scala 6523:84 lut_35.scala 6557:47]
  wire  _GEN_10670 = read_stack32_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10664; // @[lut_35.scala 6523:84 lut_35.scala 6558:47]
  wire  _GEN_10675 = read_stack31_clear == clear_ray_id & clear_valid ? 1'h0 : _T_886; // @[lut_35.scala 6485:84 lut_35.scala 6518:47]
  wire  _GEN_10676 = read_stack31_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10669; // @[lut_35.scala 6485:84 lut_35.scala 6519:47]
  wire  _GEN_10677 = read_stack31_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10670; // @[lut_35.scala 6485:84 lut_35.scala 6520:47]
  wire  _GEN_10682 = read_stack30_clear == clear_ray_id & clear_valid ? 1'h0 : _T_883; // @[lut_35.scala 6447:84 lut_35.scala 6479:47]
  wire  _GEN_10683 = read_stack30_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10675; // @[lut_35.scala 6447:84 lut_35.scala 6480:47]
  wire  _GEN_10684 = read_stack30_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10676; // @[lut_35.scala 6447:84 lut_35.scala 6481:47]
  wire  _GEN_10685 = read_stack30_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10677; // @[lut_35.scala 6447:84 lut_35.scala 6482:47]
  wire  _GEN_10690 = read_stack29_clear == clear_ray_id & clear_valid ? 1'h0 : _T_880; // @[lut_35.scala 6409:84 lut_35.scala 6440:47]
  wire  _GEN_10691 = read_stack29_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10682; // @[lut_35.scala 6409:84 lut_35.scala 6441:47]
  wire  _GEN_10692 = read_stack29_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10683; // @[lut_35.scala 6409:84 lut_35.scala 6442:47]
  wire  _GEN_10693 = read_stack29_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10684; // @[lut_35.scala 6409:84 lut_35.scala 6443:47]
  wire  _GEN_10694 = read_stack29_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10685; // @[lut_35.scala 6409:84 lut_35.scala 6444:47]
  wire  _GEN_10699 = read_stack28_clear == clear_ray_id & clear_valid ? 1'h0 : _T_877; // @[lut_35.scala 6371:84 lut_35.scala 6401:47]
  wire  _GEN_10700 = read_stack28_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10690; // @[lut_35.scala 6371:84 lut_35.scala 6402:47]
  wire  _GEN_10701 = read_stack28_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10691; // @[lut_35.scala 6371:84 lut_35.scala 6403:47]
  wire  _GEN_10702 = read_stack28_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10692; // @[lut_35.scala 6371:84 lut_35.scala 6404:47]
  wire  _GEN_10703 = read_stack28_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10693; // @[lut_35.scala 6371:84 lut_35.scala 6405:47]
  wire  _GEN_10704 = read_stack28_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10694; // @[lut_35.scala 6371:84 lut_35.scala 6406:47]
  wire  _GEN_10709 = read_stack27_clear == clear_ray_id & clear_valid ? 1'h0 : _T_874; // @[lut_35.scala 6333:84 lut_35.scala 6362:47]
  wire  _GEN_10710 = read_stack27_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10699; // @[lut_35.scala 6333:84 lut_35.scala 6363:47]
  wire  _GEN_10711 = read_stack27_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10700; // @[lut_35.scala 6333:84 lut_35.scala 6364:47]
  wire  _GEN_10712 = read_stack27_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10701; // @[lut_35.scala 6333:84 lut_35.scala 6365:47]
  wire  _GEN_10713 = read_stack27_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10702; // @[lut_35.scala 6333:84 lut_35.scala 6366:47]
  wire  _GEN_10714 = read_stack27_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10703; // @[lut_35.scala 6333:84 lut_35.scala 6367:47]
  wire  _GEN_10715 = read_stack27_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10704; // @[lut_35.scala 6333:84 lut_35.scala 6368:47]
  wire  _GEN_10720 = read_stack26_clear == clear_ray_id & clear_valid ? 1'h0 : _T_871; // @[lut_35.scala 6295:84 lut_35.scala 6323:47]
  wire  _GEN_10721 = read_stack26_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10709; // @[lut_35.scala 6295:84 lut_35.scala 6324:47]
  wire  _GEN_10722 = read_stack26_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10710; // @[lut_35.scala 6295:84 lut_35.scala 6325:47]
  wire  _GEN_10723 = read_stack26_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10711; // @[lut_35.scala 6295:84 lut_35.scala 6326:47]
  wire  _GEN_10724 = read_stack26_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10712; // @[lut_35.scala 6295:84 lut_35.scala 6327:47]
  wire  _GEN_10725 = read_stack26_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10713; // @[lut_35.scala 6295:84 lut_35.scala 6328:47]
  wire  _GEN_10726 = read_stack26_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10714; // @[lut_35.scala 6295:84 lut_35.scala 6329:47]
  wire  _GEN_10727 = read_stack26_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10715; // @[lut_35.scala 6295:84 lut_35.scala 6330:47]
  wire  _GEN_10732 = read_stack25_clear == clear_ray_id & clear_valid ? 1'h0 : _T_868; // @[lut_35.scala 6257:84 lut_35.scala 6284:47]
  wire  _GEN_10733 = read_stack25_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10720; // @[lut_35.scala 6257:84 lut_35.scala 6285:47]
  wire  _GEN_10734 = read_stack25_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10721; // @[lut_35.scala 6257:84 lut_35.scala 6286:47]
  wire  _GEN_10735 = read_stack25_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10722; // @[lut_35.scala 6257:84 lut_35.scala 6287:47]
  wire  _GEN_10736 = read_stack25_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10723; // @[lut_35.scala 6257:84 lut_35.scala 6288:47]
  wire  _GEN_10737 = read_stack25_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10724; // @[lut_35.scala 6257:84 lut_35.scala 6289:47]
  wire  _GEN_10738 = read_stack25_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10725; // @[lut_35.scala 6257:84 lut_35.scala 6290:47]
  wire  _GEN_10739 = read_stack25_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10726; // @[lut_35.scala 6257:84 lut_35.scala 6291:47]
  wire  _GEN_10740 = read_stack25_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10727; // @[lut_35.scala 6257:84 lut_35.scala 6292:47]
  wire  _GEN_10745 = read_stack24_clear == clear_ray_id & clear_valid ? 1'h0 : _T_865; // @[lut_35.scala 6219:84 lut_35.scala 6245:47]
  wire  _GEN_10746 = read_stack24_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10732; // @[lut_35.scala 6219:84 lut_35.scala 6246:47]
  wire  _GEN_10747 = read_stack24_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10733; // @[lut_35.scala 6219:84 lut_35.scala 6247:47]
  wire  _GEN_10748 = read_stack24_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10734; // @[lut_35.scala 6219:84 lut_35.scala 6248:47]
  wire  _GEN_10749 = read_stack24_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10735; // @[lut_35.scala 6219:84 lut_35.scala 6249:47]
  wire  _GEN_10750 = read_stack24_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10736; // @[lut_35.scala 6219:84 lut_35.scala 6250:47]
  wire  _GEN_10751 = read_stack24_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10737; // @[lut_35.scala 6219:84 lut_35.scala 6251:47]
  wire  _GEN_10752 = read_stack24_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10738; // @[lut_35.scala 6219:84 lut_35.scala 6252:47]
  wire  _GEN_10753 = read_stack24_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10739; // @[lut_35.scala 6219:84 lut_35.scala 6253:47]
  wire  _GEN_10754 = read_stack24_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10740; // @[lut_35.scala 6219:84 lut_35.scala 6254:47]
  wire  _GEN_10759 = read_stack23_clear == clear_ray_id & clear_valid ? 1'h0 : _T_862; // @[lut_35.scala 6181:84 lut_35.scala 6206:47]
  wire  _GEN_10760 = read_stack23_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10745; // @[lut_35.scala 6181:84 lut_35.scala 6207:47]
  wire  _GEN_10761 = read_stack23_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10746; // @[lut_35.scala 6181:84 lut_35.scala 6208:47]
  wire  _GEN_10762 = read_stack23_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10747; // @[lut_35.scala 6181:84 lut_35.scala 6209:47]
  wire  _GEN_10763 = read_stack23_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10748; // @[lut_35.scala 6181:84 lut_35.scala 6210:47]
  wire  _GEN_10764 = read_stack23_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10749; // @[lut_35.scala 6181:84 lut_35.scala 6211:47]
  wire  _GEN_10765 = read_stack23_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10750; // @[lut_35.scala 6181:84 lut_35.scala 6212:47]
  wire  _GEN_10766 = read_stack23_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10751; // @[lut_35.scala 6181:84 lut_35.scala 6213:47]
  wire  _GEN_10767 = read_stack23_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10752; // @[lut_35.scala 6181:84 lut_35.scala 6214:47]
  wire  _GEN_10768 = read_stack23_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10753; // @[lut_35.scala 6181:84 lut_35.scala 6215:47]
  wire  _GEN_10769 = read_stack23_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10754; // @[lut_35.scala 6181:84 lut_35.scala 6216:47]
  wire  _GEN_10774 = read_stack22_clear == clear_ray_id & clear_valid ? 1'h0 : _T_859; // @[lut_35.scala 6143:84 lut_35.scala 6167:47]
  wire  _GEN_10775 = read_stack22_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10759; // @[lut_35.scala 6143:84 lut_35.scala 6168:47]
  wire  _GEN_10776 = read_stack22_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10760; // @[lut_35.scala 6143:84 lut_35.scala 6169:47]
  wire  _GEN_10777 = read_stack22_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10761; // @[lut_35.scala 6143:84 lut_35.scala 6170:47]
  wire  _GEN_10778 = read_stack22_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10762; // @[lut_35.scala 6143:84 lut_35.scala 6171:47]
  wire  _GEN_10779 = read_stack22_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10763; // @[lut_35.scala 6143:84 lut_35.scala 6172:47]
  wire  _GEN_10780 = read_stack22_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10764; // @[lut_35.scala 6143:84 lut_35.scala 6173:47]
  wire  _GEN_10781 = read_stack22_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10765; // @[lut_35.scala 6143:84 lut_35.scala 6174:47]
  wire  _GEN_10782 = read_stack22_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10766; // @[lut_35.scala 6143:84 lut_35.scala 6175:47]
  wire  _GEN_10783 = read_stack22_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10767; // @[lut_35.scala 6143:84 lut_35.scala 6176:47]
  wire  _GEN_10784 = read_stack22_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10768; // @[lut_35.scala 6143:84 lut_35.scala 6177:47]
  wire  _GEN_10785 = read_stack22_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10769; // @[lut_35.scala 6143:84 lut_35.scala 6178:47]
  wire  _GEN_10790 = read_stack21_clear == clear_ray_id & clear_valid ? 1'h0 : _T_856; // @[lut_35.scala 6105:84 lut_35.scala 6128:47]
  wire  _GEN_10791 = read_stack21_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10774; // @[lut_35.scala 6105:84 lut_35.scala 6129:47]
  wire  _GEN_10792 = read_stack21_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10775; // @[lut_35.scala 6105:84 lut_35.scala 6130:47]
  wire  _GEN_10793 = read_stack21_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10776; // @[lut_35.scala 6105:84 lut_35.scala 6131:47]
  wire  _GEN_10794 = read_stack21_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10777; // @[lut_35.scala 6105:84 lut_35.scala 6132:47]
  wire  _GEN_10795 = read_stack21_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10778; // @[lut_35.scala 6105:84 lut_35.scala 6133:47]
  wire  _GEN_10796 = read_stack21_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10779; // @[lut_35.scala 6105:84 lut_35.scala 6134:47]
  wire  _GEN_10797 = read_stack21_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10780; // @[lut_35.scala 6105:84 lut_35.scala 6135:47]
  wire  _GEN_10798 = read_stack21_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10781; // @[lut_35.scala 6105:84 lut_35.scala 6136:47]
  wire  _GEN_10799 = read_stack21_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10782; // @[lut_35.scala 6105:84 lut_35.scala 6137:47]
  wire  _GEN_10800 = read_stack21_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10783; // @[lut_35.scala 6105:84 lut_35.scala 6138:47]
  wire  _GEN_10801 = read_stack21_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10784; // @[lut_35.scala 6105:84 lut_35.scala 6139:47]
  wire  _GEN_10802 = read_stack21_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10785; // @[lut_35.scala 6105:84 lut_35.scala 6140:47]
  wire  _GEN_10807 = read_stack20_clear == clear_ray_id & clear_valid ? 1'h0 : _T_853; // @[lut_35.scala 6067:84 lut_35.scala 6089:47]
  wire  _GEN_10808 = read_stack20_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10790; // @[lut_35.scala 6067:84 lut_35.scala 6090:47]
  wire  _GEN_10809 = read_stack20_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10791; // @[lut_35.scala 6067:84 lut_35.scala 6091:47]
  wire  _GEN_10810 = read_stack20_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10792; // @[lut_35.scala 6067:84 lut_35.scala 6092:47]
  wire  _GEN_10811 = read_stack20_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10793; // @[lut_35.scala 6067:84 lut_35.scala 6093:47]
  wire  _GEN_10812 = read_stack20_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10794; // @[lut_35.scala 6067:84 lut_35.scala 6094:47]
  wire  _GEN_10813 = read_stack20_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10795; // @[lut_35.scala 6067:84 lut_35.scala 6095:47]
  wire  _GEN_10814 = read_stack20_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10796; // @[lut_35.scala 6067:84 lut_35.scala 6096:47]
  wire  _GEN_10815 = read_stack20_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10797; // @[lut_35.scala 6067:84 lut_35.scala 6097:47]
  wire  _GEN_10816 = read_stack20_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10798; // @[lut_35.scala 6067:84 lut_35.scala 6098:47]
  wire  _GEN_10817 = read_stack20_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10799; // @[lut_35.scala 6067:84 lut_35.scala 6099:47]
  wire  _GEN_10818 = read_stack20_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10800; // @[lut_35.scala 6067:84 lut_35.scala 6100:47]
  wire  _GEN_10819 = read_stack20_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10801; // @[lut_35.scala 6067:84 lut_35.scala 6101:47]
  wire  _GEN_10820 = read_stack20_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10802; // @[lut_35.scala 6067:84 lut_35.scala 6102:47]
  wire  _GEN_10825 = read_stack19_clear == clear_ray_id & clear_valid ? 1'h0 : _T_850; // @[lut_35.scala 6029:84 lut_35.scala 6050:47]
  wire  _GEN_10826 = read_stack19_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10807; // @[lut_35.scala 6029:84 lut_35.scala 6051:47]
  wire  _GEN_10827 = read_stack19_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10808; // @[lut_35.scala 6029:84 lut_35.scala 6052:47]
  wire  _GEN_10828 = read_stack19_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10809; // @[lut_35.scala 6029:84 lut_35.scala 6053:47]
  wire  _GEN_10829 = read_stack19_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10810; // @[lut_35.scala 6029:84 lut_35.scala 6054:47]
  wire  _GEN_10830 = read_stack19_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10811; // @[lut_35.scala 6029:84 lut_35.scala 6055:47]
  wire  _GEN_10831 = read_stack19_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10812; // @[lut_35.scala 6029:84 lut_35.scala 6056:47]
  wire  _GEN_10832 = read_stack19_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10813; // @[lut_35.scala 6029:84 lut_35.scala 6057:47]
  wire  _GEN_10833 = read_stack19_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10814; // @[lut_35.scala 6029:84 lut_35.scala 6058:47]
  wire  _GEN_10834 = read_stack19_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10815; // @[lut_35.scala 6029:84 lut_35.scala 6059:47]
  wire  _GEN_10835 = read_stack19_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10816; // @[lut_35.scala 6029:84 lut_35.scala 6060:47]
  wire  _GEN_10836 = read_stack19_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10817; // @[lut_35.scala 6029:84 lut_35.scala 6061:47]
  wire  _GEN_10837 = read_stack19_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10818; // @[lut_35.scala 6029:84 lut_35.scala 6062:47]
  wire  _GEN_10838 = read_stack19_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10819; // @[lut_35.scala 6029:84 lut_35.scala 6063:47]
  wire  _GEN_10839 = read_stack19_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10820; // @[lut_35.scala 6029:84 lut_35.scala 6064:47]
  wire  _GEN_10844 = read_stack18_clear == clear_ray_id & clear_valid ? 1'h0 : _T_847; // @[lut_35.scala 5991:84 lut_35.scala 6011:47]
  wire  _GEN_10845 = read_stack18_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10825; // @[lut_35.scala 5991:84 lut_35.scala 6012:47]
  wire  _GEN_10846 = read_stack18_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10826; // @[lut_35.scala 5991:84 lut_35.scala 6013:47]
  wire  _GEN_10847 = read_stack18_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10827; // @[lut_35.scala 5991:84 lut_35.scala 6014:47]
  wire  _GEN_10848 = read_stack18_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10828; // @[lut_35.scala 5991:84 lut_35.scala 6015:47]
  wire  _GEN_10849 = read_stack18_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10829; // @[lut_35.scala 5991:84 lut_35.scala 6016:47]
  wire  _GEN_10850 = read_stack18_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10830; // @[lut_35.scala 5991:84 lut_35.scala 6017:47]
  wire  _GEN_10851 = read_stack18_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10831; // @[lut_35.scala 5991:84 lut_35.scala 6018:47]
  wire  _GEN_10852 = read_stack18_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10832; // @[lut_35.scala 5991:84 lut_35.scala 6019:47]
  wire  _GEN_10853 = read_stack18_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10833; // @[lut_35.scala 5991:84 lut_35.scala 6020:47]
  wire  _GEN_10854 = read_stack18_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10834; // @[lut_35.scala 5991:84 lut_35.scala 6021:47]
  wire  _GEN_10855 = read_stack18_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10835; // @[lut_35.scala 5991:84 lut_35.scala 6022:47]
  wire  _GEN_10856 = read_stack18_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10836; // @[lut_35.scala 5991:84 lut_35.scala 6023:47]
  wire  _GEN_10857 = read_stack18_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10837; // @[lut_35.scala 5991:84 lut_35.scala 6024:47]
  wire  _GEN_10858 = read_stack18_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10838; // @[lut_35.scala 5991:84 lut_35.scala 6025:47]
  wire  _GEN_10859 = read_stack18_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10839; // @[lut_35.scala 5991:84 lut_35.scala 6026:47]
  wire  _GEN_10864 = read_stack17_clear == clear_ray_id & clear_valid ? 1'h0 : _T_844; // @[lut_35.scala 5953:84 lut_35.scala 5972:47]
  wire  _GEN_10865 = read_stack17_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10844; // @[lut_35.scala 5953:84 lut_35.scala 5973:47]
  wire  _GEN_10866 = read_stack17_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10845; // @[lut_35.scala 5953:84 lut_35.scala 5974:47]
  wire  _GEN_10867 = read_stack17_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10846; // @[lut_35.scala 5953:84 lut_35.scala 5975:47]
  wire  _GEN_10868 = read_stack17_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10847; // @[lut_35.scala 5953:84 lut_35.scala 5976:47]
  wire  _GEN_10869 = read_stack17_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10848; // @[lut_35.scala 5953:84 lut_35.scala 5977:47]
  wire  _GEN_10870 = read_stack17_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10849; // @[lut_35.scala 5953:84 lut_35.scala 5978:47]
  wire  _GEN_10871 = read_stack17_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10850; // @[lut_35.scala 5953:84 lut_35.scala 5979:47]
  wire  _GEN_10872 = read_stack17_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10851; // @[lut_35.scala 5953:84 lut_35.scala 5980:47]
  wire  _GEN_10873 = read_stack17_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10852; // @[lut_35.scala 5953:84 lut_35.scala 5981:47]
  wire  _GEN_10874 = read_stack17_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10853; // @[lut_35.scala 5953:84 lut_35.scala 5982:47]
  wire  _GEN_10875 = read_stack17_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10854; // @[lut_35.scala 5953:84 lut_35.scala 5983:47]
  wire  _GEN_10876 = read_stack17_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10855; // @[lut_35.scala 5953:84 lut_35.scala 5984:47]
  wire  _GEN_10877 = read_stack17_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10856; // @[lut_35.scala 5953:84 lut_35.scala 5985:47]
  wire  _GEN_10878 = read_stack17_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10857; // @[lut_35.scala 5953:84 lut_35.scala 5986:47]
  wire  _GEN_10879 = read_stack17_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10858; // @[lut_35.scala 5953:84 lut_35.scala 5987:47]
  wire  _GEN_10880 = read_stack17_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10859; // @[lut_35.scala 5953:84 lut_35.scala 5988:47]
  wire  _GEN_10885 = read_stack16_clear == clear_ray_id & clear_valid ? 1'h0 : _T_841; // @[lut_35.scala 5915:84 lut_35.scala 5933:47]
  wire  _GEN_10886 = read_stack16_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10864; // @[lut_35.scala 5915:84 lut_35.scala 5934:47]
  wire  _GEN_10887 = read_stack16_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10865; // @[lut_35.scala 5915:84 lut_35.scala 5935:47]
  wire  _GEN_10888 = read_stack16_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10866; // @[lut_35.scala 5915:84 lut_35.scala 5936:47]
  wire  _GEN_10889 = read_stack16_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10867; // @[lut_35.scala 5915:84 lut_35.scala 5937:47]
  wire  _GEN_10890 = read_stack16_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10868; // @[lut_35.scala 5915:84 lut_35.scala 5938:47]
  wire  _GEN_10891 = read_stack16_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10869; // @[lut_35.scala 5915:84 lut_35.scala 5939:47]
  wire  _GEN_10892 = read_stack16_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10870; // @[lut_35.scala 5915:84 lut_35.scala 5940:47]
  wire  _GEN_10893 = read_stack16_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10871; // @[lut_35.scala 5915:84 lut_35.scala 5941:47]
  wire  _GEN_10894 = read_stack16_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10872; // @[lut_35.scala 5915:84 lut_35.scala 5942:47]
  wire  _GEN_10895 = read_stack16_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10873; // @[lut_35.scala 5915:84 lut_35.scala 5943:47]
  wire  _GEN_10896 = read_stack16_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10874; // @[lut_35.scala 5915:84 lut_35.scala 5944:47]
  wire  _GEN_10897 = read_stack16_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10875; // @[lut_35.scala 5915:84 lut_35.scala 5945:47]
  wire  _GEN_10898 = read_stack16_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10876; // @[lut_35.scala 5915:84 lut_35.scala 5946:47]
  wire  _GEN_10899 = read_stack16_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10877; // @[lut_35.scala 5915:84 lut_35.scala 5947:47]
  wire  _GEN_10900 = read_stack16_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10878; // @[lut_35.scala 5915:84 lut_35.scala 5948:47]
  wire  _GEN_10901 = read_stack16_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10879; // @[lut_35.scala 5915:84 lut_35.scala 5949:47]
  wire  _GEN_10902 = read_stack16_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10880; // @[lut_35.scala 5915:84 lut_35.scala 5950:47]
  wire  _GEN_10907 = read_stack15_clear == clear_ray_id & clear_valid ? 1'h0 : _T_838; // @[lut_35.scala 5877:84 lut_35.scala 5894:47]
  wire  _GEN_10908 = read_stack15_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10885; // @[lut_35.scala 5877:84 lut_35.scala 5895:47]
  wire  _GEN_10909 = read_stack15_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10886; // @[lut_35.scala 5877:84 lut_35.scala 5896:47]
  wire  _GEN_10910 = read_stack15_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10887; // @[lut_35.scala 5877:84 lut_35.scala 5897:47]
  wire  _GEN_10911 = read_stack15_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10888; // @[lut_35.scala 5877:84 lut_35.scala 5898:47]
  wire  _GEN_10912 = read_stack15_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10889; // @[lut_35.scala 5877:84 lut_35.scala 5899:47]
  wire  _GEN_10913 = read_stack15_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10890; // @[lut_35.scala 5877:84 lut_35.scala 5900:47]
  wire  _GEN_10914 = read_stack15_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10891; // @[lut_35.scala 5877:84 lut_35.scala 5901:47]
  wire  _GEN_10915 = read_stack15_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10892; // @[lut_35.scala 5877:84 lut_35.scala 5902:47]
  wire  _GEN_10916 = read_stack15_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10893; // @[lut_35.scala 5877:84 lut_35.scala 5903:47]
  wire  _GEN_10917 = read_stack15_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10894; // @[lut_35.scala 5877:84 lut_35.scala 5904:47]
  wire  _GEN_10918 = read_stack15_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10895; // @[lut_35.scala 5877:84 lut_35.scala 5905:47]
  wire  _GEN_10919 = read_stack15_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10896; // @[lut_35.scala 5877:84 lut_35.scala 5906:47]
  wire  _GEN_10920 = read_stack15_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10897; // @[lut_35.scala 5877:84 lut_35.scala 5907:47]
  wire  _GEN_10921 = read_stack15_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10898; // @[lut_35.scala 5877:84 lut_35.scala 5908:47]
  wire  _GEN_10922 = read_stack15_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10899; // @[lut_35.scala 5877:84 lut_35.scala 5909:47]
  wire  _GEN_10923 = read_stack15_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10900; // @[lut_35.scala 5877:84 lut_35.scala 5910:47]
  wire  _GEN_10924 = read_stack15_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10901; // @[lut_35.scala 5877:84 lut_35.scala 5911:47]
  wire  _GEN_10925 = read_stack15_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10902; // @[lut_35.scala 5877:84 lut_35.scala 5912:47]
  wire  _GEN_10930 = read_stack14_clear == clear_ray_id & clear_valid ? 1'h0 : _T_835; // @[lut_35.scala 5839:84 lut_35.scala 5855:47]
  wire  _GEN_10931 = read_stack14_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10907; // @[lut_35.scala 5839:84 lut_35.scala 5856:47]
  wire  _GEN_10932 = read_stack14_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10908; // @[lut_35.scala 5839:84 lut_35.scala 5857:47]
  wire  _GEN_10933 = read_stack14_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10909; // @[lut_35.scala 5839:84 lut_35.scala 5858:47]
  wire  _GEN_10934 = read_stack14_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10910; // @[lut_35.scala 5839:84 lut_35.scala 5859:47]
  wire  _GEN_10935 = read_stack14_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10911; // @[lut_35.scala 5839:84 lut_35.scala 5860:47]
  wire  _GEN_10936 = read_stack14_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10912; // @[lut_35.scala 5839:84 lut_35.scala 5861:47]
  wire  _GEN_10937 = read_stack14_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10913; // @[lut_35.scala 5839:84 lut_35.scala 5862:47]
  wire  _GEN_10938 = read_stack14_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10914; // @[lut_35.scala 5839:84 lut_35.scala 5863:47]
  wire  _GEN_10939 = read_stack14_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10915; // @[lut_35.scala 5839:84 lut_35.scala 5864:47]
  wire  _GEN_10940 = read_stack14_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10916; // @[lut_35.scala 5839:84 lut_35.scala 5865:47]
  wire  _GEN_10941 = read_stack14_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10917; // @[lut_35.scala 5839:84 lut_35.scala 5866:47]
  wire  _GEN_10942 = read_stack14_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10918; // @[lut_35.scala 5839:84 lut_35.scala 5867:47]
  wire  _GEN_10943 = read_stack14_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10919; // @[lut_35.scala 5839:84 lut_35.scala 5868:47]
  wire  _GEN_10944 = read_stack14_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10920; // @[lut_35.scala 5839:84 lut_35.scala 5869:47]
  wire  _GEN_10945 = read_stack14_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10921; // @[lut_35.scala 5839:84 lut_35.scala 5870:47]
  wire  _GEN_10946 = read_stack14_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10922; // @[lut_35.scala 5839:84 lut_35.scala 5871:47]
  wire  _GEN_10947 = read_stack14_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10923; // @[lut_35.scala 5839:84 lut_35.scala 5872:47]
  wire  _GEN_10948 = read_stack14_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10924; // @[lut_35.scala 5839:84 lut_35.scala 5873:47]
  wire  _GEN_10949 = read_stack14_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10925; // @[lut_35.scala 5839:84 lut_35.scala 5874:47]
  wire  _GEN_10954 = read_stack13_clear == clear_ray_id & clear_valid ? 1'h0 : _T_832; // @[lut_35.scala 5801:84 lut_35.scala 5816:47]
  wire  _GEN_10955 = read_stack13_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10930; // @[lut_35.scala 5801:84 lut_35.scala 5817:47]
  wire  _GEN_10956 = read_stack13_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10931; // @[lut_35.scala 5801:84 lut_35.scala 5818:47]
  wire  _GEN_10957 = read_stack13_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10932; // @[lut_35.scala 5801:84 lut_35.scala 5819:47]
  wire  _GEN_10958 = read_stack13_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10933; // @[lut_35.scala 5801:84 lut_35.scala 5820:47]
  wire  _GEN_10959 = read_stack13_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10934; // @[lut_35.scala 5801:84 lut_35.scala 5821:47]
  wire  _GEN_10960 = read_stack13_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10935; // @[lut_35.scala 5801:84 lut_35.scala 5822:47]
  wire  _GEN_10961 = read_stack13_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10936; // @[lut_35.scala 5801:84 lut_35.scala 5823:47]
  wire  _GEN_10962 = read_stack13_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10937; // @[lut_35.scala 5801:84 lut_35.scala 5824:47]
  wire  _GEN_10963 = read_stack13_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10938; // @[lut_35.scala 5801:84 lut_35.scala 5825:47]
  wire  _GEN_10964 = read_stack13_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10939; // @[lut_35.scala 5801:84 lut_35.scala 5826:47]
  wire  _GEN_10965 = read_stack13_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10940; // @[lut_35.scala 5801:84 lut_35.scala 5827:47]
  wire  _GEN_10966 = read_stack13_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10941; // @[lut_35.scala 5801:84 lut_35.scala 5828:47]
  wire  _GEN_10967 = read_stack13_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10942; // @[lut_35.scala 5801:84 lut_35.scala 5829:47]
  wire  _GEN_10968 = read_stack13_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10943; // @[lut_35.scala 5801:84 lut_35.scala 5830:47]
  wire  _GEN_10969 = read_stack13_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10944; // @[lut_35.scala 5801:84 lut_35.scala 5831:47]
  wire  _GEN_10970 = read_stack13_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10945; // @[lut_35.scala 5801:84 lut_35.scala 5832:47]
  wire  _GEN_10971 = read_stack13_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10946; // @[lut_35.scala 5801:84 lut_35.scala 5833:47]
  wire  _GEN_10972 = read_stack13_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10947; // @[lut_35.scala 5801:84 lut_35.scala 5834:47]
  wire  _GEN_10973 = read_stack13_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10948; // @[lut_35.scala 5801:84 lut_35.scala 5835:47]
  wire  _GEN_10974 = read_stack13_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10949; // @[lut_35.scala 5801:84 lut_35.scala 5836:47]
  wire  _GEN_10979 = read_stack12_clear == clear_ray_id & clear_valid ? 1'h0 : _T_829; // @[lut_35.scala 5763:84 lut_35.scala 5777:47]
  wire  _GEN_10980 = read_stack12_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10954; // @[lut_35.scala 5763:84 lut_35.scala 5778:47]
  wire  _GEN_10981 = read_stack12_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10955; // @[lut_35.scala 5763:84 lut_35.scala 5779:47]
  wire  _GEN_10982 = read_stack12_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10956; // @[lut_35.scala 5763:84 lut_35.scala 5780:47]
  wire  _GEN_10983 = read_stack12_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10957; // @[lut_35.scala 5763:84 lut_35.scala 5781:47]
  wire  _GEN_10984 = read_stack12_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10958; // @[lut_35.scala 5763:84 lut_35.scala 5782:47]
  wire  _GEN_10985 = read_stack12_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10959; // @[lut_35.scala 5763:84 lut_35.scala 5783:47]
  wire  _GEN_10986 = read_stack12_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10960; // @[lut_35.scala 5763:84 lut_35.scala 5784:47]
  wire  _GEN_10987 = read_stack12_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10961; // @[lut_35.scala 5763:84 lut_35.scala 5785:47]
  wire  _GEN_10988 = read_stack12_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10962; // @[lut_35.scala 5763:84 lut_35.scala 5786:47]
  wire  _GEN_10989 = read_stack12_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10963; // @[lut_35.scala 5763:84 lut_35.scala 5787:47]
  wire  _GEN_10990 = read_stack12_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10964; // @[lut_35.scala 5763:84 lut_35.scala 5788:47]
  wire  _GEN_10991 = read_stack12_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10965; // @[lut_35.scala 5763:84 lut_35.scala 5789:47]
  wire  _GEN_10992 = read_stack12_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10966; // @[lut_35.scala 5763:84 lut_35.scala 5790:47]
  wire  _GEN_10993 = read_stack12_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10967; // @[lut_35.scala 5763:84 lut_35.scala 5791:47]
  wire  _GEN_10994 = read_stack12_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10968; // @[lut_35.scala 5763:84 lut_35.scala 5792:47]
  wire  _GEN_10995 = read_stack12_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10969; // @[lut_35.scala 5763:84 lut_35.scala 5793:47]
  wire  _GEN_10996 = read_stack12_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10970; // @[lut_35.scala 5763:84 lut_35.scala 5794:47]
  wire  _GEN_10997 = read_stack12_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10971; // @[lut_35.scala 5763:84 lut_35.scala 5795:47]
  wire  _GEN_10998 = read_stack12_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10972; // @[lut_35.scala 5763:84 lut_35.scala 5796:47]
  wire  _GEN_10999 = read_stack12_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10973; // @[lut_35.scala 5763:84 lut_35.scala 5797:47]
  wire  _GEN_11000 = read_stack12_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10974; // @[lut_35.scala 5763:84 lut_35.scala 5798:47]
  wire  _GEN_11005 = read_stack11_clear == clear_ray_id & clear_valid ? 1'h0 : _T_826; // @[lut_35.scala 5725:84 lut_35.scala 5738:47]
  wire  _GEN_11006 = read_stack11_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10979; // @[lut_35.scala 5725:84 lut_35.scala 5739:47]
  wire  _GEN_11007 = read_stack11_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10980; // @[lut_35.scala 5725:84 lut_35.scala 5740:47]
  wire  _GEN_11008 = read_stack11_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10981; // @[lut_35.scala 5725:84 lut_35.scala 5741:47]
  wire  _GEN_11009 = read_stack11_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10982; // @[lut_35.scala 5725:84 lut_35.scala 5742:47]
  wire  _GEN_11010 = read_stack11_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10983; // @[lut_35.scala 5725:84 lut_35.scala 5743:47]
  wire  _GEN_11011 = read_stack11_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10984; // @[lut_35.scala 5725:84 lut_35.scala 5744:47]
  wire  _GEN_11012 = read_stack11_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10985; // @[lut_35.scala 5725:84 lut_35.scala 5745:47]
  wire  _GEN_11013 = read_stack11_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10986; // @[lut_35.scala 5725:84 lut_35.scala 5746:47]
  wire  _GEN_11014 = read_stack11_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10987; // @[lut_35.scala 5725:84 lut_35.scala 5747:47]
  wire  _GEN_11015 = read_stack11_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10988; // @[lut_35.scala 5725:84 lut_35.scala 5748:47]
  wire  _GEN_11016 = read_stack11_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10989; // @[lut_35.scala 5725:84 lut_35.scala 5749:47]
  wire  _GEN_11017 = read_stack11_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10990; // @[lut_35.scala 5725:84 lut_35.scala 5750:47]
  wire  _GEN_11018 = read_stack11_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10991; // @[lut_35.scala 5725:84 lut_35.scala 5751:47]
  wire  _GEN_11019 = read_stack11_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10992; // @[lut_35.scala 5725:84 lut_35.scala 5752:47]
  wire  _GEN_11020 = read_stack11_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10993; // @[lut_35.scala 5725:84 lut_35.scala 5753:47]
  wire  _GEN_11021 = read_stack11_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10994; // @[lut_35.scala 5725:84 lut_35.scala 5754:47]
  wire  _GEN_11022 = read_stack11_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10995; // @[lut_35.scala 5725:84 lut_35.scala 5755:47]
  wire  _GEN_11023 = read_stack11_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10996; // @[lut_35.scala 5725:84 lut_35.scala 5756:47]
  wire  _GEN_11024 = read_stack11_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10997; // @[lut_35.scala 5725:84 lut_35.scala 5757:47]
  wire  _GEN_11025 = read_stack11_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10998; // @[lut_35.scala 5725:84 lut_35.scala 5758:47]
  wire  _GEN_11026 = read_stack11_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_10999; // @[lut_35.scala 5725:84 lut_35.scala 5759:47]
  wire  _GEN_11027 = read_stack11_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11000; // @[lut_35.scala 5725:84 lut_35.scala 5760:47]
  wire  _GEN_11032 = read_stack10_clear == clear_ray_id & clear_valid ? 1'h0 : _T_823; // @[lut_35.scala 5687:84 lut_35.scala 5699:47]
  wire  _GEN_11033 = read_stack10_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11005; // @[lut_35.scala 5687:84 lut_35.scala 5700:47]
  wire  _GEN_11034 = read_stack10_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11006; // @[lut_35.scala 5687:84 lut_35.scala 5701:47]
  wire  _GEN_11035 = read_stack10_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11007; // @[lut_35.scala 5687:84 lut_35.scala 5702:47]
  wire  _GEN_11036 = read_stack10_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11008; // @[lut_35.scala 5687:84 lut_35.scala 5703:47]
  wire  _GEN_11037 = read_stack10_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11009; // @[lut_35.scala 5687:84 lut_35.scala 5704:47]
  wire  _GEN_11038 = read_stack10_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11010; // @[lut_35.scala 5687:84 lut_35.scala 5705:47]
  wire  _GEN_11039 = read_stack10_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11011; // @[lut_35.scala 5687:84 lut_35.scala 5706:47]
  wire  _GEN_11040 = read_stack10_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11012; // @[lut_35.scala 5687:84 lut_35.scala 5707:47]
  wire  _GEN_11041 = read_stack10_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11013; // @[lut_35.scala 5687:84 lut_35.scala 5708:47]
  wire  _GEN_11042 = read_stack10_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11014; // @[lut_35.scala 5687:84 lut_35.scala 5709:47]
  wire  _GEN_11043 = read_stack10_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11015; // @[lut_35.scala 5687:84 lut_35.scala 5710:47]
  wire  _GEN_11044 = read_stack10_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11016; // @[lut_35.scala 5687:84 lut_35.scala 5711:47]
  wire  _GEN_11045 = read_stack10_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11017; // @[lut_35.scala 5687:84 lut_35.scala 5712:47]
  wire  _GEN_11046 = read_stack10_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11018; // @[lut_35.scala 5687:84 lut_35.scala 5713:47]
  wire  _GEN_11047 = read_stack10_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11019; // @[lut_35.scala 5687:84 lut_35.scala 5714:47]
  wire  _GEN_11048 = read_stack10_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11020; // @[lut_35.scala 5687:84 lut_35.scala 5715:47]
  wire  _GEN_11049 = read_stack10_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11021; // @[lut_35.scala 5687:84 lut_35.scala 5716:47]
  wire  _GEN_11050 = read_stack10_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11022; // @[lut_35.scala 5687:84 lut_35.scala 5717:47]
  wire  _GEN_11051 = read_stack10_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11023; // @[lut_35.scala 5687:84 lut_35.scala 5718:47]
  wire  _GEN_11052 = read_stack10_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11024; // @[lut_35.scala 5687:84 lut_35.scala 5719:47]
  wire  _GEN_11053 = read_stack10_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11025; // @[lut_35.scala 5687:84 lut_35.scala 5720:47]
  wire  _GEN_11054 = read_stack10_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11026; // @[lut_35.scala 5687:84 lut_35.scala 5721:47]
  wire  _GEN_11055 = read_stack10_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11027; // @[lut_35.scala 5687:84 lut_35.scala 5722:47]
  wire  _GEN_11060 = read_stack9_clear == clear_ray_id & clear_valid ? 1'h0 : _T_820; // @[lut_35.scala 5649:83 lut_35.scala 5660:47]
  wire  _GEN_11061 = read_stack9_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11032; // @[lut_35.scala 5649:83 lut_35.scala 5661:47]
  wire  _GEN_11062 = read_stack9_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11033; // @[lut_35.scala 5649:83 lut_35.scala 5662:47]
  wire  _GEN_11063 = read_stack9_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11034; // @[lut_35.scala 5649:83 lut_35.scala 5663:47]
  wire  _GEN_11064 = read_stack9_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11035; // @[lut_35.scala 5649:83 lut_35.scala 5664:47]
  wire  _GEN_11065 = read_stack9_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11036; // @[lut_35.scala 5649:83 lut_35.scala 5665:47]
  wire  _GEN_11066 = read_stack9_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11037; // @[lut_35.scala 5649:83 lut_35.scala 5666:47]
  wire  _GEN_11067 = read_stack9_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11038; // @[lut_35.scala 5649:83 lut_35.scala 5667:47]
  wire  _GEN_11068 = read_stack9_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11039; // @[lut_35.scala 5649:83 lut_35.scala 5668:47]
  wire  _GEN_11069 = read_stack9_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11040; // @[lut_35.scala 5649:83 lut_35.scala 5669:47]
  wire  _GEN_11070 = read_stack9_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11041; // @[lut_35.scala 5649:83 lut_35.scala 5670:47]
  wire  _GEN_11071 = read_stack9_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11042; // @[lut_35.scala 5649:83 lut_35.scala 5671:47]
  wire  _GEN_11072 = read_stack9_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11043; // @[lut_35.scala 5649:83 lut_35.scala 5672:47]
  wire  _GEN_11073 = read_stack9_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11044; // @[lut_35.scala 5649:83 lut_35.scala 5673:47]
  wire  _GEN_11074 = read_stack9_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11045; // @[lut_35.scala 5649:83 lut_35.scala 5674:47]
  wire  _GEN_11075 = read_stack9_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11046; // @[lut_35.scala 5649:83 lut_35.scala 5675:47]
  wire  _GEN_11076 = read_stack9_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11047; // @[lut_35.scala 5649:83 lut_35.scala 5676:47]
  wire  _GEN_11077 = read_stack9_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11048; // @[lut_35.scala 5649:83 lut_35.scala 5677:47]
  wire  _GEN_11078 = read_stack9_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11049; // @[lut_35.scala 5649:83 lut_35.scala 5678:47]
  wire  _GEN_11079 = read_stack9_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11050; // @[lut_35.scala 5649:83 lut_35.scala 5679:47]
  wire  _GEN_11080 = read_stack9_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11051; // @[lut_35.scala 5649:83 lut_35.scala 5680:47]
  wire  _GEN_11081 = read_stack9_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11052; // @[lut_35.scala 5649:83 lut_35.scala 5681:47]
  wire  _GEN_11082 = read_stack9_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11053; // @[lut_35.scala 5649:83 lut_35.scala 5682:47]
  wire  _GEN_11083 = read_stack9_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11054; // @[lut_35.scala 5649:83 lut_35.scala 5683:47]
  wire  _GEN_11084 = read_stack9_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11055; // @[lut_35.scala 5649:83 lut_35.scala 5684:47]
  wire  _GEN_11089 = read_stack8_clear == clear_ray_id & clear_valid ? 1'h0 : _T_817; // @[lut_35.scala 5611:83 lut_35.scala 5621:46]
  wire  _GEN_11090 = read_stack8_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11060; // @[lut_35.scala 5611:83 lut_35.scala 5622:47]
  wire  _GEN_11091 = read_stack8_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11061; // @[lut_35.scala 5611:83 lut_35.scala 5623:47]
  wire  _GEN_11092 = read_stack8_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11062; // @[lut_35.scala 5611:83 lut_35.scala 5624:47]
  wire  _GEN_11093 = read_stack8_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11063; // @[lut_35.scala 5611:83 lut_35.scala 5625:47]
  wire  _GEN_11094 = read_stack8_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11064; // @[lut_35.scala 5611:83 lut_35.scala 5626:47]
  wire  _GEN_11095 = read_stack8_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11065; // @[lut_35.scala 5611:83 lut_35.scala 5627:47]
  wire  _GEN_11096 = read_stack8_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11066; // @[lut_35.scala 5611:83 lut_35.scala 5628:47]
  wire  _GEN_11097 = read_stack8_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11067; // @[lut_35.scala 5611:83 lut_35.scala 5629:47]
  wire  _GEN_11098 = read_stack8_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11068; // @[lut_35.scala 5611:83 lut_35.scala 5630:47]
  wire  _GEN_11099 = read_stack8_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11069; // @[lut_35.scala 5611:83 lut_35.scala 5631:47]
  wire  _GEN_11100 = read_stack8_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11070; // @[lut_35.scala 5611:83 lut_35.scala 5632:47]
  wire  _GEN_11101 = read_stack8_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11071; // @[lut_35.scala 5611:83 lut_35.scala 5633:47]
  wire  _GEN_11102 = read_stack8_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11072; // @[lut_35.scala 5611:83 lut_35.scala 5634:47]
  wire  _GEN_11103 = read_stack8_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11073; // @[lut_35.scala 5611:83 lut_35.scala 5635:47]
  wire  _GEN_11104 = read_stack8_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11074; // @[lut_35.scala 5611:83 lut_35.scala 5636:47]
  wire  _GEN_11105 = read_stack8_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11075; // @[lut_35.scala 5611:83 lut_35.scala 5637:47]
  wire  _GEN_11106 = read_stack8_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11076; // @[lut_35.scala 5611:83 lut_35.scala 5638:47]
  wire  _GEN_11107 = read_stack8_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11077; // @[lut_35.scala 5611:83 lut_35.scala 5639:47]
  wire  _GEN_11108 = read_stack8_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11078; // @[lut_35.scala 5611:83 lut_35.scala 5640:47]
  wire  _GEN_11109 = read_stack8_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11079; // @[lut_35.scala 5611:83 lut_35.scala 5641:47]
  wire  _GEN_11110 = read_stack8_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11080; // @[lut_35.scala 5611:83 lut_35.scala 5642:47]
  wire  _GEN_11111 = read_stack8_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11081; // @[lut_35.scala 5611:83 lut_35.scala 5643:47]
  wire  _GEN_11112 = read_stack8_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11082; // @[lut_35.scala 5611:83 lut_35.scala 5644:47]
  wire  _GEN_11113 = read_stack8_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11083; // @[lut_35.scala 5611:83 lut_35.scala 5645:47]
  wire  _GEN_11114 = read_stack8_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11084; // @[lut_35.scala 5611:83 lut_35.scala 5646:47]
  wire  _GEN_11119 = read_stack7_clear == clear_ray_id & clear_valid ? 1'h0 : _T_814; // @[lut_35.scala 5573:83 lut_35.scala 5582:46]
  wire  _GEN_11120 = read_stack7_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11089; // @[lut_35.scala 5573:83 lut_35.scala 5583:46]
  wire  _GEN_11121 = read_stack7_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11090; // @[lut_35.scala 5573:83 lut_35.scala 5584:47]
  wire  _GEN_11122 = read_stack7_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11091; // @[lut_35.scala 5573:83 lut_35.scala 5585:47]
  wire  _GEN_11123 = read_stack7_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11092; // @[lut_35.scala 5573:83 lut_35.scala 5586:47]
  wire  _GEN_11124 = read_stack7_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11093; // @[lut_35.scala 5573:83 lut_35.scala 5587:47]
  wire  _GEN_11125 = read_stack7_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11094; // @[lut_35.scala 5573:83 lut_35.scala 5588:47]
  wire  _GEN_11126 = read_stack7_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11095; // @[lut_35.scala 5573:83 lut_35.scala 5589:47]
  wire  _GEN_11127 = read_stack7_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11096; // @[lut_35.scala 5573:83 lut_35.scala 5590:47]
  wire  _GEN_11128 = read_stack7_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11097; // @[lut_35.scala 5573:83 lut_35.scala 5591:47]
  wire  _GEN_11129 = read_stack7_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11098; // @[lut_35.scala 5573:83 lut_35.scala 5592:47]
  wire  _GEN_11130 = read_stack7_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11099; // @[lut_35.scala 5573:83 lut_35.scala 5593:47]
  wire  _GEN_11131 = read_stack7_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11100; // @[lut_35.scala 5573:83 lut_35.scala 5594:47]
  wire  _GEN_11132 = read_stack7_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11101; // @[lut_35.scala 5573:83 lut_35.scala 5595:47]
  wire  _GEN_11133 = read_stack7_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11102; // @[lut_35.scala 5573:83 lut_35.scala 5596:47]
  wire  _GEN_11134 = read_stack7_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11103; // @[lut_35.scala 5573:83 lut_35.scala 5597:47]
  wire  _GEN_11135 = read_stack7_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11104; // @[lut_35.scala 5573:83 lut_35.scala 5598:47]
  wire  _GEN_11136 = read_stack7_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11105; // @[lut_35.scala 5573:83 lut_35.scala 5599:47]
  wire  _GEN_11137 = read_stack7_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11106; // @[lut_35.scala 5573:83 lut_35.scala 5600:47]
  wire  _GEN_11138 = read_stack7_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11107; // @[lut_35.scala 5573:83 lut_35.scala 5601:47]
  wire  _GEN_11139 = read_stack7_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11108; // @[lut_35.scala 5573:83 lut_35.scala 5602:47]
  wire  _GEN_11140 = read_stack7_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11109; // @[lut_35.scala 5573:83 lut_35.scala 5603:47]
  wire  _GEN_11141 = read_stack7_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11110; // @[lut_35.scala 5573:83 lut_35.scala 5604:47]
  wire  _GEN_11142 = read_stack7_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11111; // @[lut_35.scala 5573:83 lut_35.scala 5605:47]
  wire  _GEN_11143 = read_stack7_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11112; // @[lut_35.scala 5573:83 lut_35.scala 5606:47]
  wire  _GEN_11144 = read_stack7_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11113; // @[lut_35.scala 5573:83 lut_35.scala 5607:47]
  wire  _GEN_11145 = read_stack7_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11114; // @[lut_35.scala 5573:83 lut_35.scala 5608:47]
  wire  _GEN_11150 = read_stack6_clear == clear_ray_id & clear_valid ? 1'h0 : _T_811; // @[lut_35.scala 5535:83 lut_35.scala 5543:46]
  wire  _GEN_11151 = read_stack6_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11119; // @[lut_35.scala 5535:83 lut_35.scala 5544:46]
  wire  _GEN_11152 = read_stack6_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11120; // @[lut_35.scala 5535:83 lut_35.scala 5545:46]
  wire  _GEN_11153 = read_stack6_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11121; // @[lut_35.scala 5535:83 lut_35.scala 5546:47]
  wire  _GEN_11154 = read_stack6_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11122; // @[lut_35.scala 5535:83 lut_35.scala 5547:47]
  wire  _GEN_11155 = read_stack6_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11123; // @[lut_35.scala 5535:83 lut_35.scala 5548:47]
  wire  _GEN_11156 = read_stack6_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11124; // @[lut_35.scala 5535:83 lut_35.scala 5549:47]
  wire  _GEN_11157 = read_stack6_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11125; // @[lut_35.scala 5535:83 lut_35.scala 5550:47]
  wire  _GEN_11158 = read_stack6_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11126; // @[lut_35.scala 5535:83 lut_35.scala 5551:47]
  wire  _GEN_11159 = read_stack6_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11127; // @[lut_35.scala 5535:83 lut_35.scala 5552:47]
  wire  _GEN_11160 = read_stack6_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11128; // @[lut_35.scala 5535:83 lut_35.scala 5553:47]
  wire  _GEN_11161 = read_stack6_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11129; // @[lut_35.scala 5535:83 lut_35.scala 5554:47]
  wire  _GEN_11162 = read_stack6_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11130; // @[lut_35.scala 5535:83 lut_35.scala 5555:47]
  wire  _GEN_11163 = read_stack6_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11131; // @[lut_35.scala 5535:83 lut_35.scala 5556:47]
  wire  _GEN_11164 = read_stack6_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11132; // @[lut_35.scala 5535:83 lut_35.scala 5557:47]
  wire  _GEN_11165 = read_stack6_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11133; // @[lut_35.scala 5535:83 lut_35.scala 5558:47]
  wire  _GEN_11166 = read_stack6_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11134; // @[lut_35.scala 5535:83 lut_35.scala 5559:47]
  wire  _GEN_11167 = read_stack6_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11135; // @[lut_35.scala 5535:83 lut_35.scala 5560:47]
  wire  _GEN_11168 = read_stack6_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11136; // @[lut_35.scala 5535:83 lut_35.scala 5561:47]
  wire  _GEN_11169 = read_stack6_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11137; // @[lut_35.scala 5535:83 lut_35.scala 5562:47]
  wire  _GEN_11170 = read_stack6_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11138; // @[lut_35.scala 5535:83 lut_35.scala 5563:47]
  wire  _GEN_11171 = read_stack6_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11139; // @[lut_35.scala 5535:83 lut_35.scala 5564:47]
  wire  _GEN_11172 = read_stack6_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11140; // @[lut_35.scala 5535:83 lut_35.scala 5565:47]
  wire  _GEN_11173 = read_stack6_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11141; // @[lut_35.scala 5535:83 lut_35.scala 5566:47]
  wire  _GEN_11174 = read_stack6_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11142; // @[lut_35.scala 5535:83 lut_35.scala 5567:47]
  wire  _GEN_11175 = read_stack6_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11143; // @[lut_35.scala 5535:83 lut_35.scala 5568:47]
  wire  _GEN_11176 = read_stack6_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11144; // @[lut_35.scala 5535:83 lut_35.scala 5569:47]
  wire  _GEN_11177 = read_stack6_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11145; // @[lut_35.scala 5535:83 lut_35.scala 5570:47]
  wire  _GEN_11182 = read_stack5_clear == clear_ray_id & clear_valid ? 1'h0 : _T_808; // @[lut_35.scala 5497:83 lut_35.scala 5504:46]
  wire  _GEN_11183 = read_stack5_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11150; // @[lut_35.scala 5497:83 lut_35.scala 5505:46]
  wire  _GEN_11184 = read_stack5_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11151; // @[lut_35.scala 5497:83 lut_35.scala 5506:46]
  wire  _GEN_11185 = read_stack5_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11152; // @[lut_35.scala 5497:83 lut_35.scala 5507:46]
  wire  _GEN_11186 = read_stack5_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11153; // @[lut_35.scala 5497:83 lut_35.scala 5508:47]
  wire  _GEN_11187 = read_stack5_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11154; // @[lut_35.scala 5497:83 lut_35.scala 5509:47]
  wire  _GEN_11188 = read_stack5_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11155; // @[lut_35.scala 5497:83 lut_35.scala 5510:47]
  wire  _GEN_11189 = read_stack5_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11156; // @[lut_35.scala 5497:83 lut_35.scala 5511:47]
  wire  _GEN_11190 = read_stack5_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11157; // @[lut_35.scala 5497:83 lut_35.scala 5512:47]
  wire  _GEN_11191 = read_stack5_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11158; // @[lut_35.scala 5497:83 lut_35.scala 5513:47]
  wire  _GEN_11192 = read_stack5_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11159; // @[lut_35.scala 5497:83 lut_35.scala 5514:47]
  wire  _GEN_11193 = read_stack5_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11160; // @[lut_35.scala 5497:83 lut_35.scala 5515:47]
  wire  _GEN_11194 = read_stack5_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11161; // @[lut_35.scala 5497:83 lut_35.scala 5516:47]
  wire  _GEN_11195 = read_stack5_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11162; // @[lut_35.scala 5497:83 lut_35.scala 5517:47]
  wire  _GEN_11196 = read_stack5_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11163; // @[lut_35.scala 5497:83 lut_35.scala 5518:47]
  wire  _GEN_11197 = read_stack5_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11164; // @[lut_35.scala 5497:83 lut_35.scala 5519:47]
  wire  _GEN_11198 = read_stack5_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11165; // @[lut_35.scala 5497:83 lut_35.scala 5520:47]
  wire  _GEN_11199 = read_stack5_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11166; // @[lut_35.scala 5497:83 lut_35.scala 5521:47]
  wire  _GEN_11200 = read_stack5_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11167; // @[lut_35.scala 5497:83 lut_35.scala 5522:47]
  wire  _GEN_11201 = read_stack5_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11168; // @[lut_35.scala 5497:83 lut_35.scala 5523:47]
  wire  _GEN_11202 = read_stack5_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11169; // @[lut_35.scala 5497:83 lut_35.scala 5524:47]
  wire  _GEN_11203 = read_stack5_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11170; // @[lut_35.scala 5497:83 lut_35.scala 5525:47]
  wire  _GEN_11204 = read_stack5_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11171; // @[lut_35.scala 5497:83 lut_35.scala 5526:47]
  wire  _GEN_11205 = read_stack5_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11172; // @[lut_35.scala 5497:83 lut_35.scala 5527:47]
  wire  _GEN_11206 = read_stack5_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11173; // @[lut_35.scala 5497:83 lut_35.scala 5528:47]
  wire  _GEN_11207 = read_stack5_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11174; // @[lut_35.scala 5497:83 lut_35.scala 5529:47]
  wire  _GEN_11208 = read_stack5_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11175; // @[lut_35.scala 5497:83 lut_35.scala 5530:47]
  wire  _GEN_11209 = read_stack5_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11176; // @[lut_35.scala 5497:83 lut_35.scala 5531:47]
  wire  _GEN_11210 = read_stack5_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11177; // @[lut_35.scala 5497:83 lut_35.scala 5532:47]
  wire  _GEN_11215 = read_stack4_clear == clear_ray_id & clear_valid ? 1'h0 : _T_805; // @[lut_35.scala 5459:83 lut_35.scala 5465:46]
  wire  _GEN_11216 = read_stack4_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11182; // @[lut_35.scala 5459:83 lut_35.scala 5466:46]
  wire  _GEN_11217 = read_stack4_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11183; // @[lut_35.scala 5459:83 lut_35.scala 5467:46]
  wire  _GEN_11218 = read_stack4_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11184; // @[lut_35.scala 5459:83 lut_35.scala 5468:46]
  wire  _GEN_11219 = read_stack4_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11185; // @[lut_35.scala 5459:83 lut_35.scala 5469:46]
  wire  _GEN_11220 = read_stack4_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11186; // @[lut_35.scala 5459:83 lut_35.scala 5470:47]
  wire  _GEN_11221 = read_stack4_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11187; // @[lut_35.scala 5459:83 lut_35.scala 5471:47]
  wire  _GEN_11222 = read_stack4_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11188; // @[lut_35.scala 5459:83 lut_35.scala 5472:47]
  wire  _GEN_11223 = read_stack4_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11189; // @[lut_35.scala 5459:83 lut_35.scala 5473:47]
  wire  _GEN_11224 = read_stack4_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11190; // @[lut_35.scala 5459:83 lut_35.scala 5474:47]
  wire  _GEN_11225 = read_stack4_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11191; // @[lut_35.scala 5459:83 lut_35.scala 5475:47]
  wire  _GEN_11226 = read_stack4_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11192; // @[lut_35.scala 5459:83 lut_35.scala 5476:47]
  wire  _GEN_11227 = read_stack4_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11193; // @[lut_35.scala 5459:83 lut_35.scala 5477:47]
  wire  _GEN_11228 = read_stack4_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11194; // @[lut_35.scala 5459:83 lut_35.scala 5478:47]
  wire  _GEN_11229 = read_stack4_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11195; // @[lut_35.scala 5459:83 lut_35.scala 5479:47]
  wire  _GEN_11230 = read_stack4_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11196; // @[lut_35.scala 5459:83 lut_35.scala 5480:47]
  wire  _GEN_11231 = read_stack4_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11197; // @[lut_35.scala 5459:83 lut_35.scala 5481:47]
  wire  _GEN_11232 = read_stack4_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11198; // @[lut_35.scala 5459:83 lut_35.scala 5482:47]
  wire  _GEN_11233 = read_stack4_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11199; // @[lut_35.scala 5459:83 lut_35.scala 5483:47]
  wire  _GEN_11234 = read_stack4_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11200; // @[lut_35.scala 5459:83 lut_35.scala 5484:47]
  wire  _GEN_11235 = read_stack4_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11201; // @[lut_35.scala 5459:83 lut_35.scala 5485:47]
  wire  _GEN_11236 = read_stack4_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11202; // @[lut_35.scala 5459:83 lut_35.scala 5486:47]
  wire  _GEN_11237 = read_stack4_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11203; // @[lut_35.scala 5459:83 lut_35.scala 5487:47]
  wire  _GEN_11238 = read_stack4_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11204; // @[lut_35.scala 5459:83 lut_35.scala 5488:47]
  wire  _GEN_11239 = read_stack4_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11205; // @[lut_35.scala 5459:83 lut_35.scala 5489:47]
  wire  _GEN_11240 = read_stack4_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11206; // @[lut_35.scala 5459:83 lut_35.scala 5490:47]
  wire  _GEN_11241 = read_stack4_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11207; // @[lut_35.scala 5459:83 lut_35.scala 5491:47]
  wire  _GEN_11242 = read_stack4_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11208; // @[lut_35.scala 5459:83 lut_35.scala 5492:47]
  wire  _GEN_11243 = read_stack4_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11209; // @[lut_35.scala 5459:83 lut_35.scala 5493:47]
  wire  _GEN_11244 = read_stack4_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11210; // @[lut_35.scala 5459:83 lut_35.scala 5494:47]
  wire  _GEN_11249 = _T_796 ? 1'h0 : _T_802; // @[lut_35.scala 5421:83 lut_35.scala 5426:46]
  wire  _GEN_11250 = _T_796 ? 1'h0 : _GEN_11215; // @[lut_35.scala 5421:83 lut_35.scala 5427:46]
  wire  _GEN_11251 = _T_796 ? 1'h0 : _GEN_11216; // @[lut_35.scala 5421:83 lut_35.scala 5428:46]
  wire  _GEN_11252 = _T_796 ? 1'h0 : _GEN_11217; // @[lut_35.scala 5421:83 lut_35.scala 5429:46]
  wire  _GEN_11253 = _T_796 ? 1'h0 : _GEN_11218; // @[lut_35.scala 5421:83 lut_35.scala 5430:46]
  wire  _GEN_11254 = _T_796 ? 1'h0 : _GEN_11219; // @[lut_35.scala 5421:83 lut_35.scala 5431:46]
  wire  _GEN_11255 = _T_796 ? 1'h0 : _GEN_11220; // @[lut_35.scala 5421:83 lut_35.scala 5432:47]
  wire  _GEN_11256 = _T_796 ? 1'h0 : _GEN_11221; // @[lut_35.scala 5421:83 lut_35.scala 5433:47]
  wire  _GEN_11257 = _T_796 ? 1'h0 : _GEN_11222; // @[lut_35.scala 5421:83 lut_35.scala 5434:47]
  wire  _GEN_11258 = _T_796 ? 1'h0 : _GEN_11223; // @[lut_35.scala 5421:83 lut_35.scala 5435:47]
  wire  _GEN_11259 = _T_796 ? 1'h0 : _GEN_11224; // @[lut_35.scala 5421:83 lut_35.scala 5436:47]
  wire  _GEN_11260 = _T_796 ? 1'h0 : _GEN_11225; // @[lut_35.scala 5421:83 lut_35.scala 5437:47]
  wire  _GEN_11261 = _T_796 ? 1'h0 : _GEN_11226; // @[lut_35.scala 5421:83 lut_35.scala 5438:47]
  wire  _GEN_11262 = _T_796 ? 1'h0 : _GEN_11227; // @[lut_35.scala 5421:83 lut_35.scala 5439:47]
  wire  _GEN_11263 = _T_796 ? 1'h0 : _GEN_11228; // @[lut_35.scala 5421:83 lut_35.scala 5440:47]
  wire  _GEN_11264 = _T_796 ? 1'h0 : _GEN_11229; // @[lut_35.scala 5421:83 lut_35.scala 5441:47]
  wire  _GEN_11265 = _T_796 ? 1'h0 : _GEN_11230; // @[lut_35.scala 5421:83 lut_35.scala 5442:47]
  wire  _GEN_11266 = _T_796 ? 1'h0 : _GEN_11231; // @[lut_35.scala 5421:83 lut_35.scala 5443:47]
  wire  _GEN_11267 = _T_796 ? 1'h0 : _GEN_11232; // @[lut_35.scala 5421:83 lut_35.scala 5444:47]
  wire  _GEN_11268 = _T_796 ? 1'h0 : _GEN_11233; // @[lut_35.scala 5421:83 lut_35.scala 5445:47]
  wire  _GEN_11269 = _T_796 ? 1'h0 : _GEN_11234; // @[lut_35.scala 5421:83 lut_35.scala 5446:47]
  wire  _GEN_11270 = _T_796 ? 1'h0 : _GEN_11235; // @[lut_35.scala 5421:83 lut_35.scala 5447:47]
  wire  _GEN_11271 = _T_796 ? 1'h0 : _GEN_11236; // @[lut_35.scala 5421:83 lut_35.scala 5448:47]
  wire  _GEN_11272 = _T_796 ? 1'h0 : _GEN_11237; // @[lut_35.scala 5421:83 lut_35.scala 5449:47]
  wire  _GEN_11273 = _T_796 ? 1'h0 : _GEN_11238; // @[lut_35.scala 5421:83 lut_35.scala 5450:47]
  wire  _GEN_11274 = _T_796 ? 1'h0 : _GEN_11239; // @[lut_35.scala 5421:83 lut_35.scala 5451:47]
  wire  _GEN_11275 = _T_796 ? 1'h0 : _GEN_11240; // @[lut_35.scala 5421:83 lut_35.scala 5452:47]
  wire  _GEN_11276 = _T_796 ? 1'h0 : _GEN_11241; // @[lut_35.scala 5421:83 lut_35.scala 5453:47]
  wire  _GEN_11277 = _T_796 ? 1'h0 : _GEN_11242; // @[lut_35.scala 5421:83 lut_35.scala 5454:47]
  wire  _GEN_11278 = _T_796 ? 1'h0 : _GEN_11243; // @[lut_35.scala 5421:83 lut_35.scala 5455:47]
  wire  _GEN_11279 = _T_796 ? 1'h0 : _GEN_11244; // @[lut_35.scala 5421:83 lut_35.scala 5456:47]
  wire  _GEN_11284 = read_stack3_clear == clear_ray_id & clear_valid ? 1'h0 : read_stack3_clear == clear_ray_id &
    clear_valid; // @[lut_35.scala 5383:83 lut_35.scala 5387:46]
  wire  _GEN_11285 = read_stack3_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11249; // @[lut_35.scala 5383:83 lut_35.scala 5388:46]
  wire  _GEN_11286 = read_stack3_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11250; // @[lut_35.scala 5383:83 lut_35.scala 5389:46]
  wire  _GEN_11287 = read_stack3_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11251; // @[lut_35.scala 5383:83 lut_35.scala 5390:46]
  wire  _GEN_11288 = read_stack3_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11252; // @[lut_35.scala 5383:83 lut_35.scala 5391:46]
  wire  _GEN_11289 = read_stack3_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11253; // @[lut_35.scala 5383:83 lut_35.scala 5392:46]
  wire  _GEN_11290 = read_stack3_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11254; // @[lut_35.scala 5383:83 lut_35.scala 5393:46]
  wire  _GEN_11291 = read_stack3_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11255; // @[lut_35.scala 5383:83 lut_35.scala 5394:47]
  wire  _GEN_11292 = read_stack3_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11256; // @[lut_35.scala 5383:83 lut_35.scala 5395:47]
  wire  _GEN_11293 = read_stack3_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11257; // @[lut_35.scala 5383:83 lut_35.scala 5396:47]
  wire  _GEN_11294 = read_stack3_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11258; // @[lut_35.scala 5383:83 lut_35.scala 5397:47]
  wire  _GEN_11295 = read_stack3_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11259; // @[lut_35.scala 5383:83 lut_35.scala 5398:47]
  wire  _GEN_11296 = read_stack3_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11260; // @[lut_35.scala 5383:83 lut_35.scala 5399:47]
  wire  _GEN_11297 = read_stack3_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11261; // @[lut_35.scala 5383:83 lut_35.scala 5400:47]
  wire  _GEN_11298 = read_stack3_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11262; // @[lut_35.scala 5383:83 lut_35.scala 5401:47]
  wire  _GEN_11299 = read_stack3_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11263; // @[lut_35.scala 5383:83 lut_35.scala 5402:47]
  wire  _GEN_11300 = read_stack3_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11264; // @[lut_35.scala 5383:83 lut_35.scala 5403:47]
  wire  _GEN_11301 = read_stack3_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11265; // @[lut_35.scala 5383:83 lut_35.scala 5404:47]
  wire  _GEN_11302 = read_stack3_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11266; // @[lut_35.scala 5383:83 lut_35.scala 5405:47]
  wire  _GEN_11303 = read_stack3_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11267; // @[lut_35.scala 5383:83 lut_35.scala 5406:47]
  wire  _GEN_11304 = read_stack3_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11268; // @[lut_35.scala 5383:83 lut_35.scala 5407:47]
  wire  _GEN_11305 = read_stack3_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11269; // @[lut_35.scala 5383:83 lut_35.scala 5408:47]
  wire  _GEN_11306 = read_stack3_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11270; // @[lut_35.scala 5383:83 lut_35.scala 5409:47]
  wire  _GEN_11307 = read_stack3_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11271; // @[lut_35.scala 5383:83 lut_35.scala 5410:47]
  wire  _GEN_11308 = read_stack3_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11272; // @[lut_35.scala 5383:83 lut_35.scala 5411:47]
  wire  _GEN_11309 = read_stack3_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11273; // @[lut_35.scala 5383:83 lut_35.scala 5412:47]
  wire  _GEN_11310 = read_stack3_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11274; // @[lut_35.scala 5383:83 lut_35.scala 5413:47]
  wire  _GEN_11311 = read_stack3_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11275; // @[lut_35.scala 5383:83 lut_35.scala 5414:47]
  wire  _GEN_11312 = read_stack3_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11276; // @[lut_35.scala 5383:83 lut_35.scala 5415:47]
  wire  _GEN_11313 = read_stack3_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11277; // @[lut_35.scala 5383:83 lut_35.scala 5416:47]
  wire  _GEN_11314 = read_stack3_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11278; // @[lut_35.scala 5383:83 lut_35.scala 5417:47]
  wire  _GEN_11315 = read_stack3_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11279; // @[lut_35.scala 5383:83 lut_35.scala 5418:47]
  wire  _GEN_11320 = read_stack1_clear == clear_ray_id & clear_valid ? 1'h0 : _T_796; // @[lut_35.scala 5345:83 lut_35.scala 5348:46]
  wire  _GEN_11321 = read_stack1_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11284; // @[lut_35.scala 5345:83 lut_35.scala 5349:46]
  wire  _GEN_11322 = read_stack1_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11285; // @[lut_35.scala 5345:83 lut_35.scala 5350:46]
  wire  _GEN_11323 = read_stack1_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11286; // @[lut_35.scala 5345:83 lut_35.scala 5351:46]
  wire  _GEN_11324 = read_stack1_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11287; // @[lut_35.scala 5345:83 lut_35.scala 5352:46]
  wire  _GEN_11325 = read_stack1_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11288; // @[lut_35.scala 5345:83 lut_35.scala 5353:46]
  wire  _GEN_11326 = read_stack1_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11289; // @[lut_35.scala 5345:83 lut_35.scala 5354:46]
  wire  _GEN_11327 = read_stack1_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11290; // @[lut_35.scala 5345:83 lut_35.scala 5355:46]
  wire  _GEN_11328 = read_stack1_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11291; // @[lut_35.scala 5345:83 lut_35.scala 5356:47]
  wire  _GEN_11329 = read_stack1_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11292; // @[lut_35.scala 5345:83 lut_35.scala 5357:47]
  wire  _GEN_11330 = read_stack1_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11293; // @[lut_35.scala 5345:83 lut_35.scala 5358:47]
  wire  _GEN_11331 = read_stack1_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11294; // @[lut_35.scala 5345:83 lut_35.scala 5359:47]
  wire  _GEN_11332 = read_stack1_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11295; // @[lut_35.scala 5345:83 lut_35.scala 5360:47]
  wire  _GEN_11333 = read_stack1_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11296; // @[lut_35.scala 5345:83 lut_35.scala 5361:47]
  wire  _GEN_11334 = read_stack1_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11297; // @[lut_35.scala 5345:83 lut_35.scala 5362:47]
  wire  _GEN_11335 = read_stack1_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11298; // @[lut_35.scala 5345:83 lut_35.scala 5363:47]
  wire  _GEN_11336 = read_stack1_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11299; // @[lut_35.scala 5345:83 lut_35.scala 5364:47]
  wire  _GEN_11337 = read_stack1_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11300; // @[lut_35.scala 5345:83 lut_35.scala 5365:47]
  wire  _GEN_11338 = read_stack1_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11301; // @[lut_35.scala 5345:83 lut_35.scala 5366:47]
  wire  _GEN_11339 = read_stack1_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11302; // @[lut_35.scala 5345:83 lut_35.scala 5367:47]
  wire  _GEN_11340 = read_stack1_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11303; // @[lut_35.scala 5345:83 lut_35.scala 5368:47]
  wire  _GEN_11341 = read_stack1_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11304; // @[lut_35.scala 5345:83 lut_35.scala 5369:47]
  wire  _GEN_11342 = read_stack1_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11305; // @[lut_35.scala 5345:83 lut_35.scala 5370:47]
  wire  _GEN_11343 = read_stack1_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11306; // @[lut_35.scala 5345:83 lut_35.scala 5371:47]
  wire  _GEN_11344 = read_stack1_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11307; // @[lut_35.scala 5345:83 lut_35.scala 5372:47]
  wire  _GEN_11345 = read_stack1_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11308; // @[lut_35.scala 5345:83 lut_35.scala 5373:47]
  wire  _GEN_11346 = read_stack1_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11309; // @[lut_35.scala 5345:83 lut_35.scala 5374:47]
  wire  _GEN_11347 = read_stack1_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11310; // @[lut_35.scala 5345:83 lut_35.scala 5375:47]
  wire  _GEN_11348 = read_stack1_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11311; // @[lut_35.scala 5345:83 lut_35.scala 5376:47]
  wire  _GEN_11349 = read_stack1_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11312; // @[lut_35.scala 5345:83 lut_35.scala 5377:47]
  wire  _GEN_11350 = read_stack1_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11313; // @[lut_35.scala 5345:83 lut_35.scala 5378:47]
  wire  _GEN_11351 = read_stack1_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11314; // @[lut_35.scala 5345:83 lut_35.scala 5379:47]
  wire  _GEN_11352 = read_stack1_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11315; // @[lut_35.scala 5345:83 lut_35.scala 5380:47]
  wire  _GEN_11356 = read_stack0_clear == clear_ray_id & clear_valid ? 1'h0 : _T_793; // @[lut_35.scala 5307:73 lut_35.scala 5309:42]
  wire  _GEN_11357 = read_stack0_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11320; // @[lut_35.scala 5307:73 lut_35.scala 5310:42]
  wire  _GEN_11358 = read_stack0_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11321; // @[lut_35.scala 5307:73 lut_35.scala 5311:42]
  wire  _GEN_11359 = read_stack0_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11322; // @[lut_35.scala 5307:73 lut_35.scala 5312:42]
  wire  _GEN_11360 = read_stack0_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11323; // @[lut_35.scala 5307:73 lut_35.scala 5313:42]
  wire  _GEN_11361 = read_stack0_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11324; // @[lut_35.scala 5307:73 lut_35.scala 5314:42]
  wire  _GEN_11362 = read_stack0_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11325; // @[lut_35.scala 5307:73 lut_35.scala 5315:42]
  wire  _GEN_11363 = read_stack0_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11326; // @[lut_35.scala 5307:73 lut_35.scala 5316:42]
  wire  _GEN_11364 = read_stack0_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11327; // @[lut_35.scala 5307:73 lut_35.scala 5317:42]
  wire  _GEN_11365 = read_stack0_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11328; // @[lut_35.scala 5307:73 lut_35.scala 5318:43]
  wire  _GEN_11366 = read_stack0_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11329; // @[lut_35.scala 5307:73 lut_35.scala 5319:43]
  wire  _GEN_11367 = read_stack0_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11330; // @[lut_35.scala 5307:73 lut_35.scala 5320:43]
  wire  _GEN_11368 = read_stack0_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11331; // @[lut_35.scala 5307:73 lut_35.scala 5321:43]
  wire  _GEN_11369 = read_stack0_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11332; // @[lut_35.scala 5307:73 lut_35.scala 5322:43]
  wire  _GEN_11370 = read_stack0_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11333; // @[lut_35.scala 5307:73 lut_35.scala 5323:43]
  wire  _GEN_11371 = read_stack0_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11334; // @[lut_35.scala 5307:73 lut_35.scala 5324:43]
  wire  _GEN_11372 = read_stack0_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11335; // @[lut_35.scala 5307:73 lut_35.scala 5325:43]
  wire  _GEN_11373 = read_stack0_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11336; // @[lut_35.scala 5307:73 lut_35.scala 5326:43]
  wire  _GEN_11374 = read_stack0_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11337; // @[lut_35.scala 5307:73 lut_35.scala 5327:43]
  wire  _GEN_11375 = read_stack0_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11338; // @[lut_35.scala 5307:73 lut_35.scala 5328:43]
  wire  _GEN_11376 = read_stack0_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11339; // @[lut_35.scala 5307:73 lut_35.scala 5329:43]
  wire  _GEN_11377 = read_stack0_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11340; // @[lut_35.scala 5307:73 lut_35.scala 5330:43]
  wire  _GEN_11378 = read_stack0_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11341; // @[lut_35.scala 5307:73 lut_35.scala 5331:43]
  wire  _GEN_11379 = read_stack0_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11342; // @[lut_35.scala 5307:73 lut_35.scala 5332:43]
  wire  _GEN_11380 = read_stack0_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11343; // @[lut_35.scala 5307:73 lut_35.scala 5333:43]
  wire  _GEN_11381 = read_stack0_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11344; // @[lut_35.scala 5307:73 lut_35.scala 5334:43]
  wire  _GEN_11382 = read_stack0_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11345; // @[lut_35.scala 5307:73 lut_35.scala 5335:43]
  wire  _GEN_11383 = read_stack0_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11346; // @[lut_35.scala 5307:73 lut_35.scala 5336:43]
  wire  _GEN_11384 = read_stack0_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11347; // @[lut_35.scala 5307:73 lut_35.scala 5337:43]
  wire  _GEN_11385 = read_stack0_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11348; // @[lut_35.scala 5307:73 lut_35.scala 5338:43]
  wire  _GEN_11386 = read_stack0_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11349; // @[lut_35.scala 5307:73 lut_35.scala 5339:43]
  wire  _GEN_11387 = read_stack0_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11350; // @[lut_35.scala 5307:73 lut_35.scala 5340:43]
  wire  _GEN_11388 = read_stack0_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11351; // @[lut_35.scala 5307:73 lut_35.scala 5341:43]
  wire  _GEN_11389 = read_stack0_clear == clear_ray_id & clear_valid ? 1'h0 : _GEN_11352; // @[lut_35.scala 5307:73 lut_35.scala 5342:43]
  wire  _GEN_11392 = clear_1 & clear_valid & _T_790; // @[lut_35.scala 5306:51 lut_35.scala 6676:42]
  wire  _GEN_11393 = clear_1 & clear_valid & _GEN_11356; // @[lut_35.scala 5306:51 lut_35.scala 6677:42]
  wire  _GEN_11394 = clear_1 & clear_valid & _GEN_11357; // @[lut_35.scala 5306:51 lut_35.scala 6678:42]
  wire  _GEN_11395 = clear_1 & clear_valid & _GEN_11358; // @[lut_35.scala 5306:51 lut_35.scala 6679:42]
  wire  _GEN_11396 = clear_1 & clear_valid & _GEN_11359; // @[lut_35.scala 5306:51 lut_35.scala 6680:42]
  wire  _GEN_11397 = clear_1 & clear_valid & _GEN_11360; // @[lut_35.scala 5306:51 lut_35.scala 6681:42]
  wire  _GEN_11398 = clear_1 & clear_valid & _GEN_11361; // @[lut_35.scala 5306:51 lut_35.scala 6682:42]
  wire  _GEN_11399 = clear_1 & clear_valid & _GEN_11362; // @[lut_35.scala 5306:51 lut_35.scala 6683:42]
  wire  _GEN_11400 = clear_1 & clear_valid & _GEN_11363; // @[lut_35.scala 5306:51 lut_35.scala 6684:42]
  wire  _GEN_11401 = clear_1 & clear_valid & _GEN_11364; // @[lut_35.scala 5306:51 lut_35.scala 6685:42]
  wire  _GEN_11402 = clear_1 & clear_valid & _GEN_11365; // @[lut_35.scala 5306:51 lut_35.scala 6686:43]
  wire  _GEN_11403 = clear_1 & clear_valid & _GEN_11366; // @[lut_35.scala 5306:51 lut_35.scala 6687:43]
  wire  _GEN_11404 = clear_1 & clear_valid & _GEN_11367; // @[lut_35.scala 5306:51 lut_35.scala 6688:43]
  wire  _GEN_11405 = clear_1 & clear_valid & _GEN_11368; // @[lut_35.scala 5306:51 lut_35.scala 6689:43]
  wire  _GEN_11406 = clear_1 & clear_valid & _GEN_11369; // @[lut_35.scala 5306:51 lut_35.scala 6690:43]
  wire  _GEN_11407 = clear_1 & clear_valid & _GEN_11370; // @[lut_35.scala 5306:51 lut_35.scala 6691:43]
  wire  _GEN_11408 = clear_1 & clear_valid & _GEN_11371; // @[lut_35.scala 5306:51 lut_35.scala 6692:43]
  wire  _GEN_11409 = clear_1 & clear_valid & _GEN_11372; // @[lut_35.scala 5306:51 lut_35.scala 6693:43]
  wire  _GEN_11410 = clear_1 & clear_valid & _GEN_11373; // @[lut_35.scala 5306:51 lut_35.scala 6694:43]
  wire  _GEN_11411 = clear_1 & clear_valid & _GEN_11374; // @[lut_35.scala 5306:51 lut_35.scala 6695:43]
  wire  _GEN_11412 = clear_1 & clear_valid & _GEN_11375; // @[lut_35.scala 5306:51 lut_35.scala 6696:43]
  wire  _GEN_11413 = clear_1 & clear_valid & _GEN_11376; // @[lut_35.scala 5306:51 lut_35.scala 6697:43]
  wire  _GEN_11414 = clear_1 & clear_valid & _GEN_11377; // @[lut_35.scala 5306:51 lut_35.scala 6698:43]
  wire  _GEN_11415 = clear_1 & clear_valid & _GEN_11378; // @[lut_35.scala 5306:51 lut_35.scala 6699:43]
  wire  _GEN_11416 = clear_1 & clear_valid & _GEN_11379; // @[lut_35.scala 5306:51 lut_35.scala 6700:43]
  wire  _GEN_11417 = clear_1 & clear_valid & _GEN_11380; // @[lut_35.scala 5306:51 lut_35.scala 6701:43]
  wire  _GEN_11418 = clear_1 & clear_valid & _GEN_11381; // @[lut_35.scala 5306:51 lut_35.scala 6702:43]
  wire  _GEN_11419 = clear_1 & clear_valid & _GEN_11382; // @[lut_35.scala 5306:51 lut_35.scala 6703:43]
  wire  _GEN_11420 = clear_1 & clear_valid & _GEN_11383; // @[lut_35.scala 5306:51 lut_35.scala 6704:43]
  wire  _GEN_11421 = clear_1 & clear_valid & _GEN_11384; // @[lut_35.scala 5306:51 lut_35.scala 6705:43]
  wire  _GEN_11422 = clear_1 & clear_valid & _GEN_11385; // @[lut_35.scala 5306:51 lut_35.scala 6706:43]
  wire  _GEN_11423 = clear_1 & clear_valid & _GEN_11386; // @[lut_35.scala 5306:51 lut_35.scala 6707:43]
  wire  _GEN_11424 = clear_1 & clear_valid & _GEN_11387; // @[lut_35.scala 5306:51 lut_35.scala 6708:43]
  wire  _GEN_11425 = clear_1 & clear_valid & _GEN_11388; // @[lut_35.scala 5306:51 lut_35.scala 6709:43]
  wire  _GEN_11426 = clear_1 & clear_valid & _GEN_11389; // @[lut_35.scala 5306:51 lut_35.scala 6710:43]
  wire  _T_895 = dispatch_reg_0 | clear_0_1; // @[lut_35.scala 6754:33]
  wire [31:0] lo = LUT_mem_MPORT_176_data[31:0]; // @[lut_35.scala 6755:43]
  wire  _T_897 = push_mem_temp == 6'h0; // @[lut_35.scala 6756:30]
  wire  _GEN_11436 = push_mem_temp == 6'h0 ? 1'h0 : 1'h1; // @[lut_35.scala 6756:38 lut_35.scala 216:26 lut_35.scala 6759:16]
  wire  _T_901 = dispatch_reg_1 | clear_1_1; // @[lut_35.scala 6762:33]
  wire [31:0] lo_1 = LUT_mem_MPORT_181_data[31:0]; // @[lut_35.scala 6763:42]
  wire  _T_903 = push_mem_temp == 6'h1; // @[lut_35.scala 6764:30]
  wire  _GEN_11460 = push_mem_temp == 6'h1 ? 1'h0 : 1'h1; // @[lut_35.scala 6764:38 lut_35.scala 216:26 lut_35.scala 6767:16]
  wire  _T_907 = dispatch_reg_2 | clear_2_1; // @[lut_35.scala 6770:33]
  wire [31:0] lo_2 = LUT_mem_MPORT_186_data[31:0]; // @[lut_35.scala 6771:42]
  wire  _T_909 = push_mem_temp == 6'h2; // @[lut_35.scala 6772:30]
  wire  _GEN_11481 = push_mem_temp == 6'h2 ? 1'h0 : 1'h1; // @[lut_35.scala 6772:38 lut_35.scala 216:26 lut_35.scala 6775:16]
  wire  _T_913 = dispatch_reg_3 | clear_3_1; // @[lut_35.scala 6778:33]
  wire [31:0] lo_3 = LUT_mem_MPORT_191_data[31:0]; // @[lut_35.scala 6779:42]
  wire  _T_915 = push_mem_temp == 6'h3; // @[lut_35.scala 6780:30]
  wire  _GEN_11506 = push_mem_temp == 6'h3 ? 1'h0 : 1'h1; // @[lut_35.scala 6780:38 lut_35.scala 216:26 lut_35.scala 6783:16]
  wire  _T_919 = dispatch_reg_4 | clear_4_1; // @[lut_35.scala 6786:33]
  wire [31:0] lo_4 = LUT_mem_MPORT_196_data[31:0]; // @[lut_35.scala 6787:42]
  wire  _T_921 = push_mem_temp == 6'h4; // @[lut_35.scala 6788:30]
  wire  _GEN_11531 = push_mem_temp == 6'h4 ? 1'h0 : 1'h1; // @[lut_35.scala 6788:38 lut_35.scala 216:26 lut_35.scala 6791:16]
  wire  _T_925 = dispatch_reg_5 | clear_5_1; // @[lut_35.scala 6794:33]
  wire [31:0] lo_5 = LUT_mem_MPORT_201_data[31:0]; // @[lut_35.scala 6795:42]
  wire  _T_927 = push_mem_temp == 6'h5; // @[lut_35.scala 6796:30]
  wire  _GEN_11556 = push_mem_temp == 6'h5 ? 1'h0 : 1'h1; // @[lut_35.scala 6796:38 lut_35.scala 216:26 lut_35.scala 6799:16]
  wire  _T_931 = dispatch_reg_6 | clear_6_1; // @[lut_35.scala 6802:33]
  wire [31:0] lo_6 = LUT_mem_MPORT_206_data[31:0]; // @[lut_35.scala 6803:42]
  wire  _T_933 = push_mem_temp == 6'h6; // @[lut_35.scala 6804:30]
  wire  _GEN_11581 = push_mem_temp == 6'h6 ? 1'h0 : 1'h1; // @[lut_35.scala 6804:38 lut_35.scala 216:26 lut_35.scala 6807:16]
  wire  _T_937 = dispatch_reg_7 | clear_7_1; // @[lut_35.scala 6810:33]
  wire [31:0] lo_7 = LUT_mem_MPORT_211_data[31:0]; // @[lut_35.scala 6811:42]
  wire  _T_939 = push_mem_temp == 6'h7; // @[lut_35.scala 6812:30]
  wire  _GEN_11606 = push_mem_temp == 6'h7 ? 1'h0 : 1'h1; // @[lut_35.scala 6812:38 lut_35.scala 216:26 lut_35.scala 6815:16]
  wire  _T_943 = dispatch_reg_8 | clear_8_1; // @[lut_35.scala 6818:33]
  wire [31:0] lo_8 = LUT_mem_MPORT_216_data[31:0]; // @[lut_35.scala 6819:42]
  wire  _T_945 = push_mem_temp == 6'h8; // @[lut_35.scala 6820:30]
  wire  _GEN_11631 = push_mem_temp == 6'h8 ? 1'h0 : 1'h1; // @[lut_35.scala 6820:38 lut_35.scala 216:26 lut_35.scala 6823:16]
  wire  _T_949 = dispatch_reg_9 | clear_9_1; // @[lut_35.scala 6826:33]
  wire [31:0] lo_9 = LUT_mem_MPORT_221_data[31:0]; // @[lut_35.scala 6827:42]
  wire  _T_951 = push_mem_temp == 6'h9; // @[lut_35.scala 6828:30]
  wire  _GEN_11656 = push_mem_temp == 6'h9 ? 1'h0 : 1'h1; // @[lut_35.scala 6828:38 lut_35.scala 216:26 lut_35.scala 6831:16]
  wire  _T_955 = dispatch_reg_10 | clear_10_1; // @[lut_35.scala 6834:34]
  wire [31:0] lo_10 = LUT_mem_MPORT_226_data[31:0]; // @[lut_35.scala 6835:44]
  wire  _T_957 = push_mem_temp == 6'ha; // @[lut_35.scala 6836:30]
  wire  _GEN_11681 = push_mem_temp == 6'ha ? 1'h0 : 1'h1; // @[lut_35.scala 6836:39 lut_35.scala 216:26 lut_35.scala 6839:16]
  wire  _T_961 = dispatch_reg_11 | clear_11_1; // @[lut_35.scala 6842:34]
  wire [31:0] lo_11 = LUT_mem_MPORT_231_data[31:0]; // @[lut_35.scala 6843:44]
  wire  _T_963 = push_mem_temp == 6'hb; // @[lut_35.scala 6844:30]
  wire  _GEN_11706 = push_mem_temp == 6'hb ? 1'h0 : 1'h1; // @[lut_35.scala 6844:39 lut_35.scala 216:26 lut_35.scala 6847:16]
  wire  _T_967 = dispatch_reg_12 | clear_12_1; // @[lut_35.scala 6850:34]
  wire [31:0] lo_12 = LUT_mem_MPORT_236_data[31:0]; // @[lut_35.scala 6851:44]
  wire  _T_969 = push_mem_temp == 6'hc; // @[lut_35.scala 6852:30]
  wire  _GEN_11731 = push_mem_temp == 6'hc ? 1'h0 : 1'h1; // @[lut_35.scala 6852:39 lut_35.scala 216:26 lut_35.scala 6855:16]
  wire  _T_973 = dispatch_reg_13 | clear_13_1; // @[lut_35.scala 6858:34]
  wire [31:0] lo_13 = LUT_mem_MPORT_241_data[31:0]; // @[lut_35.scala 6859:44]
  wire  _T_975 = push_mem_temp == 6'hd; // @[lut_35.scala 6860:30]
  wire  _GEN_11756 = push_mem_temp == 6'hd ? 1'h0 : 1'h1; // @[lut_35.scala 6860:39 lut_35.scala 216:26 lut_35.scala 6863:16]
  wire  _T_979 = dispatch_reg_14 | clear_14_1; // @[lut_35.scala 6866:34]
  wire [31:0] lo_14 = LUT_mem_MPORT_246_data[31:0]; // @[lut_35.scala 6867:44]
  wire  _T_981 = push_mem_temp == 6'he; // @[lut_35.scala 6868:30]
  wire  _GEN_11781 = push_mem_temp == 6'he ? 1'h0 : 1'h1; // @[lut_35.scala 6868:39 lut_35.scala 216:26 lut_35.scala 6871:16]
  wire  _T_985 = dispatch_reg_15 | clear_15_1; // @[lut_35.scala 6874:34]
  wire [31:0] lo_15 = LUT_mem_MPORT_251_data[31:0]; // @[lut_35.scala 6875:44]
  wire  _T_987 = push_mem_temp == 6'hf; // @[lut_35.scala 6876:30]
  wire  _GEN_11806 = push_mem_temp == 6'hf ? 1'h0 : 1'h1; // @[lut_35.scala 6876:39 lut_35.scala 216:26 lut_35.scala 6879:16]
  wire  _T_991 = dispatch_reg_16 | clear_16_1; // @[lut_35.scala 6882:34]
  wire [31:0] lo_16 = LUT_mem_MPORT_256_data[31:0]; // @[lut_35.scala 6883:44]
  wire  _T_993 = push_mem_temp == 6'h10; // @[lut_35.scala 6884:30]
  wire  _GEN_11831 = push_mem_temp == 6'h10 ? 1'h0 : 1'h1; // @[lut_35.scala 6884:39 lut_35.scala 216:26 lut_35.scala 6887:16]
  wire  _T_997 = dispatch_reg_17 | clear_17_1; // @[lut_35.scala 6890:34]
  wire [31:0] lo_17 = LUT_mem_MPORT_261_data[31:0]; // @[lut_35.scala 6891:44]
  wire  _T_999 = push_mem_temp == 6'h11; // @[lut_35.scala 6892:30]
  wire  _GEN_11856 = push_mem_temp == 6'h11 ? 1'h0 : 1'h1; // @[lut_35.scala 6892:39 lut_35.scala 216:26 lut_35.scala 6895:16]
  wire  _T_1003 = dispatch_reg_18 | clear_18_1; // @[lut_35.scala 6898:34]
  wire [31:0] lo_18 = LUT_mem_MPORT_266_data[31:0]; // @[lut_35.scala 6899:44]
  wire  _T_1005 = push_mem_temp == 6'h12; // @[lut_35.scala 6900:30]
  wire  _GEN_11881 = push_mem_temp == 6'h12 ? 1'h0 : 1'h1; // @[lut_35.scala 6900:39 lut_35.scala 216:26 lut_35.scala 6903:16]
  wire  _T_1009 = dispatch_reg_19 | clear_19_1; // @[lut_35.scala 6906:34]
  wire [31:0] lo_19 = LUT_mem_MPORT_271_data[31:0]; // @[lut_35.scala 6907:44]
  wire  _T_1011 = push_mem_temp == 6'h13; // @[lut_35.scala 6908:30]
  wire  _GEN_11906 = push_mem_temp == 6'h13 ? 1'h0 : 1'h1; // @[lut_35.scala 6908:39 lut_35.scala 216:26 lut_35.scala 6911:16]
  wire  _T_1015 = dispatch_reg_20 | clear_20_1; // @[lut_35.scala 6914:34]
  wire [31:0] lo_20 = LUT_mem_MPORT_276_data[31:0]; // @[lut_35.scala 6915:44]
  wire  _T_1017 = push_mem_temp == 6'h14; // @[lut_35.scala 6916:30]
  wire  _GEN_11931 = push_mem_temp == 6'h14 ? 1'h0 : 1'h1; // @[lut_35.scala 6916:39 lut_35.scala 216:26 lut_35.scala 6919:16]
  wire  _T_1021 = dispatch_reg_21 | clear_21_1; // @[lut_35.scala 6922:34]
  wire [31:0] lo_21 = LUT_mem_MPORT_281_data[31:0]; // @[lut_35.scala 6923:44]
  wire  _T_1023 = push_mem_temp == 6'h15; // @[lut_35.scala 6924:30]
  wire  _GEN_11956 = push_mem_temp == 6'h15 ? 1'h0 : 1'h1; // @[lut_35.scala 6924:39 lut_35.scala 216:26 lut_35.scala 6927:16]
  wire  _T_1027 = dispatch_reg_22 | clear_22_1; // @[lut_35.scala 6930:34]
  wire [31:0] lo_22 = LUT_mem_MPORT_286_data[31:0]; // @[lut_35.scala 6931:44]
  wire  _T_1029 = push_mem_temp == 6'h16; // @[lut_35.scala 6932:30]
  wire  _GEN_11981 = push_mem_temp == 6'h16 ? 1'h0 : 1'h1; // @[lut_35.scala 6932:39 lut_35.scala 216:26 lut_35.scala 6935:16]
  wire  _T_1033 = dispatch_reg_23 | clear_23_1; // @[lut_35.scala 6938:34]
  wire [31:0] lo_23 = LUT_mem_MPORT_291_data[31:0]; // @[lut_35.scala 6939:44]
  wire  _T_1035 = push_mem_temp == 6'h17; // @[lut_35.scala 6940:30]
  wire  _GEN_12006 = push_mem_temp == 6'h17 ? 1'h0 : 1'h1; // @[lut_35.scala 6940:39 lut_35.scala 216:26 lut_35.scala 6943:16]
  wire  _T_1039 = dispatch_reg_24 | clear_24_1; // @[lut_35.scala 6946:34]
  wire [31:0] lo_24 = LUT_mem_MPORT_296_data[31:0]; // @[lut_35.scala 6947:44]
  wire  _T_1041 = push_mem_temp == 6'h18; // @[lut_35.scala 6948:30]
  wire  _GEN_12031 = push_mem_temp == 6'h18 ? 1'h0 : 1'h1; // @[lut_35.scala 6948:39 lut_35.scala 216:26 lut_35.scala 6951:16]
  wire  _T_1045 = dispatch_reg_25 | clear_25_1; // @[lut_35.scala 6954:34]
  wire [31:0] lo_25 = LUT_mem_MPORT_301_data[31:0]; // @[lut_35.scala 6955:44]
  wire  _T_1047 = push_mem_temp == 6'h19; // @[lut_35.scala 6956:30]
  wire  _GEN_12056 = push_mem_temp == 6'h19 ? 1'h0 : 1'h1; // @[lut_35.scala 6956:39 lut_35.scala 216:26 lut_35.scala 6959:16]
  wire  _T_1051 = dispatch_reg_26 | clear_26_1; // @[lut_35.scala 6962:34]
  wire [31:0] lo_26 = LUT_mem_MPORT_306_data[31:0]; // @[lut_35.scala 6963:44]
  wire  _T_1053 = push_mem_temp == 6'h1a; // @[lut_35.scala 6964:30]
  wire  _GEN_12081 = push_mem_temp == 6'h1a ? 1'h0 : 1'h1; // @[lut_35.scala 6964:39 lut_35.scala 216:26 lut_35.scala 6967:16]
  wire  _T_1057 = dispatch_reg_27 | clear_27_1; // @[lut_35.scala 6970:34]
  wire [31:0] lo_27 = LUT_mem_MPORT_311_data[31:0]; // @[lut_35.scala 6971:44]
  wire  _T_1059 = push_mem_temp == 6'h1b; // @[lut_35.scala 6972:30]
  wire  _GEN_12106 = push_mem_temp == 6'h1b ? 1'h0 : 1'h1; // @[lut_35.scala 6972:39 lut_35.scala 216:26 lut_35.scala 6975:16]
  wire  _T_1063 = dispatch_reg_28 | clear_28_1; // @[lut_35.scala 6978:34]
  wire [31:0] lo_28 = LUT_mem_MPORT_316_data[31:0]; // @[lut_35.scala 6979:44]
  wire  _T_1065 = push_mem_temp == 6'h1c; // @[lut_35.scala 6980:30]
  wire  _GEN_12131 = push_mem_temp == 6'h1c ? 1'h0 : 1'h1; // @[lut_35.scala 6980:39 lut_35.scala 216:26 lut_35.scala 6983:16]
  wire  _T_1069 = dispatch_reg_29 | clear_29_1; // @[lut_35.scala 6986:34]
  wire [31:0] lo_29 = LUT_mem_MPORT_321_data[31:0]; // @[lut_35.scala 6987:44]
  wire  _T_1071 = push_mem_temp == 6'h1d; // @[lut_35.scala 6988:30]
  wire  _GEN_12156 = push_mem_temp == 6'h1d ? 1'h0 : 1'h1; // @[lut_35.scala 6988:39 lut_35.scala 216:26 lut_35.scala 6991:16]
  wire  _T_1075 = dispatch_reg_30 | clear_30_1; // @[lut_35.scala 6994:36]
  wire [31:0] lo_30 = LUT_mem_MPORT_326_data[31:0]; // @[lut_35.scala 6995:44]
  wire  _T_1077 = push_mem_temp == 6'h1e; // @[lut_35.scala 6996:30]
  wire  _GEN_12181 = push_mem_temp == 6'h1e ? 1'h0 : 1'h1; // @[lut_35.scala 6996:39 lut_35.scala 216:26 lut_35.scala 6999:16]
  wire  _T_1081 = dispatch_reg_31 | clear_31_1; // @[lut_35.scala 7002:34]
  wire [31:0] lo_31 = LUT_mem_MPORT_331_data[31:0]; // @[lut_35.scala 7003:44]
  wire  _T_1083 = push_mem_temp == 6'h1f; // @[lut_35.scala 7004:30]
  wire  _GEN_12206 = push_mem_temp == 6'h1f ? 1'h0 : 1'h1; // @[lut_35.scala 7004:39 lut_35.scala 216:26 lut_35.scala 7007:16]
  wire  _T_1087 = dispatch_reg_32 | clear_32_1; // @[lut_35.scala 7010:34]
  wire [31:0] lo_32 = LUT_mem_MPORT_336_data[31:0]; // @[lut_35.scala 7011:44]
  wire  _T_1089 = push_mem_temp == 6'h20; // @[lut_35.scala 7012:30]
  wire  _GEN_12231 = push_mem_temp == 6'h20 ? 1'h0 : 1'h1; // @[lut_35.scala 7012:39 lut_35.scala 216:26 lut_35.scala 7015:16]
  wire  _T_1093 = dispatch_reg_33 | clear_33_1; // @[lut_35.scala 7018:34]
  wire [31:0] lo_33 = LUT_mem_MPORT_341_data[31:0]; // @[lut_35.scala 7019:44]
  wire  _T_1095 = push_mem_temp == 6'h21; // @[lut_35.scala 7020:30]
  wire  _GEN_12256 = push_mem_temp == 6'h21 ? 1'h0 : 1'h1; // @[lut_35.scala 7020:39 lut_35.scala 216:26 lut_35.scala 7023:16]
  wire  _T_1099 = dispatch_reg_34 | clear_34_1; // @[lut_35.scala 7026:34]
  wire [31:0] lo_34 = LUT_mem_MPORT_346_data[31:0]; // @[lut_35.scala 7027:44]
  wire  _T_1101 = push_mem_temp == 6'h22; // @[lut_35.scala 7028:30]
  wire  _GEN_12281 = push_mem_temp == 6'h22 ? 1'h0 : 1'h1; // @[lut_35.scala 7028:39 lut_35.scala 216:26 lut_35.scala 7031:16]
  assign LUT_mem_MPORT_addr = 6'h0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_data = LUT_mem[LUT_mem_MPORT_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_data = LUT_mem_MPORT_addr >= 6'h23 ? _RAND_1[32:0] : LUT_mem[LUT_mem_MPORT_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_1_addr = 6'h1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_1_data = LUT_mem[LUT_mem_MPORT_1_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_1_data = LUT_mem_MPORT_1_addr >= 6'h23 ? _RAND_2[32:0] : LUT_mem[LUT_mem_MPORT_1_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_2_addr = 6'h2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_2_data = LUT_mem[LUT_mem_MPORT_2_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_2_data = LUT_mem_MPORT_2_addr >= 6'h23 ? _RAND_3[32:0] : LUT_mem[LUT_mem_MPORT_2_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_3_addr = 6'h3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_3_data = LUT_mem[LUT_mem_MPORT_3_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_3_data = LUT_mem_MPORT_3_addr >= 6'h23 ? _RAND_4[32:0] : LUT_mem[LUT_mem_MPORT_3_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_4_addr = 6'h4;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_4_data = LUT_mem[LUT_mem_MPORT_4_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_4_data = LUT_mem_MPORT_4_addr >= 6'h23 ? _RAND_5[32:0] : LUT_mem[LUT_mem_MPORT_4_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_5_addr = 6'h5;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_5_data = LUT_mem[LUT_mem_MPORT_5_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_5_data = LUT_mem_MPORT_5_addr >= 6'h23 ? _RAND_6[32:0] : LUT_mem[LUT_mem_MPORT_5_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_6_addr = 6'h6;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_6_data = LUT_mem[LUT_mem_MPORT_6_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_6_data = LUT_mem_MPORT_6_addr >= 6'h23 ? _RAND_7[32:0] : LUT_mem[LUT_mem_MPORT_6_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_7_addr = 6'h7;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_7_data = LUT_mem[LUT_mem_MPORT_7_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_7_data = LUT_mem_MPORT_7_addr >= 6'h23 ? _RAND_8[32:0] : LUT_mem[LUT_mem_MPORT_7_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_8_addr = 6'h8;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_8_data = LUT_mem[LUT_mem_MPORT_8_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_8_data = LUT_mem_MPORT_8_addr >= 6'h23 ? _RAND_9[32:0] : LUT_mem[LUT_mem_MPORT_8_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_9_addr = 6'h9;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_9_data = LUT_mem[LUT_mem_MPORT_9_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_9_data = LUT_mem_MPORT_9_addr >= 6'h23 ? _RAND_10[32:0] : LUT_mem[LUT_mem_MPORT_9_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_10_addr = 6'ha;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_10_data = LUT_mem[LUT_mem_MPORT_10_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_10_data = LUT_mem_MPORT_10_addr >= 6'h23 ? _RAND_11[32:0] : LUT_mem[LUT_mem_MPORT_10_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_11_addr = 6'hb;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_11_data = LUT_mem[LUT_mem_MPORT_11_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_11_data = LUT_mem_MPORT_11_addr >= 6'h23 ? _RAND_12[32:0] : LUT_mem[LUT_mem_MPORT_11_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_12_addr = 6'hc;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_12_data = LUT_mem[LUT_mem_MPORT_12_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_12_data = LUT_mem_MPORT_12_addr >= 6'h23 ? _RAND_13[32:0] : LUT_mem[LUT_mem_MPORT_12_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_13_addr = 6'hd;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_13_data = LUT_mem[LUT_mem_MPORT_13_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_13_data = LUT_mem_MPORT_13_addr >= 6'h23 ? _RAND_14[32:0] : LUT_mem[LUT_mem_MPORT_13_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_14_addr = 6'he;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_14_data = LUT_mem[LUT_mem_MPORT_14_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_14_data = LUT_mem_MPORT_14_addr >= 6'h23 ? _RAND_15[32:0] : LUT_mem[LUT_mem_MPORT_14_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_15_addr = 6'hf;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_15_data = LUT_mem[LUT_mem_MPORT_15_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_15_data = LUT_mem_MPORT_15_addr >= 6'h23 ? _RAND_16[32:0] : LUT_mem[LUT_mem_MPORT_15_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_16_addr = 6'h10;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_16_data = LUT_mem[LUT_mem_MPORT_16_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_16_data = LUT_mem_MPORT_16_addr >= 6'h23 ? _RAND_17[32:0] : LUT_mem[LUT_mem_MPORT_16_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_17_addr = 6'h11;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_17_data = LUT_mem[LUT_mem_MPORT_17_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_17_data = LUT_mem_MPORT_17_addr >= 6'h23 ? _RAND_18[32:0] : LUT_mem[LUT_mem_MPORT_17_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_18_addr = 6'h12;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_18_data = LUT_mem[LUT_mem_MPORT_18_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_18_data = LUT_mem_MPORT_18_addr >= 6'h23 ? _RAND_19[32:0] : LUT_mem[LUT_mem_MPORT_18_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_19_addr = 6'h13;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_19_data = LUT_mem[LUT_mem_MPORT_19_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_19_data = LUT_mem_MPORT_19_addr >= 6'h23 ? _RAND_20[32:0] : LUT_mem[LUT_mem_MPORT_19_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_20_addr = 6'h14;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_20_data = LUT_mem[LUT_mem_MPORT_20_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_20_data = LUT_mem_MPORT_20_addr >= 6'h23 ? _RAND_21[32:0] : LUT_mem[LUT_mem_MPORT_20_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_21_addr = 6'h15;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_21_data = LUT_mem[LUT_mem_MPORT_21_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_21_data = LUT_mem_MPORT_21_addr >= 6'h23 ? _RAND_22[32:0] : LUT_mem[LUT_mem_MPORT_21_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_22_addr = 6'h16;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_22_data = LUT_mem[LUT_mem_MPORT_22_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_22_data = LUT_mem_MPORT_22_addr >= 6'h23 ? _RAND_23[32:0] : LUT_mem[LUT_mem_MPORT_22_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_23_addr = 6'h17;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_23_data = LUT_mem[LUT_mem_MPORT_23_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_23_data = LUT_mem_MPORT_23_addr >= 6'h23 ? _RAND_24[32:0] : LUT_mem[LUT_mem_MPORT_23_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_24_addr = 6'h18;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_24_data = LUT_mem[LUT_mem_MPORT_24_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_24_data = LUT_mem_MPORT_24_addr >= 6'h23 ? _RAND_25[32:0] : LUT_mem[LUT_mem_MPORT_24_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_25_addr = 6'h19;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_25_data = LUT_mem[LUT_mem_MPORT_25_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_25_data = LUT_mem_MPORT_25_addr >= 6'h23 ? _RAND_26[32:0] : LUT_mem[LUT_mem_MPORT_25_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_26_addr = 6'h1a;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_26_data = LUT_mem[LUT_mem_MPORT_26_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_26_data = LUT_mem_MPORT_26_addr >= 6'h23 ? _RAND_27[32:0] : LUT_mem[LUT_mem_MPORT_26_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_27_addr = 6'h1b;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_27_data = LUT_mem[LUT_mem_MPORT_27_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_27_data = LUT_mem_MPORT_27_addr >= 6'h23 ? _RAND_28[32:0] : LUT_mem[LUT_mem_MPORT_27_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_28_addr = 6'h1c;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_28_data = LUT_mem[LUT_mem_MPORT_28_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_28_data = LUT_mem_MPORT_28_addr >= 6'h23 ? _RAND_29[32:0] : LUT_mem[LUT_mem_MPORT_28_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_29_addr = 6'h1d;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_29_data = LUT_mem[LUT_mem_MPORT_29_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_29_data = LUT_mem_MPORT_29_addr >= 6'h23 ? _RAND_30[32:0] : LUT_mem[LUT_mem_MPORT_29_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_30_addr = 6'h1e;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_30_data = LUT_mem[LUT_mem_MPORT_30_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_30_data = LUT_mem_MPORT_30_addr >= 6'h23 ? _RAND_31[32:0] : LUT_mem[LUT_mem_MPORT_30_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_31_addr = 6'h1f;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_31_data = LUT_mem[LUT_mem_MPORT_31_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_31_data = LUT_mem_MPORT_31_addr >= 6'h23 ? _RAND_32[32:0] : LUT_mem[LUT_mem_MPORT_31_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_32_addr = 6'h20;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_32_data = LUT_mem[LUT_mem_MPORT_32_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_32_data = LUT_mem_MPORT_32_addr >= 6'h23 ? _RAND_33[32:0] : LUT_mem[LUT_mem_MPORT_32_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_33_addr = 6'h21;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_33_data = LUT_mem[LUT_mem_MPORT_33_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_33_data = LUT_mem_MPORT_33_addr >= 6'h23 ? _RAND_34[32:0] : LUT_mem[LUT_mem_MPORT_33_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_34_addr = 6'h22;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_34_data = LUT_mem[LUT_mem_MPORT_34_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_34_data = LUT_mem_MPORT_34_addr >= 6'h23 ? _RAND_35[32:0] : LUT_mem[LUT_mem_MPORT_34_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_35_addr = 6'h0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_35_data = LUT_mem[LUT_mem_MPORT_35_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_35_data = LUT_mem_MPORT_35_addr >= 6'h23 ? _RAND_36[32:0] : LUT_mem[LUT_mem_MPORT_35_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_36_addr = 6'h1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_36_data = LUT_mem[LUT_mem_MPORT_36_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_36_data = LUT_mem_MPORT_36_addr >= 6'h23 ? _RAND_37[32:0] : LUT_mem[LUT_mem_MPORT_36_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_37_addr = 6'h2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_37_data = LUT_mem[LUT_mem_MPORT_37_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_37_data = LUT_mem_MPORT_37_addr >= 6'h23 ? _RAND_38[32:0] : LUT_mem[LUT_mem_MPORT_37_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_38_addr = 6'h3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_38_data = LUT_mem[LUT_mem_MPORT_38_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_38_data = LUT_mem_MPORT_38_addr >= 6'h23 ? _RAND_39[32:0] : LUT_mem[LUT_mem_MPORT_38_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_39_addr = 6'h4;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_39_data = LUT_mem[LUT_mem_MPORT_39_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_39_data = LUT_mem_MPORT_39_addr >= 6'h23 ? _RAND_40[32:0] : LUT_mem[LUT_mem_MPORT_39_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_40_addr = 6'h5;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_40_data = LUT_mem[LUT_mem_MPORT_40_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_40_data = LUT_mem_MPORT_40_addr >= 6'h23 ? _RAND_41[32:0] : LUT_mem[LUT_mem_MPORT_40_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_41_addr = 6'h6;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_41_data = LUT_mem[LUT_mem_MPORT_41_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_41_data = LUT_mem_MPORT_41_addr >= 6'h23 ? _RAND_42[32:0] : LUT_mem[LUT_mem_MPORT_41_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_42_addr = 6'h7;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_42_data = LUT_mem[LUT_mem_MPORT_42_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_42_data = LUT_mem_MPORT_42_addr >= 6'h23 ? _RAND_43[32:0] : LUT_mem[LUT_mem_MPORT_42_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_43_addr = 6'h8;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_43_data = LUT_mem[LUT_mem_MPORT_43_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_43_data = LUT_mem_MPORT_43_addr >= 6'h23 ? _RAND_44[32:0] : LUT_mem[LUT_mem_MPORT_43_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_44_addr = 6'h9;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_44_data = LUT_mem[LUT_mem_MPORT_44_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_44_data = LUT_mem_MPORT_44_addr >= 6'h23 ? _RAND_45[32:0] : LUT_mem[LUT_mem_MPORT_44_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_45_addr = 6'ha;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_45_data = LUT_mem[LUT_mem_MPORT_45_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_45_data = LUT_mem_MPORT_45_addr >= 6'h23 ? _RAND_46[32:0] : LUT_mem[LUT_mem_MPORT_45_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_46_addr = 6'hb;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_46_data = LUT_mem[LUT_mem_MPORT_46_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_46_data = LUT_mem_MPORT_46_addr >= 6'h23 ? _RAND_47[32:0] : LUT_mem[LUT_mem_MPORT_46_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_47_addr = 6'hc;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_47_data = LUT_mem[LUT_mem_MPORT_47_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_47_data = LUT_mem_MPORT_47_addr >= 6'h23 ? _RAND_48[32:0] : LUT_mem[LUT_mem_MPORT_47_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_48_addr = 6'hd;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_48_data = LUT_mem[LUT_mem_MPORT_48_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_48_data = LUT_mem_MPORT_48_addr >= 6'h23 ? _RAND_49[32:0] : LUT_mem[LUT_mem_MPORT_48_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_49_addr = 6'he;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_49_data = LUT_mem[LUT_mem_MPORT_49_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_49_data = LUT_mem_MPORT_49_addr >= 6'h23 ? _RAND_50[32:0] : LUT_mem[LUT_mem_MPORT_49_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_50_addr = 6'hf;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_50_data = LUT_mem[LUT_mem_MPORT_50_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_50_data = LUT_mem_MPORT_50_addr >= 6'h23 ? _RAND_51[32:0] : LUT_mem[LUT_mem_MPORT_50_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_51_addr = 6'h10;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_51_data = LUT_mem[LUT_mem_MPORT_51_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_51_data = LUT_mem_MPORT_51_addr >= 6'h23 ? _RAND_52[32:0] : LUT_mem[LUT_mem_MPORT_51_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_52_addr = 6'h11;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_52_data = LUT_mem[LUT_mem_MPORT_52_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_52_data = LUT_mem_MPORT_52_addr >= 6'h23 ? _RAND_53[32:0] : LUT_mem[LUT_mem_MPORT_52_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_53_addr = 6'h12;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_53_data = LUT_mem[LUT_mem_MPORT_53_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_53_data = LUT_mem_MPORT_53_addr >= 6'h23 ? _RAND_54[32:0] : LUT_mem[LUT_mem_MPORT_53_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_54_addr = 6'h13;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_54_data = LUT_mem[LUT_mem_MPORT_54_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_54_data = LUT_mem_MPORT_54_addr >= 6'h23 ? _RAND_55[32:0] : LUT_mem[LUT_mem_MPORT_54_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_55_addr = 6'h14;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_55_data = LUT_mem[LUT_mem_MPORT_55_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_55_data = LUT_mem_MPORT_55_addr >= 6'h23 ? _RAND_56[32:0] : LUT_mem[LUT_mem_MPORT_55_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_56_addr = 6'h15;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_56_data = LUT_mem[LUT_mem_MPORT_56_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_56_data = LUT_mem_MPORT_56_addr >= 6'h23 ? _RAND_57[32:0] : LUT_mem[LUT_mem_MPORT_56_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_57_addr = 6'h16;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_57_data = LUT_mem[LUT_mem_MPORT_57_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_57_data = LUT_mem_MPORT_57_addr >= 6'h23 ? _RAND_58[32:0] : LUT_mem[LUT_mem_MPORT_57_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_58_addr = 6'h17;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_58_data = LUT_mem[LUT_mem_MPORT_58_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_58_data = LUT_mem_MPORT_58_addr >= 6'h23 ? _RAND_59[32:0] : LUT_mem[LUT_mem_MPORT_58_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_59_addr = 6'h18;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_59_data = LUT_mem[LUT_mem_MPORT_59_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_59_data = LUT_mem_MPORT_59_addr >= 6'h23 ? _RAND_60[32:0] : LUT_mem[LUT_mem_MPORT_59_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_60_addr = 6'h19;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_60_data = LUT_mem[LUT_mem_MPORT_60_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_60_data = LUT_mem_MPORT_60_addr >= 6'h23 ? _RAND_61[32:0] : LUT_mem[LUT_mem_MPORT_60_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_61_addr = 6'h1a;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_61_data = LUT_mem[LUT_mem_MPORT_61_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_61_data = LUT_mem_MPORT_61_addr >= 6'h23 ? _RAND_62[32:0] : LUT_mem[LUT_mem_MPORT_61_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_62_addr = 6'h1b;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_62_data = LUT_mem[LUT_mem_MPORT_62_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_62_data = LUT_mem_MPORT_62_addr >= 6'h23 ? _RAND_63[32:0] : LUT_mem[LUT_mem_MPORT_62_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_63_addr = 6'h1c;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_63_data = LUT_mem[LUT_mem_MPORT_63_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_63_data = LUT_mem_MPORT_63_addr >= 6'h23 ? _RAND_64[32:0] : LUT_mem[LUT_mem_MPORT_63_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_64_addr = 6'h1d;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_64_data = LUT_mem[LUT_mem_MPORT_64_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_64_data = LUT_mem_MPORT_64_addr >= 6'h23 ? _RAND_65[32:0] : LUT_mem[LUT_mem_MPORT_64_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_65_addr = 6'h1e;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_65_data = LUT_mem[LUT_mem_MPORT_65_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_65_data = LUT_mem_MPORT_65_addr >= 6'h23 ? _RAND_66[32:0] : LUT_mem[LUT_mem_MPORT_65_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_66_addr = 6'h1f;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_66_data = LUT_mem[LUT_mem_MPORT_66_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_66_data = LUT_mem_MPORT_66_addr >= 6'h23 ? _RAND_67[32:0] : LUT_mem[LUT_mem_MPORT_66_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_67_addr = 6'h20;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_67_data = LUT_mem[LUT_mem_MPORT_67_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_67_data = LUT_mem_MPORT_67_addr >= 6'h23 ? _RAND_68[32:0] : LUT_mem[LUT_mem_MPORT_67_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_68_addr = 6'h21;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_68_data = LUT_mem[LUT_mem_MPORT_68_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_68_data = LUT_mem_MPORT_68_addr >= 6'h23 ? _RAND_69[32:0] : LUT_mem[LUT_mem_MPORT_68_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_69_addr = 6'h22;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_69_data = LUT_mem[LUT_mem_MPORT_69_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_69_data = LUT_mem_MPORT_69_addr >= 6'h23 ? _RAND_70[32:0] : LUT_mem[LUT_mem_MPORT_69_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_70_addr = 6'h0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_70_data = LUT_mem[LUT_mem_MPORT_70_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_70_data = LUT_mem_MPORT_70_addr >= 6'h23 ? _RAND_71[32:0] : LUT_mem[LUT_mem_MPORT_70_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_71_addr = 6'h1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_71_data = LUT_mem[LUT_mem_MPORT_71_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_71_data = LUT_mem_MPORT_71_addr >= 6'h23 ? _RAND_72[32:0] : LUT_mem[LUT_mem_MPORT_71_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_72_addr = 6'h2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_72_data = LUT_mem[LUT_mem_MPORT_72_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_72_data = LUT_mem_MPORT_72_addr >= 6'h23 ? _RAND_73[32:0] : LUT_mem[LUT_mem_MPORT_72_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_73_addr = 6'h3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_73_data = LUT_mem[LUT_mem_MPORT_73_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_73_data = LUT_mem_MPORT_73_addr >= 6'h23 ? _RAND_74[32:0] : LUT_mem[LUT_mem_MPORT_73_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_74_addr = 6'h4;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_74_data = LUT_mem[LUT_mem_MPORT_74_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_74_data = LUT_mem_MPORT_74_addr >= 6'h23 ? _RAND_75[32:0] : LUT_mem[LUT_mem_MPORT_74_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_75_addr = 6'h5;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_75_data = LUT_mem[LUT_mem_MPORT_75_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_75_data = LUT_mem_MPORT_75_addr >= 6'h23 ? _RAND_76[32:0] : LUT_mem[LUT_mem_MPORT_75_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_76_addr = 6'h6;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_76_data = LUT_mem[LUT_mem_MPORT_76_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_76_data = LUT_mem_MPORT_76_addr >= 6'h23 ? _RAND_77[32:0] : LUT_mem[LUT_mem_MPORT_76_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_77_addr = 6'h7;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_77_data = LUT_mem[LUT_mem_MPORT_77_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_77_data = LUT_mem_MPORT_77_addr >= 6'h23 ? _RAND_78[32:0] : LUT_mem[LUT_mem_MPORT_77_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_78_addr = 6'h8;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_78_data = LUT_mem[LUT_mem_MPORT_78_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_78_data = LUT_mem_MPORT_78_addr >= 6'h23 ? _RAND_79[32:0] : LUT_mem[LUT_mem_MPORT_78_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_79_addr = 6'h9;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_79_data = LUT_mem[LUT_mem_MPORT_79_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_79_data = LUT_mem_MPORT_79_addr >= 6'h23 ? _RAND_80[32:0] : LUT_mem[LUT_mem_MPORT_79_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_80_addr = 6'ha;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_80_data = LUT_mem[LUT_mem_MPORT_80_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_80_data = LUT_mem_MPORT_80_addr >= 6'h23 ? _RAND_81[32:0] : LUT_mem[LUT_mem_MPORT_80_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_81_addr = 6'hb;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_81_data = LUT_mem[LUT_mem_MPORT_81_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_81_data = LUT_mem_MPORT_81_addr >= 6'h23 ? _RAND_82[32:0] : LUT_mem[LUT_mem_MPORT_81_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_82_addr = 6'hc;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_82_data = LUT_mem[LUT_mem_MPORT_82_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_82_data = LUT_mem_MPORT_82_addr >= 6'h23 ? _RAND_83[32:0] : LUT_mem[LUT_mem_MPORT_82_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_83_addr = 6'hd;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_83_data = LUT_mem[LUT_mem_MPORT_83_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_83_data = LUT_mem_MPORT_83_addr >= 6'h23 ? _RAND_84[32:0] : LUT_mem[LUT_mem_MPORT_83_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_84_addr = 6'he;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_84_data = LUT_mem[LUT_mem_MPORT_84_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_84_data = LUT_mem_MPORT_84_addr >= 6'h23 ? _RAND_85[32:0] : LUT_mem[LUT_mem_MPORT_84_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_85_addr = 6'hf;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_85_data = LUT_mem[LUT_mem_MPORT_85_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_85_data = LUT_mem_MPORT_85_addr >= 6'h23 ? _RAND_86[32:0] : LUT_mem[LUT_mem_MPORT_85_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_86_addr = 6'h10;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_86_data = LUT_mem[LUT_mem_MPORT_86_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_86_data = LUT_mem_MPORT_86_addr >= 6'h23 ? _RAND_87[32:0] : LUT_mem[LUT_mem_MPORT_86_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_87_addr = 6'h11;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_87_data = LUT_mem[LUT_mem_MPORT_87_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_87_data = LUT_mem_MPORT_87_addr >= 6'h23 ? _RAND_88[32:0] : LUT_mem[LUT_mem_MPORT_87_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_88_addr = 6'h12;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_88_data = LUT_mem[LUT_mem_MPORT_88_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_88_data = LUT_mem_MPORT_88_addr >= 6'h23 ? _RAND_89[32:0] : LUT_mem[LUT_mem_MPORT_88_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_89_addr = 6'h13;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_89_data = LUT_mem[LUT_mem_MPORT_89_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_89_data = LUT_mem_MPORT_89_addr >= 6'h23 ? _RAND_90[32:0] : LUT_mem[LUT_mem_MPORT_89_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_90_addr = 6'h14;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_90_data = LUT_mem[LUT_mem_MPORT_90_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_90_data = LUT_mem_MPORT_90_addr >= 6'h23 ? _RAND_91[32:0] : LUT_mem[LUT_mem_MPORT_90_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_91_addr = 6'h15;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_91_data = LUT_mem[LUT_mem_MPORT_91_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_91_data = LUT_mem_MPORT_91_addr >= 6'h23 ? _RAND_92[32:0] : LUT_mem[LUT_mem_MPORT_91_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_92_addr = 6'h16;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_92_data = LUT_mem[LUT_mem_MPORT_92_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_92_data = LUT_mem_MPORT_92_addr >= 6'h23 ? _RAND_93[32:0] : LUT_mem[LUT_mem_MPORT_92_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_93_addr = 6'h17;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_93_data = LUT_mem[LUT_mem_MPORT_93_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_93_data = LUT_mem_MPORT_93_addr >= 6'h23 ? _RAND_94[32:0] : LUT_mem[LUT_mem_MPORT_93_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_94_addr = 6'h18;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_94_data = LUT_mem[LUT_mem_MPORT_94_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_94_data = LUT_mem_MPORT_94_addr >= 6'h23 ? _RAND_95[32:0] : LUT_mem[LUT_mem_MPORT_94_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_95_addr = 6'h19;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_95_data = LUT_mem[LUT_mem_MPORT_95_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_95_data = LUT_mem_MPORT_95_addr >= 6'h23 ? _RAND_96[32:0] : LUT_mem[LUT_mem_MPORT_95_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_96_addr = 6'h1a;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_96_data = LUT_mem[LUT_mem_MPORT_96_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_96_data = LUT_mem_MPORT_96_addr >= 6'h23 ? _RAND_97[32:0] : LUT_mem[LUT_mem_MPORT_96_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_97_addr = 6'h1b;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_97_data = LUT_mem[LUT_mem_MPORT_97_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_97_data = LUT_mem_MPORT_97_addr >= 6'h23 ? _RAND_98[32:0] : LUT_mem[LUT_mem_MPORT_97_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_98_addr = 6'h1c;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_98_data = LUT_mem[LUT_mem_MPORT_98_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_98_data = LUT_mem_MPORT_98_addr >= 6'h23 ? _RAND_99[32:0] : LUT_mem[LUT_mem_MPORT_98_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_99_addr = 6'h1d;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_99_data = LUT_mem[LUT_mem_MPORT_99_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_99_data = LUT_mem_MPORT_99_addr >= 6'h23 ? _RAND_100[32:0] : LUT_mem[LUT_mem_MPORT_99_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_100_addr = 6'h1e;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_100_data = LUT_mem[LUT_mem_MPORT_100_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_100_data = LUT_mem_MPORT_100_addr >= 6'h23 ? _RAND_101[32:0] : LUT_mem[LUT_mem_MPORT_100_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_101_addr = 6'h1f;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_101_data = LUT_mem[LUT_mem_MPORT_101_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_101_data = LUT_mem_MPORT_101_addr >= 6'h23 ? _RAND_102[32:0] : LUT_mem[LUT_mem_MPORT_101_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_102_addr = 6'h20;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_102_data = LUT_mem[LUT_mem_MPORT_102_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_102_data = LUT_mem_MPORT_102_addr >= 6'h23 ? _RAND_103[32:0] : LUT_mem[LUT_mem_MPORT_102_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_103_addr = 6'h21;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_103_data = LUT_mem[LUT_mem_MPORT_103_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_103_data = LUT_mem_MPORT_103_addr >= 6'h23 ? _RAND_104[32:0] : LUT_mem[LUT_mem_MPORT_103_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_104_addr = 6'h22;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_104_data = LUT_mem[LUT_mem_MPORT_104_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_104_data = LUT_mem_MPORT_104_addr >= 6'h23 ? _RAND_105[32:0] : LUT_mem[LUT_mem_MPORT_104_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_105_addr = 6'h0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_105_data = LUT_mem[LUT_mem_MPORT_105_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_105_data = LUT_mem_MPORT_105_addr >= 6'h23 ? _RAND_106[32:0] : LUT_mem[LUT_mem_MPORT_105_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_106_addr = 6'h1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_106_data = LUT_mem[LUT_mem_MPORT_106_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_106_data = LUT_mem_MPORT_106_addr >= 6'h23 ? _RAND_107[32:0] : LUT_mem[LUT_mem_MPORT_106_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_107_addr = 6'h2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_107_data = LUT_mem[LUT_mem_MPORT_107_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_107_data = LUT_mem_MPORT_107_addr >= 6'h23 ? _RAND_108[32:0] : LUT_mem[LUT_mem_MPORT_107_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_108_addr = 6'h3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_108_data = LUT_mem[LUT_mem_MPORT_108_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_108_data = LUT_mem_MPORT_108_addr >= 6'h23 ? _RAND_109[32:0] : LUT_mem[LUT_mem_MPORT_108_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_109_addr = 6'h4;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_109_data = LUT_mem[LUT_mem_MPORT_109_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_109_data = LUT_mem_MPORT_109_addr >= 6'h23 ? _RAND_110[32:0] : LUT_mem[LUT_mem_MPORT_109_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_110_addr = 6'h5;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_110_data = LUT_mem[LUT_mem_MPORT_110_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_110_data = LUT_mem_MPORT_110_addr >= 6'h23 ? _RAND_111[32:0] : LUT_mem[LUT_mem_MPORT_110_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_111_addr = 6'h6;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_111_data = LUT_mem[LUT_mem_MPORT_111_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_111_data = LUT_mem_MPORT_111_addr >= 6'h23 ? _RAND_112[32:0] : LUT_mem[LUT_mem_MPORT_111_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_112_addr = 6'h7;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_112_data = LUT_mem[LUT_mem_MPORT_112_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_112_data = LUT_mem_MPORT_112_addr >= 6'h23 ? _RAND_113[32:0] : LUT_mem[LUT_mem_MPORT_112_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_113_addr = 6'h8;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_113_data = LUT_mem[LUT_mem_MPORT_113_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_113_data = LUT_mem_MPORT_113_addr >= 6'h23 ? _RAND_114[32:0] : LUT_mem[LUT_mem_MPORT_113_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_114_addr = 6'h9;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_114_data = LUT_mem[LUT_mem_MPORT_114_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_114_data = LUT_mem_MPORT_114_addr >= 6'h23 ? _RAND_115[32:0] : LUT_mem[LUT_mem_MPORT_114_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_115_addr = 6'ha;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_115_data = LUT_mem[LUT_mem_MPORT_115_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_115_data = LUT_mem_MPORT_115_addr >= 6'h23 ? _RAND_116[32:0] : LUT_mem[LUT_mem_MPORT_115_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_116_addr = 6'hb;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_116_data = LUT_mem[LUT_mem_MPORT_116_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_116_data = LUT_mem_MPORT_116_addr >= 6'h23 ? _RAND_117[32:0] : LUT_mem[LUT_mem_MPORT_116_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_117_addr = 6'hc;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_117_data = LUT_mem[LUT_mem_MPORT_117_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_117_data = LUT_mem_MPORT_117_addr >= 6'h23 ? _RAND_118[32:0] : LUT_mem[LUT_mem_MPORT_117_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_118_addr = 6'hd;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_118_data = LUT_mem[LUT_mem_MPORT_118_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_118_data = LUT_mem_MPORT_118_addr >= 6'h23 ? _RAND_119[32:0] : LUT_mem[LUT_mem_MPORT_118_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_119_addr = 6'he;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_119_data = LUT_mem[LUT_mem_MPORT_119_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_119_data = LUT_mem_MPORT_119_addr >= 6'h23 ? _RAND_120[32:0] : LUT_mem[LUT_mem_MPORT_119_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_120_addr = 6'hf;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_120_data = LUT_mem[LUT_mem_MPORT_120_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_120_data = LUT_mem_MPORT_120_addr >= 6'h23 ? _RAND_121[32:0] : LUT_mem[LUT_mem_MPORT_120_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_121_addr = 6'h10;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_121_data = LUT_mem[LUT_mem_MPORT_121_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_121_data = LUT_mem_MPORT_121_addr >= 6'h23 ? _RAND_122[32:0] : LUT_mem[LUT_mem_MPORT_121_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_122_addr = 6'h11;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_122_data = LUT_mem[LUT_mem_MPORT_122_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_122_data = LUT_mem_MPORT_122_addr >= 6'h23 ? _RAND_123[32:0] : LUT_mem[LUT_mem_MPORT_122_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_123_addr = 6'h12;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_123_data = LUT_mem[LUT_mem_MPORT_123_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_123_data = LUT_mem_MPORT_123_addr >= 6'h23 ? _RAND_124[32:0] : LUT_mem[LUT_mem_MPORT_123_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_124_addr = 6'h13;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_124_data = LUT_mem[LUT_mem_MPORT_124_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_124_data = LUT_mem_MPORT_124_addr >= 6'h23 ? _RAND_125[32:0] : LUT_mem[LUT_mem_MPORT_124_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_125_addr = 6'h14;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_125_data = LUT_mem[LUT_mem_MPORT_125_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_125_data = LUT_mem_MPORT_125_addr >= 6'h23 ? _RAND_126[32:0] : LUT_mem[LUT_mem_MPORT_125_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_126_addr = 6'h15;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_126_data = LUT_mem[LUT_mem_MPORT_126_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_126_data = LUT_mem_MPORT_126_addr >= 6'h23 ? _RAND_127[32:0] : LUT_mem[LUT_mem_MPORT_126_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_127_addr = 6'h16;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_127_data = LUT_mem[LUT_mem_MPORT_127_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_127_data = LUT_mem_MPORT_127_addr >= 6'h23 ? _RAND_128[32:0] : LUT_mem[LUT_mem_MPORT_127_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_128_addr = 6'h17;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_128_data = LUT_mem[LUT_mem_MPORT_128_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_128_data = LUT_mem_MPORT_128_addr >= 6'h23 ? _RAND_129[32:0] : LUT_mem[LUT_mem_MPORT_128_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_129_addr = 6'h18;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_129_data = LUT_mem[LUT_mem_MPORT_129_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_129_data = LUT_mem_MPORT_129_addr >= 6'h23 ? _RAND_130[32:0] : LUT_mem[LUT_mem_MPORT_129_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_130_addr = 6'h19;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_130_data = LUT_mem[LUT_mem_MPORT_130_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_130_data = LUT_mem_MPORT_130_addr >= 6'h23 ? _RAND_131[32:0] : LUT_mem[LUT_mem_MPORT_130_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_131_addr = 6'h1a;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_131_data = LUT_mem[LUT_mem_MPORT_131_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_131_data = LUT_mem_MPORT_131_addr >= 6'h23 ? _RAND_132[32:0] : LUT_mem[LUT_mem_MPORT_131_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_132_addr = 6'h1b;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_132_data = LUT_mem[LUT_mem_MPORT_132_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_132_data = LUT_mem_MPORT_132_addr >= 6'h23 ? _RAND_133[32:0] : LUT_mem[LUT_mem_MPORT_132_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_133_addr = 6'h1c;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_133_data = LUT_mem[LUT_mem_MPORT_133_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_133_data = LUT_mem_MPORT_133_addr >= 6'h23 ? _RAND_134[32:0] : LUT_mem[LUT_mem_MPORT_133_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_134_addr = 6'h1d;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_134_data = LUT_mem[LUT_mem_MPORT_134_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_134_data = LUT_mem_MPORT_134_addr >= 6'h23 ? _RAND_135[32:0] : LUT_mem[LUT_mem_MPORT_134_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_135_addr = 6'h1e;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_135_data = LUT_mem[LUT_mem_MPORT_135_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_135_data = LUT_mem_MPORT_135_addr >= 6'h23 ? _RAND_136[32:0] : LUT_mem[LUT_mem_MPORT_135_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_136_addr = 6'h1f;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_136_data = LUT_mem[LUT_mem_MPORT_136_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_136_data = LUT_mem_MPORT_136_addr >= 6'h23 ? _RAND_137[32:0] : LUT_mem[LUT_mem_MPORT_136_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_137_addr = 6'h20;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_137_data = LUT_mem[LUT_mem_MPORT_137_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_137_data = LUT_mem_MPORT_137_addr >= 6'h23 ? _RAND_138[32:0] : LUT_mem[LUT_mem_MPORT_137_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_138_addr = 6'h21;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_138_data = LUT_mem[LUT_mem_MPORT_138_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_138_data = LUT_mem_MPORT_138_addr >= 6'h23 ? _RAND_139[32:0] : LUT_mem[LUT_mem_MPORT_138_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_139_addr = 6'h22;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_139_data = LUT_mem[LUT_mem_MPORT_139_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_139_data = LUT_mem_MPORT_139_addr >= 6'h23 ? _RAND_140[32:0] : LUT_mem[LUT_mem_MPORT_139_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_140_addr = 6'h0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_140_data = LUT_mem[LUT_mem_MPORT_140_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_140_data = LUT_mem_MPORT_140_addr >= 6'h23 ? _RAND_141[32:0] : LUT_mem[LUT_mem_MPORT_140_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_141_addr = 6'h1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_141_data = LUT_mem[LUT_mem_MPORT_141_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_141_data = LUT_mem_MPORT_141_addr >= 6'h23 ? _RAND_142[32:0] : LUT_mem[LUT_mem_MPORT_141_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_142_addr = 6'h2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_142_data = LUT_mem[LUT_mem_MPORT_142_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_142_data = LUT_mem_MPORT_142_addr >= 6'h23 ? _RAND_143[32:0] : LUT_mem[LUT_mem_MPORT_142_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_143_addr = 6'h3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_143_data = LUT_mem[LUT_mem_MPORT_143_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_143_data = LUT_mem_MPORT_143_addr >= 6'h23 ? _RAND_144[32:0] : LUT_mem[LUT_mem_MPORT_143_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_144_addr = 6'h4;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_144_data = LUT_mem[LUT_mem_MPORT_144_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_144_data = LUT_mem_MPORT_144_addr >= 6'h23 ? _RAND_145[32:0] : LUT_mem[LUT_mem_MPORT_144_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_145_addr = 6'h5;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_145_data = LUT_mem[LUT_mem_MPORT_145_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_145_data = LUT_mem_MPORT_145_addr >= 6'h23 ? _RAND_146[32:0] : LUT_mem[LUT_mem_MPORT_145_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_146_addr = 6'h6;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_146_data = LUT_mem[LUT_mem_MPORT_146_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_146_data = LUT_mem_MPORT_146_addr >= 6'h23 ? _RAND_147[32:0] : LUT_mem[LUT_mem_MPORT_146_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_147_addr = 6'h7;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_147_data = LUT_mem[LUT_mem_MPORT_147_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_147_data = LUT_mem_MPORT_147_addr >= 6'h23 ? _RAND_148[32:0] : LUT_mem[LUT_mem_MPORT_147_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_148_addr = 6'h8;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_148_data = LUT_mem[LUT_mem_MPORT_148_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_148_data = LUT_mem_MPORT_148_addr >= 6'h23 ? _RAND_149[32:0] : LUT_mem[LUT_mem_MPORT_148_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_149_addr = 6'h9;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_149_data = LUT_mem[LUT_mem_MPORT_149_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_149_data = LUT_mem_MPORT_149_addr >= 6'h23 ? _RAND_150[32:0] : LUT_mem[LUT_mem_MPORT_149_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_150_addr = 6'ha;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_150_data = LUT_mem[LUT_mem_MPORT_150_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_150_data = LUT_mem_MPORT_150_addr >= 6'h23 ? _RAND_151[32:0] : LUT_mem[LUT_mem_MPORT_150_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_151_addr = 6'hb;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_151_data = LUT_mem[LUT_mem_MPORT_151_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_151_data = LUT_mem_MPORT_151_addr >= 6'h23 ? _RAND_152[32:0] : LUT_mem[LUT_mem_MPORT_151_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_152_addr = 6'hc;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_152_data = LUT_mem[LUT_mem_MPORT_152_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_152_data = LUT_mem_MPORT_152_addr >= 6'h23 ? _RAND_153[32:0] : LUT_mem[LUT_mem_MPORT_152_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_153_addr = 6'hd;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_153_data = LUT_mem[LUT_mem_MPORT_153_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_153_data = LUT_mem_MPORT_153_addr >= 6'h23 ? _RAND_154[32:0] : LUT_mem[LUT_mem_MPORT_153_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_154_addr = 6'he;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_154_data = LUT_mem[LUT_mem_MPORT_154_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_154_data = LUT_mem_MPORT_154_addr >= 6'h23 ? _RAND_155[32:0] : LUT_mem[LUT_mem_MPORT_154_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_155_addr = 6'hf;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_155_data = LUT_mem[LUT_mem_MPORT_155_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_155_data = LUT_mem_MPORT_155_addr >= 6'h23 ? _RAND_156[32:0] : LUT_mem[LUT_mem_MPORT_155_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_156_addr = 6'h10;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_156_data = LUT_mem[LUT_mem_MPORT_156_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_156_data = LUT_mem_MPORT_156_addr >= 6'h23 ? _RAND_157[32:0] : LUT_mem[LUT_mem_MPORT_156_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_157_addr = 6'h11;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_157_data = LUT_mem[LUT_mem_MPORT_157_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_157_data = LUT_mem_MPORT_157_addr >= 6'h23 ? _RAND_158[32:0] : LUT_mem[LUT_mem_MPORT_157_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_158_addr = 6'h12;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_158_data = LUT_mem[LUT_mem_MPORT_158_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_158_data = LUT_mem_MPORT_158_addr >= 6'h23 ? _RAND_159[32:0] : LUT_mem[LUT_mem_MPORT_158_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_159_addr = 6'h13;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_159_data = LUT_mem[LUT_mem_MPORT_159_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_159_data = LUT_mem_MPORT_159_addr >= 6'h23 ? _RAND_160[32:0] : LUT_mem[LUT_mem_MPORT_159_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_160_addr = 6'h14;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_160_data = LUT_mem[LUT_mem_MPORT_160_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_160_data = LUT_mem_MPORT_160_addr >= 6'h23 ? _RAND_161[32:0] : LUT_mem[LUT_mem_MPORT_160_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_161_addr = 6'h15;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_161_data = LUT_mem[LUT_mem_MPORT_161_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_161_data = LUT_mem_MPORT_161_addr >= 6'h23 ? _RAND_162[32:0] : LUT_mem[LUT_mem_MPORT_161_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_162_addr = 6'h16;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_162_data = LUT_mem[LUT_mem_MPORT_162_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_162_data = LUT_mem_MPORT_162_addr >= 6'h23 ? _RAND_163[32:0] : LUT_mem[LUT_mem_MPORT_162_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_163_addr = 6'h17;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_163_data = LUT_mem[LUT_mem_MPORT_163_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_163_data = LUT_mem_MPORT_163_addr >= 6'h23 ? _RAND_164[32:0] : LUT_mem[LUT_mem_MPORT_163_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_164_addr = 6'h18;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_164_data = LUT_mem[LUT_mem_MPORT_164_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_164_data = LUT_mem_MPORT_164_addr >= 6'h23 ? _RAND_165[32:0] : LUT_mem[LUT_mem_MPORT_164_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_165_addr = 6'h19;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_165_data = LUT_mem[LUT_mem_MPORT_165_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_165_data = LUT_mem_MPORT_165_addr >= 6'h23 ? _RAND_166[32:0] : LUT_mem[LUT_mem_MPORT_165_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_166_addr = 6'h1a;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_166_data = LUT_mem[LUT_mem_MPORT_166_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_166_data = LUT_mem_MPORT_166_addr >= 6'h23 ? _RAND_167[32:0] : LUT_mem[LUT_mem_MPORT_166_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_167_addr = 6'h1b;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_167_data = LUT_mem[LUT_mem_MPORT_167_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_167_data = LUT_mem_MPORT_167_addr >= 6'h23 ? _RAND_168[32:0] : LUT_mem[LUT_mem_MPORT_167_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_168_addr = 6'h1c;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_168_data = LUT_mem[LUT_mem_MPORT_168_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_168_data = LUT_mem_MPORT_168_addr >= 6'h23 ? _RAND_169[32:0] : LUT_mem[LUT_mem_MPORT_168_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_169_addr = 6'h1d;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_169_data = LUT_mem[LUT_mem_MPORT_169_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_169_data = LUT_mem_MPORT_169_addr >= 6'h23 ? _RAND_170[32:0] : LUT_mem[LUT_mem_MPORT_169_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_170_addr = 6'h1e;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_170_data = LUT_mem[LUT_mem_MPORT_170_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_170_data = LUT_mem_MPORT_170_addr >= 6'h23 ? _RAND_171[32:0] : LUT_mem[LUT_mem_MPORT_170_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_171_addr = 6'h1f;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_171_data = LUT_mem[LUT_mem_MPORT_171_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_171_data = LUT_mem_MPORT_171_addr >= 6'h23 ? _RAND_172[32:0] : LUT_mem[LUT_mem_MPORT_171_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_172_addr = 6'h20;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_172_data = LUT_mem[LUT_mem_MPORT_172_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_172_data = LUT_mem_MPORT_172_addr >= 6'h23 ? _RAND_173[32:0] : LUT_mem[LUT_mem_MPORT_172_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_173_addr = 6'h21;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_173_data = LUT_mem[LUT_mem_MPORT_173_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_173_data = LUT_mem_MPORT_173_addr >= 6'h23 ? _RAND_174[32:0] : LUT_mem[LUT_mem_MPORT_173_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_174_addr = 6'h22;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_174_data = LUT_mem[LUT_mem_MPORT_174_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_174_data = LUT_mem_MPORT_174_addr >= 6'h23 ? _RAND_175[32:0] : LUT_mem[LUT_mem_MPORT_174_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_176_addr = 6'h0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_176_data = LUT_mem[LUT_mem_MPORT_176_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_176_data = LUT_mem_MPORT_176_addr >= 6'h23 ? _RAND_176[32:0] : LUT_mem[LUT_mem_MPORT_176_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_179_addr = 6'h0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_179_data = LUT_mem[LUT_mem_MPORT_179_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_179_data = LUT_mem_MPORT_179_addr >= 6'h23 ? _RAND_177[32:0] : LUT_mem[LUT_mem_MPORT_179_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_181_addr = 6'h1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_181_data = LUT_mem[LUT_mem_MPORT_181_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_181_data = LUT_mem_MPORT_181_addr >= 6'h23 ? _RAND_178[32:0] : LUT_mem[LUT_mem_MPORT_181_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_184_addr = 6'h1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_184_data = LUT_mem[LUT_mem_MPORT_184_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_184_data = LUT_mem_MPORT_184_addr >= 6'h23 ? _RAND_179[32:0] : LUT_mem[LUT_mem_MPORT_184_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_186_addr = 6'h2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_186_data = LUT_mem[LUT_mem_MPORT_186_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_186_data = LUT_mem_MPORT_186_addr >= 6'h23 ? _RAND_180[32:0] : LUT_mem[LUT_mem_MPORT_186_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_189_addr = 6'h2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_189_data = LUT_mem[LUT_mem_MPORT_189_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_189_data = LUT_mem_MPORT_189_addr >= 6'h23 ? _RAND_181[32:0] : LUT_mem[LUT_mem_MPORT_189_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_191_addr = 6'h3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_191_data = LUT_mem[LUT_mem_MPORT_191_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_191_data = LUT_mem_MPORT_191_addr >= 6'h23 ? _RAND_182[32:0] : LUT_mem[LUT_mem_MPORT_191_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_194_addr = 6'h3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_194_data = LUT_mem[LUT_mem_MPORT_194_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_194_data = LUT_mem_MPORT_194_addr >= 6'h23 ? _RAND_183[32:0] : LUT_mem[LUT_mem_MPORT_194_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_196_addr = 6'h4;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_196_data = LUT_mem[LUT_mem_MPORT_196_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_196_data = LUT_mem_MPORT_196_addr >= 6'h23 ? _RAND_184[32:0] : LUT_mem[LUT_mem_MPORT_196_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_199_addr = 6'h4;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_199_data = LUT_mem[LUT_mem_MPORT_199_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_199_data = LUT_mem_MPORT_199_addr >= 6'h23 ? _RAND_185[32:0] : LUT_mem[LUT_mem_MPORT_199_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_201_addr = 6'h5;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_201_data = LUT_mem[LUT_mem_MPORT_201_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_201_data = LUT_mem_MPORT_201_addr >= 6'h23 ? _RAND_186[32:0] : LUT_mem[LUT_mem_MPORT_201_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_204_addr = 6'h5;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_204_data = LUT_mem[LUT_mem_MPORT_204_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_204_data = LUT_mem_MPORT_204_addr >= 6'h23 ? _RAND_187[32:0] : LUT_mem[LUT_mem_MPORT_204_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_206_addr = 6'h6;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_206_data = LUT_mem[LUT_mem_MPORT_206_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_206_data = LUT_mem_MPORT_206_addr >= 6'h23 ? _RAND_188[32:0] : LUT_mem[LUT_mem_MPORT_206_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_209_addr = 6'h6;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_209_data = LUT_mem[LUT_mem_MPORT_209_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_209_data = LUT_mem_MPORT_209_addr >= 6'h23 ? _RAND_189[32:0] : LUT_mem[LUT_mem_MPORT_209_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_211_addr = 6'h7;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_211_data = LUT_mem[LUT_mem_MPORT_211_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_211_data = LUT_mem_MPORT_211_addr >= 6'h23 ? _RAND_190[32:0] : LUT_mem[LUT_mem_MPORT_211_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_214_addr = 6'h7;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_214_data = LUT_mem[LUT_mem_MPORT_214_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_214_data = LUT_mem_MPORT_214_addr >= 6'h23 ? _RAND_191[32:0] : LUT_mem[LUT_mem_MPORT_214_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_216_addr = 6'h8;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_216_data = LUT_mem[LUT_mem_MPORT_216_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_216_data = LUT_mem_MPORT_216_addr >= 6'h23 ? _RAND_192[32:0] : LUT_mem[LUT_mem_MPORT_216_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_219_addr = 6'h8;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_219_data = LUT_mem[LUT_mem_MPORT_219_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_219_data = LUT_mem_MPORT_219_addr >= 6'h23 ? _RAND_193[32:0] : LUT_mem[LUT_mem_MPORT_219_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_221_addr = 6'h9;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_221_data = LUT_mem[LUT_mem_MPORT_221_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_221_data = LUT_mem_MPORT_221_addr >= 6'h23 ? _RAND_194[32:0] : LUT_mem[LUT_mem_MPORT_221_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_224_addr = 6'h9;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_224_data = LUT_mem[LUT_mem_MPORT_224_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_224_data = LUT_mem_MPORT_224_addr >= 6'h23 ? _RAND_195[32:0] : LUT_mem[LUT_mem_MPORT_224_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_226_addr = 6'ha;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_226_data = LUT_mem[LUT_mem_MPORT_226_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_226_data = LUT_mem_MPORT_226_addr >= 6'h23 ? _RAND_196[32:0] : LUT_mem[LUT_mem_MPORT_226_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_229_addr = 6'ha;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_229_data = LUT_mem[LUT_mem_MPORT_229_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_229_data = LUT_mem_MPORT_229_addr >= 6'h23 ? _RAND_197[32:0] : LUT_mem[LUT_mem_MPORT_229_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_231_addr = 6'hb;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_231_data = LUT_mem[LUT_mem_MPORT_231_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_231_data = LUT_mem_MPORT_231_addr >= 6'h23 ? _RAND_198[32:0] : LUT_mem[LUT_mem_MPORT_231_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_234_addr = 6'hb;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_234_data = LUT_mem[LUT_mem_MPORT_234_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_234_data = LUT_mem_MPORT_234_addr >= 6'h23 ? _RAND_199[32:0] : LUT_mem[LUT_mem_MPORT_234_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_236_addr = 6'hc;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_236_data = LUT_mem[LUT_mem_MPORT_236_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_236_data = LUT_mem_MPORT_236_addr >= 6'h23 ? _RAND_200[32:0] : LUT_mem[LUT_mem_MPORT_236_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_239_addr = 6'hc;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_239_data = LUT_mem[LUT_mem_MPORT_239_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_239_data = LUT_mem_MPORT_239_addr >= 6'h23 ? _RAND_201[32:0] : LUT_mem[LUT_mem_MPORT_239_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_241_addr = 6'hd;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_241_data = LUT_mem[LUT_mem_MPORT_241_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_241_data = LUT_mem_MPORT_241_addr >= 6'h23 ? _RAND_202[32:0] : LUT_mem[LUT_mem_MPORT_241_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_244_addr = 6'hd;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_244_data = LUT_mem[LUT_mem_MPORT_244_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_244_data = LUT_mem_MPORT_244_addr >= 6'h23 ? _RAND_203[32:0] : LUT_mem[LUT_mem_MPORT_244_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_246_addr = 6'he;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_246_data = LUT_mem[LUT_mem_MPORT_246_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_246_data = LUT_mem_MPORT_246_addr >= 6'h23 ? _RAND_204[32:0] : LUT_mem[LUT_mem_MPORT_246_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_249_addr = 6'he;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_249_data = LUT_mem[LUT_mem_MPORT_249_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_249_data = LUT_mem_MPORT_249_addr >= 6'h23 ? _RAND_205[32:0] : LUT_mem[LUT_mem_MPORT_249_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_251_addr = 6'hf;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_251_data = LUT_mem[LUT_mem_MPORT_251_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_251_data = LUT_mem_MPORT_251_addr >= 6'h23 ? _RAND_206[32:0] : LUT_mem[LUT_mem_MPORT_251_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_254_addr = 6'hf;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_254_data = LUT_mem[LUT_mem_MPORT_254_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_254_data = LUT_mem_MPORT_254_addr >= 6'h23 ? _RAND_207[32:0] : LUT_mem[LUT_mem_MPORT_254_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_256_addr = 6'h10;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_256_data = LUT_mem[LUT_mem_MPORT_256_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_256_data = LUT_mem_MPORT_256_addr >= 6'h23 ? _RAND_208[32:0] : LUT_mem[LUT_mem_MPORT_256_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_259_addr = 6'h10;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_259_data = LUT_mem[LUT_mem_MPORT_259_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_259_data = LUT_mem_MPORT_259_addr >= 6'h23 ? _RAND_209[32:0] : LUT_mem[LUT_mem_MPORT_259_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_261_addr = 6'h11;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_261_data = LUT_mem[LUT_mem_MPORT_261_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_261_data = LUT_mem_MPORT_261_addr >= 6'h23 ? _RAND_210[32:0] : LUT_mem[LUT_mem_MPORT_261_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_264_addr = 6'h11;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_264_data = LUT_mem[LUT_mem_MPORT_264_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_264_data = LUT_mem_MPORT_264_addr >= 6'h23 ? _RAND_211[32:0] : LUT_mem[LUT_mem_MPORT_264_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_266_addr = 6'h12;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_266_data = LUT_mem[LUT_mem_MPORT_266_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_266_data = LUT_mem_MPORT_266_addr >= 6'h23 ? _RAND_212[32:0] : LUT_mem[LUT_mem_MPORT_266_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_269_addr = 6'h12;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_269_data = LUT_mem[LUT_mem_MPORT_269_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_269_data = LUT_mem_MPORT_269_addr >= 6'h23 ? _RAND_213[32:0] : LUT_mem[LUT_mem_MPORT_269_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_271_addr = 6'h13;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_271_data = LUT_mem[LUT_mem_MPORT_271_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_271_data = LUT_mem_MPORT_271_addr >= 6'h23 ? _RAND_214[32:0] : LUT_mem[LUT_mem_MPORT_271_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_274_addr = 6'h13;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_274_data = LUT_mem[LUT_mem_MPORT_274_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_274_data = LUT_mem_MPORT_274_addr >= 6'h23 ? _RAND_215[32:0] : LUT_mem[LUT_mem_MPORT_274_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_276_addr = 6'h14;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_276_data = LUT_mem[LUT_mem_MPORT_276_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_276_data = LUT_mem_MPORT_276_addr >= 6'h23 ? _RAND_216[32:0] : LUT_mem[LUT_mem_MPORT_276_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_279_addr = 6'h14;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_279_data = LUT_mem[LUT_mem_MPORT_279_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_279_data = LUT_mem_MPORT_279_addr >= 6'h23 ? _RAND_217[32:0] : LUT_mem[LUT_mem_MPORT_279_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_281_addr = 6'h15;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_281_data = LUT_mem[LUT_mem_MPORT_281_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_281_data = LUT_mem_MPORT_281_addr >= 6'h23 ? _RAND_218[32:0] : LUT_mem[LUT_mem_MPORT_281_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_284_addr = 6'h15;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_284_data = LUT_mem[LUT_mem_MPORT_284_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_284_data = LUT_mem_MPORT_284_addr >= 6'h23 ? _RAND_219[32:0] : LUT_mem[LUT_mem_MPORT_284_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_286_addr = 6'h16;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_286_data = LUT_mem[LUT_mem_MPORT_286_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_286_data = LUT_mem_MPORT_286_addr >= 6'h23 ? _RAND_220[32:0] : LUT_mem[LUT_mem_MPORT_286_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_289_addr = 6'h16;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_289_data = LUT_mem[LUT_mem_MPORT_289_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_289_data = LUT_mem_MPORT_289_addr >= 6'h23 ? _RAND_221[32:0] : LUT_mem[LUT_mem_MPORT_289_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_291_addr = 6'h17;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_291_data = LUT_mem[LUT_mem_MPORT_291_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_291_data = LUT_mem_MPORT_291_addr >= 6'h23 ? _RAND_222[32:0] : LUT_mem[LUT_mem_MPORT_291_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_294_addr = 6'h17;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_294_data = LUT_mem[LUT_mem_MPORT_294_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_294_data = LUT_mem_MPORT_294_addr >= 6'h23 ? _RAND_223[32:0] : LUT_mem[LUT_mem_MPORT_294_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_296_addr = 6'h18;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_296_data = LUT_mem[LUT_mem_MPORT_296_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_296_data = LUT_mem_MPORT_296_addr >= 6'h23 ? _RAND_224[32:0] : LUT_mem[LUT_mem_MPORT_296_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_299_addr = 6'h18;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_299_data = LUT_mem[LUT_mem_MPORT_299_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_299_data = LUT_mem_MPORT_299_addr >= 6'h23 ? _RAND_225[32:0] : LUT_mem[LUT_mem_MPORT_299_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_301_addr = 6'h19;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_301_data = LUT_mem[LUT_mem_MPORT_301_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_301_data = LUT_mem_MPORT_301_addr >= 6'h23 ? _RAND_226[32:0] : LUT_mem[LUT_mem_MPORT_301_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_304_addr = 6'h19;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_304_data = LUT_mem[LUT_mem_MPORT_304_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_304_data = LUT_mem_MPORT_304_addr >= 6'h23 ? _RAND_227[32:0] : LUT_mem[LUT_mem_MPORT_304_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_306_addr = 6'h1a;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_306_data = LUT_mem[LUT_mem_MPORT_306_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_306_data = LUT_mem_MPORT_306_addr >= 6'h23 ? _RAND_228[32:0] : LUT_mem[LUT_mem_MPORT_306_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_309_addr = 6'h1a;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_309_data = LUT_mem[LUT_mem_MPORT_309_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_309_data = LUT_mem_MPORT_309_addr >= 6'h23 ? _RAND_229[32:0] : LUT_mem[LUT_mem_MPORT_309_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_311_addr = 6'h1b;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_311_data = LUT_mem[LUT_mem_MPORT_311_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_311_data = LUT_mem_MPORT_311_addr >= 6'h23 ? _RAND_230[32:0] : LUT_mem[LUT_mem_MPORT_311_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_314_addr = 6'h1b;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_314_data = LUT_mem[LUT_mem_MPORT_314_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_314_data = LUT_mem_MPORT_314_addr >= 6'h23 ? _RAND_231[32:0] : LUT_mem[LUT_mem_MPORT_314_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_316_addr = 6'h1c;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_316_data = LUT_mem[LUT_mem_MPORT_316_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_316_data = LUT_mem_MPORT_316_addr >= 6'h23 ? _RAND_232[32:0] : LUT_mem[LUT_mem_MPORT_316_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_319_addr = 6'h1c;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_319_data = LUT_mem[LUT_mem_MPORT_319_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_319_data = LUT_mem_MPORT_319_addr >= 6'h23 ? _RAND_233[32:0] : LUT_mem[LUT_mem_MPORT_319_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_321_addr = 6'h1d;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_321_data = LUT_mem[LUT_mem_MPORT_321_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_321_data = LUT_mem_MPORT_321_addr >= 6'h23 ? _RAND_234[32:0] : LUT_mem[LUT_mem_MPORT_321_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_324_addr = 6'h1d;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_324_data = LUT_mem[LUT_mem_MPORT_324_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_324_data = LUT_mem_MPORT_324_addr >= 6'h23 ? _RAND_235[32:0] : LUT_mem[LUT_mem_MPORT_324_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_326_addr = 6'h1e;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_326_data = LUT_mem[LUT_mem_MPORT_326_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_326_data = LUT_mem_MPORT_326_addr >= 6'h23 ? _RAND_236[32:0] : LUT_mem[LUT_mem_MPORT_326_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_329_addr = 6'h1e;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_329_data = LUT_mem[LUT_mem_MPORT_329_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_329_data = LUT_mem_MPORT_329_addr >= 6'h23 ? _RAND_237[32:0] : LUT_mem[LUT_mem_MPORT_329_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_331_addr = 6'h1f;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_331_data = LUT_mem[LUT_mem_MPORT_331_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_331_data = LUT_mem_MPORT_331_addr >= 6'h23 ? _RAND_238[32:0] : LUT_mem[LUT_mem_MPORT_331_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_334_addr = 6'h1f;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_334_data = LUT_mem[LUT_mem_MPORT_334_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_334_data = LUT_mem_MPORT_334_addr >= 6'h23 ? _RAND_239[32:0] : LUT_mem[LUT_mem_MPORT_334_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_336_addr = 6'h20;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_336_data = LUT_mem[LUT_mem_MPORT_336_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_336_data = LUT_mem_MPORT_336_addr >= 6'h23 ? _RAND_240[32:0] : LUT_mem[LUT_mem_MPORT_336_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_339_addr = 6'h20;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_339_data = LUT_mem[LUT_mem_MPORT_339_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_339_data = LUT_mem_MPORT_339_addr >= 6'h23 ? _RAND_241[32:0] : LUT_mem[LUT_mem_MPORT_339_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_341_addr = 6'h21;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_341_data = LUT_mem[LUT_mem_MPORT_341_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_341_data = LUT_mem_MPORT_341_addr >= 6'h23 ? _RAND_242[32:0] : LUT_mem[LUT_mem_MPORT_341_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_344_addr = 6'h21;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_344_data = LUT_mem[LUT_mem_MPORT_344_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_344_data = LUT_mem_MPORT_344_addr >= 6'h23 ? _RAND_243[32:0] : LUT_mem[LUT_mem_MPORT_344_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_346_addr = 6'h22;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_346_data = LUT_mem[LUT_mem_MPORT_346_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_346_data = LUT_mem_MPORT_346_addr >= 6'h23 ? _RAND_244[32:0] : LUT_mem[LUT_mem_MPORT_346_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_349_addr = 6'h22;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_349_data = LUT_mem[LUT_mem_MPORT_349_addr]; // @[lut_35.scala 216:26]
  `else
  assign LUT_mem_MPORT_349_data = LUT_mem_MPORT_349_addr >= 6'h23 ? _RAND_245[32:0] : LUT_mem[LUT_mem_MPORT_349_addr]; // @[lut_35.scala 216:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_175_data = {1'h0,lo};
  assign LUT_mem_MPORT_175_addr = 6'h0;
  assign LUT_mem_MPORT_175_mask = 1'h1;
  assign LUT_mem_MPORT_175_en = dispatch_reg_0 | clear_0_1;
  assign LUT_mem_MPORT_177_data = {1'h1,push_id_temp};
  assign LUT_mem_MPORT_177_addr = 6'h0;
  assign LUT_mem_MPORT_177_mask = 1'h1;
  assign LUT_mem_MPORT_177_en = _T_895 ? 1'h0 : _T_897;
  assign LUT_mem_MPORT_178_data = LUT_mem_MPORT_179_data;
  assign LUT_mem_MPORT_178_addr = 6'h0;
  assign LUT_mem_MPORT_178_mask = 1'h1;
  assign LUT_mem_MPORT_178_en = _T_895 ? 1'h0 : _GEN_11436;
  assign LUT_mem_MPORT_180_data = {1'h0,lo_1};
  assign LUT_mem_MPORT_180_addr = 6'h1;
  assign LUT_mem_MPORT_180_mask = 1'h1;
  assign LUT_mem_MPORT_180_en = dispatch_reg_1 | clear_1_1;
  assign LUT_mem_MPORT_182_data = {1'h1,push_id_temp};
  assign LUT_mem_MPORT_182_addr = 6'h1;
  assign LUT_mem_MPORT_182_mask = 1'h1;
  assign LUT_mem_MPORT_182_en = _T_901 ? 1'h0 : _T_903;
  assign LUT_mem_MPORT_183_data = LUT_mem_MPORT_184_data;
  assign LUT_mem_MPORT_183_addr = 6'h1;
  assign LUT_mem_MPORT_183_mask = 1'h1;
  assign LUT_mem_MPORT_183_en = _T_901 ? 1'h0 : _GEN_11460;
  assign LUT_mem_MPORT_185_data = {1'h0,lo_2};
  assign LUT_mem_MPORT_185_addr = 6'h2;
  assign LUT_mem_MPORT_185_mask = 1'h1;
  assign LUT_mem_MPORT_185_en = dispatch_reg_2 | clear_2_1;
  assign LUT_mem_MPORT_187_data = {1'h1,push_id_temp};
  assign LUT_mem_MPORT_187_addr = 6'h2;
  assign LUT_mem_MPORT_187_mask = 1'h1;
  assign LUT_mem_MPORT_187_en = _T_907 ? 1'h0 : _T_909;
  assign LUT_mem_MPORT_188_data = LUT_mem_MPORT_189_data;
  assign LUT_mem_MPORT_188_addr = 6'h2;
  assign LUT_mem_MPORT_188_mask = 1'h1;
  assign LUT_mem_MPORT_188_en = _T_907 ? 1'h0 : _GEN_11481;
  assign LUT_mem_MPORT_190_data = {1'h0,lo_3};
  assign LUT_mem_MPORT_190_addr = 6'h3;
  assign LUT_mem_MPORT_190_mask = 1'h1;
  assign LUT_mem_MPORT_190_en = dispatch_reg_3 | clear_3_1;
  assign LUT_mem_MPORT_192_data = {1'h1,push_id_temp};
  assign LUT_mem_MPORT_192_addr = 6'h3;
  assign LUT_mem_MPORT_192_mask = 1'h1;
  assign LUT_mem_MPORT_192_en = _T_913 ? 1'h0 : _T_915;
  assign LUT_mem_MPORT_193_data = LUT_mem_MPORT_194_data;
  assign LUT_mem_MPORT_193_addr = 6'h3;
  assign LUT_mem_MPORT_193_mask = 1'h1;
  assign LUT_mem_MPORT_193_en = _T_913 ? 1'h0 : _GEN_11506;
  assign LUT_mem_MPORT_195_data = {1'h0,lo_4};
  assign LUT_mem_MPORT_195_addr = 6'h4;
  assign LUT_mem_MPORT_195_mask = 1'h1;
  assign LUT_mem_MPORT_195_en = dispatch_reg_4 | clear_4_1;
  assign LUT_mem_MPORT_197_data = {1'h1,push_id_temp};
  assign LUT_mem_MPORT_197_addr = 6'h4;
  assign LUT_mem_MPORT_197_mask = 1'h1;
  assign LUT_mem_MPORT_197_en = _T_919 ? 1'h0 : _T_921;
  assign LUT_mem_MPORT_198_data = LUT_mem_MPORT_199_data;
  assign LUT_mem_MPORT_198_addr = 6'h4;
  assign LUT_mem_MPORT_198_mask = 1'h1;
  assign LUT_mem_MPORT_198_en = _T_919 ? 1'h0 : _GEN_11531;
  assign LUT_mem_MPORT_200_data = {1'h0,lo_5};
  assign LUT_mem_MPORT_200_addr = 6'h5;
  assign LUT_mem_MPORT_200_mask = 1'h1;
  assign LUT_mem_MPORT_200_en = dispatch_reg_5 | clear_5_1;
  assign LUT_mem_MPORT_202_data = {1'h1,push_id_temp};
  assign LUT_mem_MPORT_202_addr = 6'h5;
  assign LUT_mem_MPORT_202_mask = 1'h1;
  assign LUT_mem_MPORT_202_en = _T_925 ? 1'h0 : _T_927;
  assign LUT_mem_MPORT_203_data = LUT_mem_MPORT_204_data;
  assign LUT_mem_MPORT_203_addr = 6'h5;
  assign LUT_mem_MPORT_203_mask = 1'h1;
  assign LUT_mem_MPORT_203_en = _T_925 ? 1'h0 : _GEN_11556;
  assign LUT_mem_MPORT_205_data = {1'h0,lo_6};
  assign LUT_mem_MPORT_205_addr = 6'h6;
  assign LUT_mem_MPORT_205_mask = 1'h1;
  assign LUT_mem_MPORT_205_en = dispatch_reg_6 | clear_6_1;
  assign LUT_mem_MPORT_207_data = {1'h1,push_id_temp};
  assign LUT_mem_MPORT_207_addr = 6'h6;
  assign LUT_mem_MPORT_207_mask = 1'h1;
  assign LUT_mem_MPORT_207_en = _T_931 ? 1'h0 : _T_933;
  assign LUT_mem_MPORT_208_data = LUT_mem_MPORT_209_data;
  assign LUT_mem_MPORT_208_addr = 6'h6;
  assign LUT_mem_MPORT_208_mask = 1'h1;
  assign LUT_mem_MPORT_208_en = _T_931 ? 1'h0 : _GEN_11581;
  assign LUT_mem_MPORT_210_data = {1'h0,lo_7};
  assign LUT_mem_MPORT_210_addr = 6'h7;
  assign LUT_mem_MPORT_210_mask = 1'h1;
  assign LUT_mem_MPORT_210_en = dispatch_reg_7 | clear_7_1;
  assign LUT_mem_MPORT_212_data = {1'h1,push_id_temp};
  assign LUT_mem_MPORT_212_addr = 6'h7;
  assign LUT_mem_MPORT_212_mask = 1'h1;
  assign LUT_mem_MPORT_212_en = _T_937 ? 1'h0 : _T_939;
  assign LUT_mem_MPORT_213_data = LUT_mem_MPORT_214_data;
  assign LUT_mem_MPORT_213_addr = 6'h7;
  assign LUT_mem_MPORT_213_mask = 1'h1;
  assign LUT_mem_MPORT_213_en = _T_937 ? 1'h0 : _GEN_11606;
  assign LUT_mem_MPORT_215_data = {1'h0,lo_8};
  assign LUT_mem_MPORT_215_addr = 6'h8;
  assign LUT_mem_MPORT_215_mask = 1'h1;
  assign LUT_mem_MPORT_215_en = dispatch_reg_8 | clear_8_1;
  assign LUT_mem_MPORT_217_data = {1'h1,push_id_temp};
  assign LUT_mem_MPORT_217_addr = 6'h8;
  assign LUT_mem_MPORT_217_mask = 1'h1;
  assign LUT_mem_MPORT_217_en = _T_943 ? 1'h0 : _T_945;
  assign LUT_mem_MPORT_218_data = LUT_mem_MPORT_219_data;
  assign LUT_mem_MPORT_218_addr = 6'h8;
  assign LUT_mem_MPORT_218_mask = 1'h1;
  assign LUT_mem_MPORT_218_en = _T_943 ? 1'h0 : _GEN_11631;
  assign LUT_mem_MPORT_220_data = {1'h0,lo_9};
  assign LUT_mem_MPORT_220_addr = 6'h9;
  assign LUT_mem_MPORT_220_mask = 1'h1;
  assign LUT_mem_MPORT_220_en = dispatch_reg_9 | clear_9_1;
  assign LUT_mem_MPORT_222_data = {1'h1,push_id_temp};
  assign LUT_mem_MPORT_222_addr = 6'h9;
  assign LUT_mem_MPORT_222_mask = 1'h1;
  assign LUT_mem_MPORT_222_en = _T_949 ? 1'h0 : _T_951;
  assign LUT_mem_MPORT_223_data = LUT_mem_MPORT_224_data;
  assign LUT_mem_MPORT_223_addr = 6'h9;
  assign LUT_mem_MPORT_223_mask = 1'h1;
  assign LUT_mem_MPORT_223_en = _T_949 ? 1'h0 : _GEN_11656;
  assign LUT_mem_MPORT_225_data = {1'h0,lo_10};
  assign LUT_mem_MPORT_225_addr = 6'ha;
  assign LUT_mem_MPORT_225_mask = 1'h1;
  assign LUT_mem_MPORT_225_en = dispatch_reg_10 | clear_10_1;
  assign LUT_mem_MPORT_227_data = {1'h1,push_id_temp};
  assign LUT_mem_MPORT_227_addr = 6'ha;
  assign LUT_mem_MPORT_227_mask = 1'h1;
  assign LUT_mem_MPORT_227_en = _T_955 ? 1'h0 : _T_957;
  assign LUT_mem_MPORT_228_data = LUT_mem_MPORT_229_data;
  assign LUT_mem_MPORT_228_addr = 6'ha;
  assign LUT_mem_MPORT_228_mask = 1'h1;
  assign LUT_mem_MPORT_228_en = _T_955 ? 1'h0 : _GEN_11681;
  assign LUT_mem_MPORT_230_data = {1'h0,lo_11};
  assign LUT_mem_MPORT_230_addr = 6'hb;
  assign LUT_mem_MPORT_230_mask = 1'h1;
  assign LUT_mem_MPORT_230_en = dispatch_reg_11 | clear_11_1;
  assign LUT_mem_MPORT_232_data = {1'h1,push_id_temp};
  assign LUT_mem_MPORT_232_addr = 6'hb;
  assign LUT_mem_MPORT_232_mask = 1'h1;
  assign LUT_mem_MPORT_232_en = _T_961 ? 1'h0 : _T_963;
  assign LUT_mem_MPORT_233_data = LUT_mem_MPORT_234_data;
  assign LUT_mem_MPORT_233_addr = 6'hb;
  assign LUT_mem_MPORT_233_mask = 1'h1;
  assign LUT_mem_MPORT_233_en = _T_961 ? 1'h0 : _GEN_11706;
  assign LUT_mem_MPORT_235_data = {1'h0,lo_12};
  assign LUT_mem_MPORT_235_addr = 6'hc;
  assign LUT_mem_MPORT_235_mask = 1'h1;
  assign LUT_mem_MPORT_235_en = dispatch_reg_12 | clear_12_1;
  assign LUT_mem_MPORT_237_data = {1'h1,push_id_temp};
  assign LUT_mem_MPORT_237_addr = 6'hc;
  assign LUT_mem_MPORT_237_mask = 1'h1;
  assign LUT_mem_MPORT_237_en = _T_967 ? 1'h0 : _T_969;
  assign LUT_mem_MPORT_238_data = LUT_mem_MPORT_239_data;
  assign LUT_mem_MPORT_238_addr = 6'hc;
  assign LUT_mem_MPORT_238_mask = 1'h1;
  assign LUT_mem_MPORT_238_en = _T_967 ? 1'h0 : _GEN_11731;
  assign LUT_mem_MPORT_240_data = {1'h0,lo_13};
  assign LUT_mem_MPORT_240_addr = 6'hd;
  assign LUT_mem_MPORT_240_mask = 1'h1;
  assign LUT_mem_MPORT_240_en = dispatch_reg_13 | clear_13_1;
  assign LUT_mem_MPORT_242_data = {1'h1,push_id_temp};
  assign LUT_mem_MPORT_242_addr = 6'hd;
  assign LUT_mem_MPORT_242_mask = 1'h1;
  assign LUT_mem_MPORT_242_en = _T_973 ? 1'h0 : _T_975;
  assign LUT_mem_MPORT_243_data = LUT_mem_MPORT_244_data;
  assign LUT_mem_MPORT_243_addr = 6'hd;
  assign LUT_mem_MPORT_243_mask = 1'h1;
  assign LUT_mem_MPORT_243_en = _T_973 ? 1'h0 : _GEN_11756;
  assign LUT_mem_MPORT_245_data = {1'h0,lo_14};
  assign LUT_mem_MPORT_245_addr = 6'he;
  assign LUT_mem_MPORT_245_mask = 1'h1;
  assign LUT_mem_MPORT_245_en = dispatch_reg_14 | clear_14_1;
  assign LUT_mem_MPORT_247_data = {1'h1,push_id_temp};
  assign LUT_mem_MPORT_247_addr = 6'he;
  assign LUT_mem_MPORT_247_mask = 1'h1;
  assign LUT_mem_MPORT_247_en = _T_979 ? 1'h0 : _T_981;
  assign LUT_mem_MPORT_248_data = LUT_mem_MPORT_249_data;
  assign LUT_mem_MPORT_248_addr = 6'he;
  assign LUT_mem_MPORT_248_mask = 1'h1;
  assign LUT_mem_MPORT_248_en = _T_979 ? 1'h0 : _GEN_11781;
  assign LUT_mem_MPORT_250_data = {1'h0,lo_15};
  assign LUT_mem_MPORT_250_addr = 6'hf;
  assign LUT_mem_MPORT_250_mask = 1'h1;
  assign LUT_mem_MPORT_250_en = dispatch_reg_15 | clear_15_1;
  assign LUT_mem_MPORT_252_data = {1'h1,push_id_temp};
  assign LUT_mem_MPORT_252_addr = 6'hf;
  assign LUT_mem_MPORT_252_mask = 1'h1;
  assign LUT_mem_MPORT_252_en = _T_985 ? 1'h0 : _T_987;
  assign LUT_mem_MPORT_253_data = LUT_mem_MPORT_254_data;
  assign LUT_mem_MPORT_253_addr = 6'hf;
  assign LUT_mem_MPORT_253_mask = 1'h1;
  assign LUT_mem_MPORT_253_en = _T_985 ? 1'h0 : _GEN_11806;
  assign LUT_mem_MPORT_255_data = {1'h0,lo_16};
  assign LUT_mem_MPORT_255_addr = 6'h10;
  assign LUT_mem_MPORT_255_mask = 1'h1;
  assign LUT_mem_MPORT_255_en = dispatch_reg_16 | clear_16_1;
  assign LUT_mem_MPORT_257_data = {1'h1,push_id_temp};
  assign LUT_mem_MPORT_257_addr = 6'h10;
  assign LUT_mem_MPORT_257_mask = 1'h1;
  assign LUT_mem_MPORT_257_en = _T_991 ? 1'h0 : _T_993;
  assign LUT_mem_MPORT_258_data = LUT_mem_MPORT_259_data;
  assign LUT_mem_MPORT_258_addr = 6'h10;
  assign LUT_mem_MPORT_258_mask = 1'h1;
  assign LUT_mem_MPORT_258_en = _T_991 ? 1'h0 : _GEN_11831;
  assign LUT_mem_MPORT_260_data = {1'h0,lo_17};
  assign LUT_mem_MPORT_260_addr = 6'h11;
  assign LUT_mem_MPORT_260_mask = 1'h1;
  assign LUT_mem_MPORT_260_en = dispatch_reg_17 | clear_17_1;
  assign LUT_mem_MPORT_262_data = {1'h1,push_id_temp};
  assign LUT_mem_MPORT_262_addr = 6'h11;
  assign LUT_mem_MPORT_262_mask = 1'h1;
  assign LUT_mem_MPORT_262_en = _T_997 ? 1'h0 : _T_999;
  assign LUT_mem_MPORT_263_data = LUT_mem_MPORT_264_data;
  assign LUT_mem_MPORT_263_addr = 6'h11;
  assign LUT_mem_MPORT_263_mask = 1'h1;
  assign LUT_mem_MPORT_263_en = _T_997 ? 1'h0 : _GEN_11856;
  assign LUT_mem_MPORT_265_data = {1'h0,lo_18};
  assign LUT_mem_MPORT_265_addr = 6'h12;
  assign LUT_mem_MPORT_265_mask = 1'h1;
  assign LUT_mem_MPORT_265_en = dispatch_reg_18 | clear_18_1;
  assign LUT_mem_MPORT_267_data = {1'h1,push_id_temp};
  assign LUT_mem_MPORT_267_addr = 6'h12;
  assign LUT_mem_MPORT_267_mask = 1'h1;
  assign LUT_mem_MPORT_267_en = _T_1003 ? 1'h0 : _T_1005;
  assign LUT_mem_MPORT_268_data = LUT_mem_MPORT_269_data;
  assign LUT_mem_MPORT_268_addr = 6'h12;
  assign LUT_mem_MPORT_268_mask = 1'h1;
  assign LUT_mem_MPORT_268_en = _T_1003 ? 1'h0 : _GEN_11881;
  assign LUT_mem_MPORT_270_data = {1'h0,lo_19};
  assign LUT_mem_MPORT_270_addr = 6'h13;
  assign LUT_mem_MPORT_270_mask = 1'h1;
  assign LUT_mem_MPORT_270_en = dispatch_reg_19 | clear_19_1;
  assign LUT_mem_MPORT_272_data = {1'h1,push_id_temp};
  assign LUT_mem_MPORT_272_addr = 6'h13;
  assign LUT_mem_MPORT_272_mask = 1'h1;
  assign LUT_mem_MPORT_272_en = _T_1009 ? 1'h0 : _T_1011;
  assign LUT_mem_MPORT_273_data = LUT_mem_MPORT_274_data;
  assign LUT_mem_MPORT_273_addr = 6'h13;
  assign LUT_mem_MPORT_273_mask = 1'h1;
  assign LUT_mem_MPORT_273_en = _T_1009 ? 1'h0 : _GEN_11906;
  assign LUT_mem_MPORT_275_data = {1'h0,lo_20};
  assign LUT_mem_MPORT_275_addr = 6'h14;
  assign LUT_mem_MPORT_275_mask = 1'h1;
  assign LUT_mem_MPORT_275_en = dispatch_reg_20 | clear_20_1;
  assign LUT_mem_MPORT_277_data = {1'h1,push_id_temp};
  assign LUT_mem_MPORT_277_addr = 6'h14;
  assign LUT_mem_MPORT_277_mask = 1'h1;
  assign LUT_mem_MPORT_277_en = _T_1015 ? 1'h0 : _T_1017;
  assign LUT_mem_MPORT_278_data = LUT_mem_MPORT_279_data;
  assign LUT_mem_MPORT_278_addr = 6'h14;
  assign LUT_mem_MPORT_278_mask = 1'h1;
  assign LUT_mem_MPORT_278_en = _T_1015 ? 1'h0 : _GEN_11931;
  assign LUT_mem_MPORT_280_data = {1'h0,lo_21};
  assign LUT_mem_MPORT_280_addr = 6'h15;
  assign LUT_mem_MPORT_280_mask = 1'h1;
  assign LUT_mem_MPORT_280_en = dispatch_reg_21 | clear_21_1;
  assign LUT_mem_MPORT_282_data = {1'h1,push_id_temp};
  assign LUT_mem_MPORT_282_addr = 6'h15;
  assign LUT_mem_MPORT_282_mask = 1'h1;
  assign LUT_mem_MPORT_282_en = _T_1021 ? 1'h0 : _T_1023;
  assign LUT_mem_MPORT_283_data = LUT_mem_MPORT_284_data;
  assign LUT_mem_MPORT_283_addr = 6'h15;
  assign LUT_mem_MPORT_283_mask = 1'h1;
  assign LUT_mem_MPORT_283_en = _T_1021 ? 1'h0 : _GEN_11956;
  assign LUT_mem_MPORT_285_data = {1'h0,lo_22};
  assign LUT_mem_MPORT_285_addr = 6'h16;
  assign LUT_mem_MPORT_285_mask = 1'h1;
  assign LUT_mem_MPORT_285_en = dispatch_reg_22 | clear_22_1;
  assign LUT_mem_MPORT_287_data = {1'h1,push_id_temp};
  assign LUT_mem_MPORT_287_addr = 6'h16;
  assign LUT_mem_MPORT_287_mask = 1'h1;
  assign LUT_mem_MPORT_287_en = _T_1027 ? 1'h0 : _T_1029;
  assign LUT_mem_MPORT_288_data = LUT_mem_MPORT_289_data;
  assign LUT_mem_MPORT_288_addr = 6'h16;
  assign LUT_mem_MPORT_288_mask = 1'h1;
  assign LUT_mem_MPORT_288_en = _T_1027 ? 1'h0 : _GEN_11981;
  assign LUT_mem_MPORT_290_data = {1'h0,lo_23};
  assign LUT_mem_MPORT_290_addr = 6'h17;
  assign LUT_mem_MPORT_290_mask = 1'h1;
  assign LUT_mem_MPORT_290_en = dispatch_reg_23 | clear_23_1;
  assign LUT_mem_MPORT_292_data = {1'h1,push_id_temp};
  assign LUT_mem_MPORT_292_addr = 6'h17;
  assign LUT_mem_MPORT_292_mask = 1'h1;
  assign LUT_mem_MPORT_292_en = _T_1033 ? 1'h0 : _T_1035;
  assign LUT_mem_MPORT_293_data = LUT_mem_MPORT_294_data;
  assign LUT_mem_MPORT_293_addr = 6'h17;
  assign LUT_mem_MPORT_293_mask = 1'h1;
  assign LUT_mem_MPORT_293_en = _T_1033 ? 1'h0 : _GEN_12006;
  assign LUT_mem_MPORT_295_data = {1'h0,lo_24};
  assign LUT_mem_MPORT_295_addr = 6'h18;
  assign LUT_mem_MPORT_295_mask = 1'h1;
  assign LUT_mem_MPORT_295_en = dispatch_reg_24 | clear_24_1;
  assign LUT_mem_MPORT_297_data = {1'h1,push_id_temp};
  assign LUT_mem_MPORT_297_addr = 6'h18;
  assign LUT_mem_MPORT_297_mask = 1'h1;
  assign LUT_mem_MPORT_297_en = _T_1039 ? 1'h0 : _T_1041;
  assign LUT_mem_MPORT_298_data = LUT_mem_MPORT_299_data;
  assign LUT_mem_MPORT_298_addr = 6'h18;
  assign LUT_mem_MPORT_298_mask = 1'h1;
  assign LUT_mem_MPORT_298_en = _T_1039 ? 1'h0 : _GEN_12031;
  assign LUT_mem_MPORT_300_data = {1'h0,lo_25};
  assign LUT_mem_MPORT_300_addr = 6'h19;
  assign LUT_mem_MPORT_300_mask = 1'h1;
  assign LUT_mem_MPORT_300_en = dispatch_reg_25 | clear_25_1;
  assign LUT_mem_MPORT_302_data = {1'h1,push_id_temp};
  assign LUT_mem_MPORT_302_addr = 6'h19;
  assign LUT_mem_MPORT_302_mask = 1'h1;
  assign LUT_mem_MPORT_302_en = _T_1045 ? 1'h0 : _T_1047;
  assign LUT_mem_MPORT_303_data = LUT_mem_MPORT_304_data;
  assign LUT_mem_MPORT_303_addr = 6'h19;
  assign LUT_mem_MPORT_303_mask = 1'h1;
  assign LUT_mem_MPORT_303_en = _T_1045 ? 1'h0 : _GEN_12056;
  assign LUT_mem_MPORT_305_data = {1'h0,lo_26};
  assign LUT_mem_MPORT_305_addr = 6'h1a;
  assign LUT_mem_MPORT_305_mask = 1'h1;
  assign LUT_mem_MPORT_305_en = dispatch_reg_26 | clear_26_1;
  assign LUT_mem_MPORT_307_data = {1'h1,push_id_temp};
  assign LUT_mem_MPORT_307_addr = 6'h1a;
  assign LUT_mem_MPORT_307_mask = 1'h1;
  assign LUT_mem_MPORT_307_en = _T_1051 ? 1'h0 : _T_1053;
  assign LUT_mem_MPORT_308_data = LUT_mem_MPORT_309_data;
  assign LUT_mem_MPORT_308_addr = 6'h1a;
  assign LUT_mem_MPORT_308_mask = 1'h1;
  assign LUT_mem_MPORT_308_en = _T_1051 ? 1'h0 : _GEN_12081;
  assign LUT_mem_MPORT_310_data = {1'h0,lo_27};
  assign LUT_mem_MPORT_310_addr = 6'h1b;
  assign LUT_mem_MPORT_310_mask = 1'h1;
  assign LUT_mem_MPORT_310_en = dispatch_reg_27 | clear_27_1;
  assign LUT_mem_MPORT_312_data = {1'h1,push_id_temp};
  assign LUT_mem_MPORT_312_addr = 6'h1b;
  assign LUT_mem_MPORT_312_mask = 1'h1;
  assign LUT_mem_MPORT_312_en = _T_1057 ? 1'h0 : _T_1059;
  assign LUT_mem_MPORT_313_data = LUT_mem_MPORT_314_data;
  assign LUT_mem_MPORT_313_addr = 6'h1b;
  assign LUT_mem_MPORT_313_mask = 1'h1;
  assign LUT_mem_MPORT_313_en = _T_1057 ? 1'h0 : _GEN_12106;
  assign LUT_mem_MPORT_315_data = {1'h0,lo_28};
  assign LUT_mem_MPORT_315_addr = 6'h1c;
  assign LUT_mem_MPORT_315_mask = 1'h1;
  assign LUT_mem_MPORT_315_en = dispatch_reg_28 | clear_28_1;
  assign LUT_mem_MPORT_317_data = {1'h1,push_id_temp};
  assign LUT_mem_MPORT_317_addr = 6'h1c;
  assign LUT_mem_MPORT_317_mask = 1'h1;
  assign LUT_mem_MPORT_317_en = _T_1063 ? 1'h0 : _T_1065;
  assign LUT_mem_MPORT_318_data = LUT_mem_MPORT_319_data;
  assign LUT_mem_MPORT_318_addr = 6'h1c;
  assign LUT_mem_MPORT_318_mask = 1'h1;
  assign LUT_mem_MPORT_318_en = _T_1063 ? 1'h0 : _GEN_12131;
  assign LUT_mem_MPORT_320_data = {1'h0,lo_29};
  assign LUT_mem_MPORT_320_addr = 6'h1d;
  assign LUT_mem_MPORT_320_mask = 1'h1;
  assign LUT_mem_MPORT_320_en = dispatch_reg_29 | clear_29_1;
  assign LUT_mem_MPORT_322_data = {1'h1,push_id_temp};
  assign LUT_mem_MPORT_322_addr = 6'h1d;
  assign LUT_mem_MPORT_322_mask = 1'h1;
  assign LUT_mem_MPORT_322_en = _T_1069 ? 1'h0 : _T_1071;
  assign LUT_mem_MPORT_323_data = LUT_mem_MPORT_324_data;
  assign LUT_mem_MPORT_323_addr = 6'h1d;
  assign LUT_mem_MPORT_323_mask = 1'h1;
  assign LUT_mem_MPORT_323_en = _T_1069 ? 1'h0 : _GEN_12156;
  assign LUT_mem_MPORT_325_data = {1'h0,lo_30};
  assign LUT_mem_MPORT_325_addr = 6'h1e;
  assign LUT_mem_MPORT_325_mask = 1'h1;
  assign LUT_mem_MPORT_325_en = dispatch_reg_30 | clear_30_1;
  assign LUT_mem_MPORT_327_data = {1'h1,push_id_temp};
  assign LUT_mem_MPORT_327_addr = 6'h1e;
  assign LUT_mem_MPORT_327_mask = 1'h1;
  assign LUT_mem_MPORT_327_en = _T_1075 ? 1'h0 : _T_1077;
  assign LUT_mem_MPORT_328_data = LUT_mem_MPORT_329_data;
  assign LUT_mem_MPORT_328_addr = 6'h1e;
  assign LUT_mem_MPORT_328_mask = 1'h1;
  assign LUT_mem_MPORT_328_en = _T_1075 ? 1'h0 : _GEN_12181;
  assign LUT_mem_MPORT_330_data = {1'h0,lo_31};
  assign LUT_mem_MPORT_330_addr = 6'h1f;
  assign LUT_mem_MPORT_330_mask = 1'h1;
  assign LUT_mem_MPORT_330_en = dispatch_reg_31 | clear_31_1;
  assign LUT_mem_MPORT_332_data = {1'h1,push_id_temp};
  assign LUT_mem_MPORT_332_addr = 6'h1f;
  assign LUT_mem_MPORT_332_mask = 1'h1;
  assign LUT_mem_MPORT_332_en = _T_1081 ? 1'h0 : _T_1083;
  assign LUT_mem_MPORT_333_data = LUT_mem_MPORT_334_data;
  assign LUT_mem_MPORT_333_addr = 6'h1f;
  assign LUT_mem_MPORT_333_mask = 1'h1;
  assign LUT_mem_MPORT_333_en = _T_1081 ? 1'h0 : _GEN_12206;
  assign LUT_mem_MPORT_335_data = {1'h0,lo_32};
  assign LUT_mem_MPORT_335_addr = 6'h20;
  assign LUT_mem_MPORT_335_mask = 1'h1;
  assign LUT_mem_MPORT_335_en = dispatch_reg_32 | clear_32_1;
  assign LUT_mem_MPORT_337_data = {1'h1,push_id_temp};
  assign LUT_mem_MPORT_337_addr = 6'h20;
  assign LUT_mem_MPORT_337_mask = 1'h1;
  assign LUT_mem_MPORT_337_en = _T_1087 ? 1'h0 : _T_1089;
  assign LUT_mem_MPORT_338_data = LUT_mem_MPORT_339_data;
  assign LUT_mem_MPORT_338_addr = 6'h20;
  assign LUT_mem_MPORT_338_mask = 1'h1;
  assign LUT_mem_MPORT_338_en = _T_1087 ? 1'h0 : _GEN_12231;
  assign LUT_mem_MPORT_340_data = {1'h0,lo_33};
  assign LUT_mem_MPORT_340_addr = 6'h21;
  assign LUT_mem_MPORT_340_mask = 1'h1;
  assign LUT_mem_MPORT_340_en = dispatch_reg_33 | clear_33_1;
  assign LUT_mem_MPORT_342_data = {1'h1,push_id_temp};
  assign LUT_mem_MPORT_342_addr = 6'h21;
  assign LUT_mem_MPORT_342_mask = 1'h1;
  assign LUT_mem_MPORT_342_en = _T_1093 ? 1'h0 : _T_1095;
  assign LUT_mem_MPORT_343_data = LUT_mem_MPORT_344_data;
  assign LUT_mem_MPORT_343_addr = 6'h21;
  assign LUT_mem_MPORT_343_mask = 1'h1;
  assign LUT_mem_MPORT_343_en = _T_1093 ? 1'h0 : _GEN_12256;
  assign LUT_mem_MPORT_345_data = {1'h0,lo_34};
  assign LUT_mem_MPORT_345_addr = 6'h22;
  assign LUT_mem_MPORT_345_mask = 1'h1;
  assign LUT_mem_MPORT_345_en = dispatch_reg_34 | clear_34_1;
  assign LUT_mem_MPORT_347_data = {1'h1,push_id_temp};
  assign LUT_mem_MPORT_347_addr = 6'h22;
  assign LUT_mem_MPORT_347_mask = 1'h1;
  assign LUT_mem_MPORT_347_en = _T_1099 ? 1'h0 : _T_1101;
  assign LUT_mem_MPORT_348_data = LUT_mem_MPORT_349_data;
  assign LUT_mem_MPORT_348_addr = 6'h22;
  assign LUT_mem_MPORT_348_mask = 1'h1;
  assign LUT_mem_MPORT_348_en = _T_1099 ? 1'h0 : _GEN_12281;
  assign io_ray_id_pop_out = pop_ray_id_2; // @[lut_35.scala 5170:46]
  assign io_hitT_out = pop_hitT_2; // @[lut_35.scala 5171:56]
  assign io_pop_0 = pop_0_1; // @[lut_35.scala 5128:57]
  assign io_pop_1 = pop_1_1; // @[lut_35.scala 5129:57]
  assign io_pop_2 = pop_2_1; // @[lut_35.scala 5130:57]
  assign io_pop_3 = pop_3_1; // @[lut_35.scala 5131:57]
  assign io_pop_4 = pop_4_1; // @[lut_35.scala 5132:57]
  assign io_pop_5 = pop_5_1; // @[lut_35.scala 5133:57]
  assign io_pop_6 = pop_6_1; // @[lut_35.scala 5134:57]
  assign io_pop_7 = pop_7_1; // @[lut_35.scala 5135:57]
  assign io_pop_8 = pop_8_1; // @[lut_35.scala 5136:57]
  assign io_pop_9 = pop_9_1; // @[lut_35.scala 5137:57]
  assign io_pop_10 = pop_10_1; // @[lut_35.scala 5139:58]
  assign io_pop_11 = pop_11_1; // @[lut_35.scala 5140:58]
  assign io_pop_12 = pop_12_1; // @[lut_35.scala 5141:58]
  assign io_pop_13 = pop_13_1; // @[lut_35.scala 5142:58]
  assign io_pop_14 = pop_14_1; // @[lut_35.scala 5143:58]
  assign io_pop_15 = pop_15_1; // @[lut_35.scala 5144:58]
  assign io_pop_16 = pop_16_1; // @[lut_35.scala 5145:58]
  assign io_pop_17 = pop_17_1; // @[lut_35.scala 5146:58]
  assign io_pop_18 = pop_18_1; // @[lut_35.scala 5147:58]
  assign io_pop_19 = pop_19_1; // @[lut_35.scala 5148:58]
  assign io_pop_20 = pop_20_1; // @[lut_35.scala 5150:58]
  assign io_pop_21 = pop_21_1; // @[lut_35.scala 5151:58]
  assign io_pop_22 = pop_22_1; // @[lut_35.scala 5152:58]
  assign io_pop_23 = pop_23_1; // @[lut_35.scala 5153:58]
  assign io_pop_24 = pop_24_1; // @[lut_35.scala 5154:58]
  assign io_pop_25 = pop_25_1; // @[lut_35.scala 5155:58]
  assign io_pop_26 = pop_26_1; // @[lut_35.scala 5156:58]
  assign io_pop_27 = pop_27_1; // @[lut_35.scala 5157:58]
  assign io_pop_28 = pop_28_1; // @[lut_35.scala 5158:58]
  assign io_pop_29 = pop_29_1; // @[lut_35.scala 5159:58]
  assign io_pop_30 = pop_30_1; // @[lut_35.scala 5161:58]
  assign io_pop_31 = pop_31_1; // @[lut_35.scala 5162:58]
  assign io_pop_32 = pop_32_1; // @[lut_35.scala 5163:58]
  assign io_pop_33 = pop_33_1; // @[lut_35.scala 5164:58]
  assign io_pop_34 = pop_34_1; // @[lut_35.scala 5165:58]
  assign io_pop_en = pop_valid_2; // @[lut_35.scala 5169:55]
  assign io_push_0 = push_0_1; // @[lut_35.scala 3455:51]
  assign io_push_1 = push_1_1; // @[lut_35.scala 3456:51]
  assign io_push_2 = push_2_1; // @[lut_35.scala 3457:51]
  assign io_push_3 = push_3_1; // @[lut_35.scala 3458:51]
  assign io_push_4 = push_4_1; // @[lut_35.scala 3459:51]
  assign io_push_5 = push_5_1; // @[lut_35.scala 3460:51]
  assign io_push_6 = push_6_1; // @[lut_35.scala 3461:51]
  assign io_push_7 = push_7_1; // @[lut_35.scala 3462:51]
  assign io_push_8 = push_8_1; // @[lut_35.scala 3463:51]
  assign io_push_9 = push_9_1; // @[lut_35.scala 3464:51]
  assign io_push_10 = push_10_1; // @[lut_35.scala 3465:52]
  assign io_push_11 = push_11_1; // @[lut_35.scala 3466:52]
  assign io_push_12 = push_12_1; // @[lut_35.scala 3467:52]
  assign io_push_13 = push_13_1; // @[lut_35.scala 3468:52]
  assign io_push_14 = push_14_1; // @[lut_35.scala 3469:52]
  assign io_push_15 = push_15_1; // @[lut_35.scala 3470:52]
  assign io_push_16 = push_16_1; // @[lut_35.scala 3471:52]
  assign io_push_17 = push_17_1; // @[lut_35.scala 3472:52]
  assign io_push_18 = push_18_1; // @[lut_35.scala 3473:52]
  assign io_push_19 = push_19_1; // @[lut_35.scala 3474:52]
  assign io_push_20 = push_20_1; // @[lut_35.scala 3475:52]
  assign io_push_21 = push_21_1; // @[lut_35.scala 3476:52]
  assign io_push_22 = push_22_1; // @[lut_35.scala 3477:52]
  assign io_push_23 = push_23_1; // @[lut_35.scala 3478:52]
  assign io_push_24 = push_24_1; // @[lut_35.scala 3479:52]
  assign io_push_25 = push_25_1; // @[lut_35.scala 3480:52]
  assign io_push_26 = push_26_1; // @[lut_35.scala 3481:52]
  assign io_push_27 = push_27_1; // @[lut_35.scala 3482:52]
  assign io_push_28 = push_28_1; // @[lut_35.scala 3483:52]
  assign io_push_29 = push_29_1; // @[lut_35.scala 3484:52]
  assign io_push_30 = push_30_1; // @[lut_35.scala 3485:52]
  assign io_push_31 = push_31_1; // @[lut_35.scala 3486:52]
  assign io_push_32 = push_32_1; // @[lut_35.scala 3487:52]
  assign io_push_33 = push_33_1; // @[lut_35.scala 3488:52]
  assign io_push_34 = push_34_1; // @[lut_35.scala 3489:52]
  assign io_clear_0 = clear_0_1; // @[lut_35.scala 6713:59]
  assign io_clear_1 = clear_1_1; // @[lut_35.scala 6714:59]
  assign io_clear_2 = clear_2_1; // @[lut_35.scala 6715:59]
  assign io_clear_3 = clear_3_1; // @[lut_35.scala 6716:59]
  assign io_clear_4 = clear_4_1; // @[lut_35.scala 6717:59]
  assign io_clear_5 = clear_5_1; // @[lut_35.scala 6718:59]
  assign io_clear_6 = clear_6_1; // @[lut_35.scala 6719:59]
  assign io_clear_7 = clear_7_1; // @[lut_35.scala 6720:59]
  assign io_clear_8 = clear_8_1; // @[lut_35.scala 6721:59]
  assign io_clear_9 = clear_9_1; // @[lut_35.scala 6722:59]
  assign io_clear_10 = clear_10_1; // @[lut_35.scala 6724:60]
  assign io_clear_11 = clear_11_1; // @[lut_35.scala 6725:60]
  assign io_clear_12 = clear_12_1; // @[lut_35.scala 6726:60]
  assign io_clear_13 = clear_13_1; // @[lut_35.scala 6727:60]
  assign io_clear_14 = clear_14_1; // @[lut_35.scala 6728:60]
  assign io_clear_15 = clear_15_1; // @[lut_35.scala 6729:60]
  assign io_clear_16 = clear_16_1; // @[lut_35.scala 6730:60]
  assign io_clear_17 = clear_17_1; // @[lut_35.scala 6731:60]
  assign io_clear_18 = clear_18_1; // @[lut_35.scala 6732:60]
  assign io_clear_19 = clear_19_1; // @[lut_35.scala 6733:60]
  assign io_clear_20 = clear_20_1; // @[lut_35.scala 6735:60]
  assign io_clear_21 = clear_21_1; // @[lut_35.scala 6736:60]
  assign io_clear_22 = clear_22_1; // @[lut_35.scala 6737:60]
  assign io_clear_23 = clear_23_1; // @[lut_35.scala 6738:60]
  assign io_clear_24 = clear_24_1; // @[lut_35.scala 6739:60]
  assign io_clear_25 = clear_25_1; // @[lut_35.scala 6740:60]
  assign io_clear_26 = clear_26_1; // @[lut_35.scala 6741:60]
  assign io_clear_27 = clear_27_1; // @[lut_35.scala 6742:60]
  assign io_clear_28 = clear_28_1; // @[lut_35.scala 6743:60]
  assign io_clear_29 = clear_29_1; // @[lut_35.scala 6744:60]
  assign io_clear_30 = clear_30_1; // @[lut_35.scala 6746:60]
  assign io_clear_31 = clear_31_1; // @[lut_35.scala 6747:60]
  assign io_clear_32 = clear_32_1; // @[lut_35.scala 6748:60]
  assign io_clear_33 = clear_33_1; // @[lut_35.scala 6749:60]
  assign io_clear_34 = clear_34_1; // @[lut_35.scala 6750:60]
  assign io_push_en = push_valid_2; // @[lut_35.scala 3492:50]
  assign io_no_match = no_match_2; // @[lut_35.scala 3648:41]
  always @(posedge clock) begin
    if(LUT_mem_MPORT_175_en & LUT_mem_MPORT_175_mask) begin
      LUT_mem[LUT_mem_MPORT_175_addr] <= LUT_mem_MPORT_175_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_177_en & LUT_mem_MPORT_177_mask) begin
      LUT_mem[LUT_mem_MPORT_177_addr] <= LUT_mem_MPORT_177_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_178_en & LUT_mem_MPORT_178_mask) begin
      LUT_mem[LUT_mem_MPORT_178_addr] <= LUT_mem_MPORT_178_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_180_en & LUT_mem_MPORT_180_mask) begin
      LUT_mem[LUT_mem_MPORT_180_addr] <= LUT_mem_MPORT_180_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_182_en & LUT_mem_MPORT_182_mask) begin
      LUT_mem[LUT_mem_MPORT_182_addr] <= LUT_mem_MPORT_182_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_183_en & LUT_mem_MPORT_183_mask) begin
      LUT_mem[LUT_mem_MPORT_183_addr] <= LUT_mem_MPORT_183_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_185_en & LUT_mem_MPORT_185_mask) begin
      LUT_mem[LUT_mem_MPORT_185_addr] <= LUT_mem_MPORT_185_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_187_en & LUT_mem_MPORT_187_mask) begin
      LUT_mem[LUT_mem_MPORT_187_addr] <= LUT_mem_MPORT_187_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_188_en & LUT_mem_MPORT_188_mask) begin
      LUT_mem[LUT_mem_MPORT_188_addr] <= LUT_mem_MPORT_188_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_190_en & LUT_mem_MPORT_190_mask) begin
      LUT_mem[LUT_mem_MPORT_190_addr] <= LUT_mem_MPORT_190_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_192_en & LUT_mem_MPORT_192_mask) begin
      LUT_mem[LUT_mem_MPORT_192_addr] <= LUT_mem_MPORT_192_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_193_en & LUT_mem_MPORT_193_mask) begin
      LUT_mem[LUT_mem_MPORT_193_addr] <= LUT_mem_MPORT_193_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_195_en & LUT_mem_MPORT_195_mask) begin
      LUT_mem[LUT_mem_MPORT_195_addr] <= LUT_mem_MPORT_195_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_197_en & LUT_mem_MPORT_197_mask) begin
      LUT_mem[LUT_mem_MPORT_197_addr] <= LUT_mem_MPORT_197_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_198_en & LUT_mem_MPORT_198_mask) begin
      LUT_mem[LUT_mem_MPORT_198_addr] <= LUT_mem_MPORT_198_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_200_en & LUT_mem_MPORT_200_mask) begin
      LUT_mem[LUT_mem_MPORT_200_addr] <= LUT_mem_MPORT_200_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_202_en & LUT_mem_MPORT_202_mask) begin
      LUT_mem[LUT_mem_MPORT_202_addr] <= LUT_mem_MPORT_202_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_203_en & LUT_mem_MPORT_203_mask) begin
      LUT_mem[LUT_mem_MPORT_203_addr] <= LUT_mem_MPORT_203_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_205_en & LUT_mem_MPORT_205_mask) begin
      LUT_mem[LUT_mem_MPORT_205_addr] <= LUT_mem_MPORT_205_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_207_en & LUT_mem_MPORT_207_mask) begin
      LUT_mem[LUT_mem_MPORT_207_addr] <= LUT_mem_MPORT_207_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_208_en & LUT_mem_MPORT_208_mask) begin
      LUT_mem[LUT_mem_MPORT_208_addr] <= LUT_mem_MPORT_208_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_210_en & LUT_mem_MPORT_210_mask) begin
      LUT_mem[LUT_mem_MPORT_210_addr] <= LUT_mem_MPORT_210_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_212_en & LUT_mem_MPORT_212_mask) begin
      LUT_mem[LUT_mem_MPORT_212_addr] <= LUT_mem_MPORT_212_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_213_en & LUT_mem_MPORT_213_mask) begin
      LUT_mem[LUT_mem_MPORT_213_addr] <= LUT_mem_MPORT_213_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_215_en & LUT_mem_MPORT_215_mask) begin
      LUT_mem[LUT_mem_MPORT_215_addr] <= LUT_mem_MPORT_215_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_217_en & LUT_mem_MPORT_217_mask) begin
      LUT_mem[LUT_mem_MPORT_217_addr] <= LUT_mem_MPORT_217_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_218_en & LUT_mem_MPORT_218_mask) begin
      LUT_mem[LUT_mem_MPORT_218_addr] <= LUT_mem_MPORT_218_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_220_en & LUT_mem_MPORT_220_mask) begin
      LUT_mem[LUT_mem_MPORT_220_addr] <= LUT_mem_MPORT_220_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_222_en & LUT_mem_MPORT_222_mask) begin
      LUT_mem[LUT_mem_MPORT_222_addr] <= LUT_mem_MPORT_222_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_223_en & LUT_mem_MPORT_223_mask) begin
      LUT_mem[LUT_mem_MPORT_223_addr] <= LUT_mem_MPORT_223_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_225_en & LUT_mem_MPORT_225_mask) begin
      LUT_mem[LUT_mem_MPORT_225_addr] <= LUT_mem_MPORT_225_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_227_en & LUT_mem_MPORT_227_mask) begin
      LUT_mem[LUT_mem_MPORT_227_addr] <= LUT_mem_MPORT_227_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_228_en & LUT_mem_MPORT_228_mask) begin
      LUT_mem[LUT_mem_MPORT_228_addr] <= LUT_mem_MPORT_228_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_230_en & LUT_mem_MPORT_230_mask) begin
      LUT_mem[LUT_mem_MPORT_230_addr] <= LUT_mem_MPORT_230_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_232_en & LUT_mem_MPORT_232_mask) begin
      LUT_mem[LUT_mem_MPORT_232_addr] <= LUT_mem_MPORT_232_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_233_en & LUT_mem_MPORT_233_mask) begin
      LUT_mem[LUT_mem_MPORT_233_addr] <= LUT_mem_MPORT_233_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_235_en & LUT_mem_MPORT_235_mask) begin
      LUT_mem[LUT_mem_MPORT_235_addr] <= LUT_mem_MPORT_235_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_237_en & LUT_mem_MPORT_237_mask) begin
      LUT_mem[LUT_mem_MPORT_237_addr] <= LUT_mem_MPORT_237_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_238_en & LUT_mem_MPORT_238_mask) begin
      LUT_mem[LUT_mem_MPORT_238_addr] <= LUT_mem_MPORT_238_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_240_en & LUT_mem_MPORT_240_mask) begin
      LUT_mem[LUT_mem_MPORT_240_addr] <= LUT_mem_MPORT_240_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_242_en & LUT_mem_MPORT_242_mask) begin
      LUT_mem[LUT_mem_MPORT_242_addr] <= LUT_mem_MPORT_242_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_243_en & LUT_mem_MPORT_243_mask) begin
      LUT_mem[LUT_mem_MPORT_243_addr] <= LUT_mem_MPORT_243_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_245_en & LUT_mem_MPORT_245_mask) begin
      LUT_mem[LUT_mem_MPORT_245_addr] <= LUT_mem_MPORT_245_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_247_en & LUT_mem_MPORT_247_mask) begin
      LUT_mem[LUT_mem_MPORT_247_addr] <= LUT_mem_MPORT_247_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_248_en & LUT_mem_MPORT_248_mask) begin
      LUT_mem[LUT_mem_MPORT_248_addr] <= LUT_mem_MPORT_248_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_250_en & LUT_mem_MPORT_250_mask) begin
      LUT_mem[LUT_mem_MPORT_250_addr] <= LUT_mem_MPORT_250_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_252_en & LUT_mem_MPORT_252_mask) begin
      LUT_mem[LUT_mem_MPORT_252_addr] <= LUT_mem_MPORT_252_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_253_en & LUT_mem_MPORT_253_mask) begin
      LUT_mem[LUT_mem_MPORT_253_addr] <= LUT_mem_MPORT_253_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_255_en & LUT_mem_MPORT_255_mask) begin
      LUT_mem[LUT_mem_MPORT_255_addr] <= LUT_mem_MPORT_255_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_257_en & LUT_mem_MPORT_257_mask) begin
      LUT_mem[LUT_mem_MPORT_257_addr] <= LUT_mem_MPORT_257_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_258_en & LUT_mem_MPORT_258_mask) begin
      LUT_mem[LUT_mem_MPORT_258_addr] <= LUT_mem_MPORT_258_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_260_en & LUT_mem_MPORT_260_mask) begin
      LUT_mem[LUT_mem_MPORT_260_addr] <= LUT_mem_MPORT_260_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_262_en & LUT_mem_MPORT_262_mask) begin
      LUT_mem[LUT_mem_MPORT_262_addr] <= LUT_mem_MPORT_262_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_263_en & LUT_mem_MPORT_263_mask) begin
      LUT_mem[LUT_mem_MPORT_263_addr] <= LUT_mem_MPORT_263_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_265_en & LUT_mem_MPORT_265_mask) begin
      LUT_mem[LUT_mem_MPORT_265_addr] <= LUT_mem_MPORT_265_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_267_en & LUT_mem_MPORT_267_mask) begin
      LUT_mem[LUT_mem_MPORT_267_addr] <= LUT_mem_MPORT_267_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_268_en & LUT_mem_MPORT_268_mask) begin
      LUT_mem[LUT_mem_MPORT_268_addr] <= LUT_mem_MPORT_268_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_270_en & LUT_mem_MPORT_270_mask) begin
      LUT_mem[LUT_mem_MPORT_270_addr] <= LUT_mem_MPORT_270_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_272_en & LUT_mem_MPORT_272_mask) begin
      LUT_mem[LUT_mem_MPORT_272_addr] <= LUT_mem_MPORT_272_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_273_en & LUT_mem_MPORT_273_mask) begin
      LUT_mem[LUT_mem_MPORT_273_addr] <= LUT_mem_MPORT_273_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_275_en & LUT_mem_MPORT_275_mask) begin
      LUT_mem[LUT_mem_MPORT_275_addr] <= LUT_mem_MPORT_275_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_277_en & LUT_mem_MPORT_277_mask) begin
      LUT_mem[LUT_mem_MPORT_277_addr] <= LUT_mem_MPORT_277_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_278_en & LUT_mem_MPORT_278_mask) begin
      LUT_mem[LUT_mem_MPORT_278_addr] <= LUT_mem_MPORT_278_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_280_en & LUT_mem_MPORT_280_mask) begin
      LUT_mem[LUT_mem_MPORT_280_addr] <= LUT_mem_MPORT_280_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_282_en & LUT_mem_MPORT_282_mask) begin
      LUT_mem[LUT_mem_MPORT_282_addr] <= LUT_mem_MPORT_282_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_283_en & LUT_mem_MPORT_283_mask) begin
      LUT_mem[LUT_mem_MPORT_283_addr] <= LUT_mem_MPORT_283_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_285_en & LUT_mem_MPORT_285_mask) begin
      LUT_mem[LUT_mem_MPORT_285_addr] <= LUT_mem_MPORT_285_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_287_en & LUT_mem_MPORT_287_mask) begin
      LUT_mem[LUT_mem_MPORT_287_addr] <= LUT_mem_MPORT_287_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_288_en & LUT_mem_MPORT_288_mask) begin
      LUT_mem[LUT_mem_MPORT_288_addr] <= LUT_mem_MPORT_288_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_290_en & LUT_mem_MPORT_290_mask) begin
      LUT_mem[LUT_mem_MPORT_290_addr] <= LUT_mem_MPORT_290_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_292_en & LUT_mem_MPORT_292_mask) begin
      LUT_mem[LUT_mem_MPORT_292_addr] <= LUT_mem_MPORT_292_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_293_en & LUT_mem_MPORT_293_mask) begin
      LUT_mem[LUT_mem_MPORT_293_addr] <= LUT_mem_MPORT_293_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_295_en & LUT_mem_MPORT_295_mask) begin
      LUT_mem[LUT_mem_MPORT_295_addr] <= LUT_mem_MPORT_295_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_297_en & LUT_mem_MPORT_297_mask) begin
      LUT_mem[LUT_mem_MPORT_297_addr] <= LUT_mem_MPORT_297_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_298_en & LUT_mem_MPORT_298_mask) begin
      LUT_mem[LUT_mem_MPORT_298_addr] <= LUT_mem_MPORT_298_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_300_en & LUT_mem_MPORT_300_mask) begin
      LUT_mem[LUT_mem_MPORT_300_addr] <= LUT_mem_MPORT_300_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_302_en & LUT_mem_MPORT_302_mask) begin
      LUT_mem[LUT_mem_MPORT_302_addr] <= LUT_mem_MPORT_302_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_303_en & LUT_mem_MPORT_303_mask) begin
      LUT_mem[LUT_mem_MPORT_303_addr] <= LUT_mem_MPORT_303_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_305_en & LUT_mem_MPORT_305_mask) begin
      LUT_mem[LUT_mem_MPORT_305_addr] <= LUT_mem_MPORT_305_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_307_en & LUT_mem_MPORT_307_mask) begin
      LUT_mem[LUT_mem_MPORT_307_addr] <= LUT_mem_MPORT_307_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_308_en & LUT_mem_MPORT_308_mask) begin
      LUT_mem[LUT_mem_MPORT_308_addr] <= LUT_mem_MPORT_308_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_310_en & LUT_mem_MPORT_310_mask) begin
      LUT_mem[LUT_mem_MPORT_310_addr] <= LUT_mem_MPORT_310_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_312_en & LUT_mem_MPORT_312_mask) begin
      LUT_mem[LUT_mem_MPORT_312_addr] <= LUT_mem_MPORT_312_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_313_en & LUT_mem_MPORT_313_mask) begin
      LUT_mem[LUT_mem_MPORT_313_addr] <= LUT_mem_MPORT_313_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_315_en & LUT_mem_MPORT_315_mask) begin
      LUT_mem[LUT_mem_MPORT_315_addr] <= LUT_mem_MPORT_315_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_317_en & LUT_mem_MPORT_317_mask) begin
      LUT_mem[LUT_mem_MPORT_317_addr] <= LUT_mem_MPORT_317_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_318_en & LUT_mem_MPORT_318_mask) begin
      LUT_mem[LUT_mem_MPORT_318_addr] <= LUT_mem_MPORT_318_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_320_en & LUT_mem_MPORT_320_mask) begin
      LUT_mem[LUT_mem_MPORT_320_addr] <= LUT_mem_MPORT_320_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_322_en & LUT_mem_MPORT_322_mask) begin
      LUT_mem[LUT_mem_MPORT_322_addr] <= LUT_mem_MPORT_322_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_323_en & LUT_mem_MPORT_323_mask) begin
      LUT_mem[LUT_mem_MPORT_323_addr] <= LUT_mem_MPORT_323_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_325_en & LUT_mem_MPORT_325_mask) begin
      LUT_mem[LUT_mem_MPORT_325_addr] <= LUT_mem_MPORT_325_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_327_en & LUT_mem_MPORT_327_mask) begin
      LUT_mem[LUT_mem_MPORT_327_addr] <= LUT_mem_MPORT_327_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_328_en & LUT_mem_MPORT_328_mask) begin
      LUT_mem[LUT_mem_MPORT_328_addr] <= LUT_mem_MPORT_328_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_330_en & LUT_mem_MPORT_330_mask) begin
      LUT_mem[LUT_mem_MPORT_330_addr] <= LUT_mem_MPORT_330_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_332_en & LUT_mem_MPORT_332_mask) begin
      LUT_mem[LUT_mem_MPORT_332_addr] <= LUT_mem_MPORT_332_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_333_en & LUT_mem_MPORT_333_mask) begin
      LUT_mem[LUT_mem_MPORT_333_addr] <= LUT_mem_MPORT_333_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_335_en & LUT_mem_MPORT_335_mask) begin
      LUT_mem[LUT_mem_MPORT_335_addr] <= LUT_mem_MPORT_335_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_337_en & LUT_mem_MPORT_337_mask) begin
      LUT_mem[LUT_mem_MPORT_337_addr] <= LUT_mem_MPORT_337_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_338_en & LUT_mem_MPORT_338_mask) begin
      LUT_mem[LUT_mem_MPORT_338_addr] <= LUT_mem_MPORT_338_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_340_en & LUT_mem_MPORT_340_mask) begin
      LUT_mem[LUT_mem_MPORT_340_addr] <= LUT_mem_MPORT_340_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_342_en & LUT_mem_MPORT_342_mask) begin
      LUT_mem[LUT_mem_MPORT_342_addr] <= LUT_mem_MPORT_342_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_343_en & LUT_mem_MPORT_343_mask) begin
      LUT_mem[LUT_mem_MPORT_343_addr] <= LUT_mem_MPORT_343_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_345_en & LUT_mem_MPORT_345_mask) begin
      LUT_mem[LUT_mem_MPORT_345_addr] <= LUT_mem_MPORT_345_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_347_en & LUT_mem_MPORT_347_mask) begin
      LUT_mem[LUT_mem_MPORT_347_addr] <= LUT_mem_MPORT_347_data; // @[lut_35.scala 216:26]
    end
    if(LUT_mem_MPORT_348_en & LUT_mem_MPORT_348_mask) begin
      LUT_mem[LUT_mem_MPORT_348_addr] <= LUT_mem_MPORT_348_data; // @[lut_35.scala 216:26]
    end
    if (reset) begin // @[lut_35.scala 217:30]
      read_stack0 <= 32'h0; // @[lut_35.scala 217:30]
    end else begin
      read_stack0 <= LUT_mem_MPORT_data[31:0]; // @[lut_35.scala 455:26]
    end
    if (reset) begin // @[lut_35.scala 218:30]
      read_stack1 <= 32'h0; // @[lut_35.scala 218:30]
    end else begin
      read_stack1 <= LUT_mem_MPORT_1_data[31:0]; // @[lut_35.scala 456:26]
    end
    if (reset) begin // @[lut_35.scala 219:30]
      read_stack2 <= 32'h0; // @[lut_35.scala 219:30]
    end else begin
      read_stack2 <= LUT_mem_MPORT_2_data[31:0]; // @[lut_35.scala 457:26]
    end
    if (reset) begin // @[lut_35.scala 220:30]
      read_stack3 <= 32'h0; // @[lut_35.scala 220:30]
    end else begin
      read_stack3 <= LUT_mem_MPORT_3_data[31:0]; // @[lut_35.scala 458:26]
    end
    if (reset) begin // @[lut_35.scala 221:30]
      read_stack4 <= 32'h0; // @[lut_35.scala 221:30]
    end else begin
      read_stack4 <= LUT_mem_MPORT_4_data[31:0]; // @[lut_35.scala 459:26]
    end
    if (reset) begin // @[lut_35.scala 222:30]
      read_stack5 <= 32'h0; // @[lut_35.scala 222:30]
    end else begin
      read_stack5 <= LUT_mem_MPORT_5_data[31:0]; // @[lut_35.scala 460:26]
    end
    if (reset) begin // @[lut_35.scala 223:30]
      read_stack6 <= 32'h0; // @[lut_35.scala 223:30]
    end else begin
      read_stack6 <= LUT_mem_MPORT_6_data[31:0]; // @[lut_35.scala 461:26]
    end
    if (reset) begin // @[lut_35.scala 224:30]
      read_stack7 <= 32'h0; // @[lut_35.scala 224:30]
    end else begin
      read_stack7 <= LUT_mem_MPORT_7_data[31:0]; // @[lut_35.scala 462:26]
    end
    if (reset) begin // @[lut_35.scala 225:30]
      read_stack8 <= 32'h0; // @[lut_35.scala 225:30]
    end else begin
      read_stack8 <= LUT_mem_MPORT_8_data[31:0]; // @[lut_35.scala 463:26]
    end
    if (reset) begin // @[lut_35.scala 226:30]
      read_stack9 <= 32'h0; // @[lut_35.scala 226:30]
    end else begin
      read_stack9 <= LUT_mem_MPORT_9_data[31:0]; // @[lut_35.scala 464:26]
    end
    if (reset) begin // @[lut_35.scala 227:31]
      read_stack10 <= 32'h0; // @[lut_35.scala 227:31]
    end else begin
      read_stack10 <= LUT_mem_MPORT_10_data[31:0]; // @[lut_35.scala 465:27]
    end
    if (reset) begin // @[lut_35.scala 228:31]
      read_stack11 <= 32'h0; // @[lut_35.scala 228:31]
    end else begin
      read_stack11 <= LUT_mem_MPORT_11_data[31:0]; // @[lut_35.scala 466:27]
    end
    if (reset) begin // @[lut_35.scala 229:31]
      read_stack12 <= 32'h0; // @[lut_35.scala 229:31]
    end else begin
      read_stack12 <= LUT_mem_MPORT_12_data[31:0]; // @[lut_35.scala 467:27]
    end
    if (reset) begin // @[lut_35.scala 230:31]
      read_stack13 <= 32'h0; // @[lut_35.scala 230:31]
    end else begin
      read_stack13 <= LUT_mem_MPORT_13_data[31:0]; // @[lut_35.scala 468:27]
    end
    if (reset) begin // @[lut_35.scala 231:31]
      read_stack14 <= 32'h0; // @[lut_35.scala 231:31]
    end else begin
      read_stack14 <= LUT_mem_MPORT_14_data[31:0]; // @[lut_35.scala 469:27]
    end
    if (reset) begin // @[lut_35.scala 232:31]
      read_stack15 <= 32'h0; // @[lut_35.scala 232:31]
    end else begin
      read_stack15 <= LUT_mem_MPORT_15_data[31:0]; // @[lut_35.scala 470:27]
    end
    if (reset) begin // @[lut_35.scala 233:31]
      read_stack16 <= 32'h0; // @[lut_35.scala 233:31]
    end else begin
      read_stack16 <= LUT_mem_MPORT_16_data[31:0]; // @[lut_35.scala 471:27]
    end
    if (reset) begin // @[lut_35.scala 234:31]
      read_stack17 <= 32'h0; // @[lut_35.scala 234:31]
    end else begin
      read_stack17 <= LUT_mem_MPORT_17_data[31:0]; // @[lut_35.scala 472:27]
    end
    if (reset) begin // @[lut_35.scala 235:31]
      read_stack18 <= 32'h0; // @[lut_35.scala 235:31]
    end else begin
      read_stack18 <= LUT_mem_MPORT_18_data[31:0]; // @[lut_35.scala 473:27]
    end
    if (reset) begin // @[lut_35.scala 236:31]
      read_stack19 <= 32'h0; // @[lut_35.scala 236:31]
    end else begin
      read_stack19 <= LUT_mem_MPORT_19_data[31:0]; // @[lut_35.scala 474:27]
    end
    if (reset) begin // @[lut_35.scala 237:31]
      read_stack20 <= 32'h0; // @[lut_35.scala 237:31]
    end else begin
      read_stack20 <= LUT_mem_MPORT_20_data[31:0]; // @[lut_35.scala 475:27]
    end
    if (reset) begin // @[lut_35.scala 238:31]
      read_stack21 <= 32'h0; // @[lut_35.scala 238:31]
    end else begin
      read_stack21 <= LUT_mem_MPORT_21_data[31:0]; // @[lut_35.scala 476:27]
    end
    if (reset) begin // @[lut_35.scala 239:31]
      read_stack22 <= 32'h0; // @[lut_35.scala 239:31]
    end else begin
      read_stack22 <= LUT_mem_MPORT_22_data[31:0]; // @[lut_35.scala 477:27]
    end
    if (reset) begin // @[lut_35.scala 240:31]
      read_stack23 <= 32'h0; // @[lut_35.scala 240:31]
    end else begin
      read_stack23 <= LUT_mem_MPORT_23_data[31:0]; // @[lut_35.scala 478:27]
    end
    if (reset) begin // @[lut_35.scala 241:31]
      read_stack24 <= 32'h0; // @[lut_35.scala 241:31]
    end else begin
      read_stack24 <= LUT_mem_MPORT_24_data[31:0]; // @[lut_35.scala 479:27]
    end
    if (reset) begin // @[lut_35.scala 242:31]
      read_stack25 <= 32'h0; // @[lut_35.scala 242:31]
    end else begin
      read_stack25 <= LUT_mem_MPORT_25_data[31:0]; // @[lut_35.scala 480:27]
    end
    if (reset) begin // @[lut_35.scala 243:31]
      read_stack26 <= 32'h0; // @[lut_35.scala 243:31]
    end else begin
      read_stack26 <= LUT_mem_MPORT_26_data[31:0]; // @[lut_35.scala 481:27]
    end
    if (reset) begin // @[lut_35.scala 244:31]
      read_stack27 <= 32'h0; // @[lut_35.scala 244:31]
    end else begin
      read_stack27 <= LUT_mem_MPORT_27_data[31:0]; // @[lut_35.scala 482:27]
    end
    if (reset) begin // @[lut_35.scala 245:31]
      read_stack28 <= 32'h0; // @[lut_35.scala 245:31]
    end else begin
      read_stack28 <= LUT_mem_MPORT_28_data[31:0]; // @[lut_35.scala 483:27]
    end
    if (reset) begin // @[lut_35.scala 246:31]
      read_stack29 <= 32'h0; // @[lut_35.scala 246:31]
    end else begin
      read_stack29 <= LUT_mem_MPORT_29_data[31:0]; // @[lut_35.scala 484:27]
    end
    if (reset) begin // @[lut_35.scala 247:31]
      read_stack30 <= 32'h0; // @[lut_35.scala 247:31]
    end else begin
      read_stack30 <= LUT_mem_MPORT_30_data[31:0]; // @[lut_35.scala 485:27]
    end
    if (reset) begin // @[lut_35.scala 248:31]
      read_stack31 <= 32'h0; // @[lut_35.scala 248:31]
    end else begin
      read_stack31 <= LUT_mem_MPORT_31_data[31:0]; // @[lut_35.scala 486:27]
    end
    if (reset) begin // @[lut_35.scala 249:31]
      read_stack32 <= 32'h0; // @[lut_35.scala 249:31]
    end else begin
      read_stack32 <= LUT_mem_MPORT_32_data[31:0]; // @[lut_35.scala 487:27]
    end
    if (reset) begin // @[lut_35.scala 250:31]
      read_stack33 <= 32'h0; // @[lut_35.scala 250:31]
    end else begin
      read_stack33 <= LUT_mem_MPORT_33_data[31:0]; // @[lut_35.scala 488:27]
    end
    if (reset) begin // @[lut_35.scala 251:31]
      read_stack34 <= 32'h0; // @[lut_35.scala 251:31]
    end else begin
      read_stack34 <= LUT_mem_MPORT_34_data[31:0]; // @[lut_35.scala 489:27]
    end
    if (reset) begin // @[lut_35.scala 253:31]
      push_0_1 <= 1'h0; // @[lut_35.scala 253:31]
    end else begin
      push_0_1 <= _GEN_9564;
    end
    if (reset) begin // @[lut_35.scala 254:31]
      push_1_1 <= 1'h0; // @[lut_35.scala 254:31]
    end else begin
      push_1_1 <= _GEN_9565;
    end
    if (reset) begin // @[lut_35.scala 255:31]
      push_2_1 <= 1'h0; // @[lut_35.scala 255:31]
    end else begin
      push_2_1 <= _GEN_9566;
    end
    if (reset) begin // @[lut_35.scala 256:31]
      push_3_1 <= 1'h0; // @[lut_35.scala 256:31]
    end else begin
      push_3_1 <= _GEN_9567;
    end
    if (reset) begin // @[lut_35.scala 257:31]
      push_4_1 <= 1'h0; // @[lut_35.scala 257:31]
    end else begin
      push_4_1 <= _GEN_9568;
    end
    if (reset) begin // @[lut_35.scala 258:31]
      push_5_1 <= 1'h0; // @[lut_35.scala 258:31]
    end else begin
      push_5_1 <= _GEN_9569;
    end
    if (reset) begin // @[lut_35.scala 259:31]
      push_6_1 <= 1'h0; // @[lut_35.scala 259:31]
    end else begin
      push_6_1 <= _GEN_9570;
    end
    if (reset) begin // @[lut_35.scala 260:31]
      push_7_1 <= 1'h0; // @[lut_35.scala 260:31]
    end else begin
      push_7_1 <= _GEN_9571;
    end
    if (reset) begin // @[lut_35.scala 261:31]
      push_8_1 <= 1'h0; // @[lut_35.scala 261:31]
    end else begin
      push_8_1 <= _GEN_9572;
    end
    if (reset) begin // @[lut_35.scala 262:31]
      push_9_1 <= 1'h0; // @[lut_35.scala 262:31]
    end else begin
      push_9_1 <= _GEN_9573;
    end
    if (reset) begin // @[lut_35.scala 263:32]
      push_10_1 <= 1'h0; // @[lut_35.scala 263:32]
    end else begin
      push_10_1 <= _GEN_9574;
    end
    if (reset) begin // @[lut_35.scala 264:32]
      push_11_1 <= 1'h0; // @[lut_35.scala 264:32]
    end else begin
      push_11_1 <= _GEN_9575;
    end
    if (reset) begin // @[lut_35.scala 265:32]
      push_12_1 <= 1'h0; // @[lut_35.scala 265:32]
    end else begin
      push_12_1 <= _GEN_9576;
    end
    if (reset) begin // @[lut_35.scala 266:32]
      push_13_1 <= 1'h0; // @[lut_35.scala 266:32]
    end else begin
      push_13_1 <= _GEN_9577;
    end
    if (reset) begin // @[lut_35.scala 267:32]
      push_14_1 <= 1'h0; // @[lut_35.scala 267:32]
    end else begin
      push_14_1 <= _GEN_9578;
    end
    if (reset) begin // @[lut_35.scala 268:32]
      push_15_1 <= 1'h0; // @[lut_35.scala 268:32]
    end else begin
      push_15_1 <= _GEN_9579;
    end
    if (reset) begin // @[lut_35.scala 269:32]
      push_16_1 <= 1'h0; // @[lut_35.scala 269:32]
    end else begin
      push_16_1 <= _GEN_9580;
    end
    if (reset) begin // @[lut_35.scala 270:32]
      push_17_1 <= 1'h0; // @[lut_35.scala 270:32]
    end else begin
      push_17_1 <= _GEN_9581;
    end
    if (reset) begin // @[lut_35.scala 271:32]
      push_18_1 <= 1'h0; // @[lut_35.scala 271:32]
    end else begin
      push_18_1 <= _GEN_9582;
    end
    if (reset) begin // @[lut_35.scala 272:32]
      push_19_1 <= 1'h0; // @[lut_35.scala 272:32]
    end else begin
      push_19_1 <= _GEN_9583;
    end
    if (reset) begin // @[lut_35.scala 273:32]
      push_20_1 <= 1'h0; // @[lut_35.scala 273:32]
    end else begin
      push_20_1 <= _GEN_9584;
    end
    if (reset) begin // @[lut_35.scala 274:32]
      push_21_1 <= 1'h0; // @[lut_35.scala 274:32]
    end else begin
      push_21_1 <= _GEN_9585;
    end
    if (reset) begin // @[lut_35.scala 275:32]
      push_22_1 <= 1'h0; // @[lut_35.scala 275:32]
    end else begin
      push_22_1 <= _GEN_9586;
    end
    if (reset) begin // @[lut_35.scala 276:32]
      push_23_1 <= 1'h0; // @[lut_35.scala 276:32]
    end else begin
      push_23_1 <= _GEN_9587;
    end
    if (reset) begin // @[lut_35.scala 277:32]
      push_24_1 <= 1'h0; // @[lut_35.scala 277:32]
    end else begin
      push_24_1 <= _GEN_9588;
    end
    if (reset) begin // @[lut_35.scala 278:32]
      push_25_1 <= 1'h0; // @[lut_35.scala 278:32]
    end else begin
      push_25_1 <= _GEN_9589;
    end
    if (reset) begin // @[lut_35.scala 279:32]
      push_26_1 <= 1'h0; // @[lut_35.scala 279:32]
    end else begin
      push_26_1 <= _GEN_9590;
    end
    if (reset) begin // @[lut_35.scala 280:32]
      push_27_1 <= 1'h0; // @[lut_35.scala 280:32]
    end else begin
      push_27_1 <= _GEN_9591;
    end
    if (reset) begin // @[lut_35.scala 281:32]
      push_28_1 <= 1'h0; // @[lut_35.scala 281:32]
    end else begin
      push_28_1 <= _GEN_9592;
    end
    if (reset) begin // @[lut_35.scala 282:32]
      push_29_1 <= 1'h0; // @[lut_35.scala 282:32]
    end else begin
      push_29_1 <= _GEN_9593;
    end
    if (reset) begin // @[lut_35.scala 283:32]
      push_30_1 <= 1'h0; // @[lut_35.scala 283:32]
    end else begin
      push_30_1 <= _GEN_9594;
    end
    if (reset) begin // @[lut_35.scala 284:32]
      push_31_1 <= 1'h0; // @[lut_35.scala 284:32]
    end else begin
      push_31_1 <= _GEN_9595;
    end
    if (reset) begin // @[lut_35.scala 285:32]
      push_32_1 <= 1'h0; // @[lut_35.scala 285:32]
    end else begin
      push_32_1 <= _GEN_9596;
    end
    if (reset) begin // @[lut_35.scala 286:32]
      push_33_1 <= 1'h0; // @[lut_35.scala 286:32]
    end else begin
      push_33_1 <= _GEN_9597;
    end
    if (reset) begin // @[lut_35.scala 287:32]
      push_34_1 <= 1'h0; // @[lut_35.scala 287:32]
    end else begin
      push_34_1 <= _GEN_9598;
    end
    if (reset) begin // @[lut_35.scala 291:40]
      push_1 <= 1'h0; // @[lut_35.scala 291:40]
    end else begin
      push_1 <= _T_36;
    end
    if (reset) begin // @[lut_35.scala 292:41]
      push_valid <= 1'h0; // @[lut_35.scala 292:41]
    end else begin
      push_valid <= _GEN_3;
    end
    if (reset) begin // @[lut_35.scala 294:41]
      push_ray_id <= 32'h0; // @[lut_35.scala 294:41]
    end else if (io_push & io_push_valid) begin // @[lut_35.scala 501:46]
      push_ray_id <= io_ray_id_push; // @[lut_35.scala 505:26]
    end
    if (reset) begin // @[lut_35.scala 334:41]
      push_valid_2 <= 1'h0; // @[lut_35.scala 334:41]
    end else begin
      push_valid_2 <= _GEN_9599;
    end
    if (reset) begin // @[lut_35.scala 340:33]
      dispatch_reg_0 <= 1'h0; // @[lut_35.scala 340:33]
    end else begin
      dispatch_reg_0 <= io_dispatch_0; // @[lut_35.scala 377:25]
    end
    if (reset) begin // @[lut_35.scala 341:33]
      dispatch_reg_1 <= 1'h0; // @[lut_35.scala 341:33]
    end else begin
      dispatch_reg_1 <= io_dispatch_1; // @[lut_35.scala 378:25]
    end
    if (reset) begin // @[lut_35.scala 342:33]
      dispatch_reg_2 <= 1'h0; // @[lut_35.scala 342:33]
    end else begin
      dispatch_reg_2 <= io_dispatch_2; // @[lut_35.scala 379:25]
    end
    if (reset) begin // @[lut_35.scala 343:33]
      dispatch_reg_3 <= 1'h0; // @[lut_35.scala 343:33]
    end else begin
      dispatch_reg_3 <= io_dispatch_3; // @[lut_35.scala 380:25]
    end
    if (reset) begin // @[lut_35.scala 344:33]
      dispatch_reg_4 <= 1'h0; // @[lut_35.scala 344:33]
    end else begin
      dispatch_reg_4 <= io_dispatch_4; // @[lut_35.scala 381:25]
    end
    if (reset) begin // @[lut_35.scala 345:33]
      dispatch_reg_5 <= 1'h0; // @[lut_35.scala 345:33]
    end else begin
      dispatch_reg_5 <= io_dispatch_5; // @[lut_35.scala 382:25]
    end
    if (reset) begin // @[lut_35.scala 346:33]
      dispatch_reg_6 <= 1'h0; // @[lut_35.scala 346:33]
    end else begin
      dispatch_reg_6 <= io_dispatch_6; // @[lut_35.scala 383:25]
    end
    if (reset) begin // @[lut_35.scala 347:33]
      dispatch_reg_7 <= 1'h0; // @[lut_35.scala 347:33]
    end else begin
      dispatch_reg_7 <= io_dispatch_7; // @[lut_35.scala 384:25]
    end
    if (reset) begin // @[lut_35.scala 348:33]
      dispatch_reg_8 <= 1'h0; // @[lut_35.scala 348:33]
    end else begin
      dispatch_reg_8 <= io_dispatch_8; // @[lut_35.scala 385:25]
    end
    if (reset) begin // @[lut_35.scala 349:33]
      dispatch_reg_9 <= 1'h0; // @[lut_35.scala 349:33]
    end else begin
      dispatch_reg_9 <= io_dispatch_9; // @[lut_35.scala 386:25]
    end
    if (reset) begin // @[lut_35.scala 350:34]
      dispatch_reg_10 <= 1'h0; // @[lut_35.scala 350:34]
    end else begin
      dispatch_reg_10 <= io_dispatch_10; // @[lut_35.scala 387:26]
    end
    if (reset) begin // @[lut_35.scala 351:34]
      dispatch_reg_11 <= 1'h0; // @[lut_35.scala 351:34]
    end else begin
      dispatch_reg_11 <= io_dispatch_11; // @[lut_35.scala 388:26]
    end
    if (reset) begin // @[lut_35.scala 352:34]
      dispatch_reg_12 <= 1'h0; // @[lut_35.scala 352:34]
    end else begin
      dispatch_reg_12 <= io_dispatch_12; // @[lut_35.scala 389:26]
    end
    if (reset) begin // @[lut_35.scala 353:34]
      dispatch_reg_13 <= 1'h0; // @[lut_35.scala 353:34]
    end else begin
      dispatch_reg_13 <= io_dispatch_13; // @[lut_35.scala 390:26]
    end
    if (reset) begin // @[lut_35.scala 354:34]
      dispatch_reg_14 <= 1'h0; // @[lut_35.scala 354:34]
    end else begin
      dispatch_reg_14 <= io_dispatch_14; // @[lut_35.scala 391:26]
    end
    if (reset) begin // @[lut_35.scala 355:34]
      dispatch_reg_15 <= 1'h0; // @[lut_35.scala 355:34]
    end else begin
      dispatch_reg_15 <= io_dispatch_15; // @[lut_35.scala 392:26]
    end
    if (reset) begin // @[lut_35.scala 356:34]
      dispatch_reg_16 <= 1'h0; // @[lut_35.scala 356:34]
    end else begin
      dispatch_reg_16 <= io_dispatch_16; // @[lut_35.scala 393:26]
    end
    if (reset) begin // @[lut_35.scala 357:34]
      dispatch_reg_17 <= 1'h0; // @[lut_35.scala 357:34]
    end else begin
      dispatch_reg_17 <= io_dispatch_17; // @[lut_35.scala 394:26]
    end
    if (reset) begin // @[lut_35.scala 358:34]
      dispatch_reg_18 <= 1'h0; // @[lut_35.scala 358:34]
    end else begin
      dispatch_reg_18 <= io_dispatch_18; // @[lut_35.scala 395:26]
    end
    if (reset) begin // @[lut_35.scala 359:34]
      dispatch_reg_19 <= 1'h0; // @[lut_35.scala 359:34]
    end else begin
      dispatch_reg_19 <= io_dispatch_19; // @[lut_35.scala 396:26]
    end
    if (reset) begin // @[lut_35.scala 360:34]
      dispatch_reg_20 <= 1'h0; // @[lut_35.scala 360:34]
    end else begin
      dispatch_reg_20 <= io_dispatch_20; // @[lut_35.scala 397:26]
    end
    if (reset) begin // @[lut_35.scala 361:34]
      dispatch_reg_21 <= 1'h0; // @[lut_35.scala 361:34]
    end else begin
      dispatch_reg_21 <= io_dispatch_21; // @[lut_35.scala 398:26]
    end
    if (reset) begin // @[lut_35.scala 362:34]
      dispatch_reg_22 <= 1'h0; // @[lut_35.scala 362:34]
    end else begin
      dispatch_reg_22 <= io_dispatch_22; // @[lut_35.scala 399:26]
    end
    if (reset) begin // @[lut_35.scala 363:34]
      dispatch_reg_23 <= 1'h0; // @[lut_35.scala 363:34]
    end else begin
      dispatch_reg_23 <= io_dispatch_23; // @[lut_35.scala 400:26]
    end
    if (reset) begin // @[lut_35.scala 364:34]
      dispatch_reg_24 <= 1'h0; // @[lut_35.scala 364:34]
    end else begin
      dispatch_reg_24 <= io_dispatch_24; // @[lut_35.scala 401:26]
    end
    if (reset) begin // @[lut_35.scala 365:34]
      dispatch_reg_25 <= 1'h0; // @[lut_35.scala 365:34]
    end else begin
      dispatch_reg_25 <= io_dispatch_25; // @[lut_35.scala 402:26]
    end
    if (reset) begin // @[lut_35.scala 366:34]
      dispatch_reg_26 <= 1'h0; // @[lut_35.scala 366:34]
    end else begin
      dispatch_reg_26 <= io_dispatch_26; // @[lut_35.scala 403:26]
    end
    if (reset) begin // @[lut_35.scala 367:34]
      dispatch_reg_27 <= 1'h0; // @[lut_35.scala 367:34]
    end else begin
      dispatch_reg_27 <= io_dispatch_27; // @[lut_35.scala 404:26]
    end
    if (reset) begin // @[lut_35.scala 368:34]
      dispatch_reg_28 <= 1'h0; // @[lut_35.scala 368:34]
    end else begin
      dispatch_reg_28 <= io_dispatch_28; // @[lut_35.scala 405:26]
    end
    if (reset) begin // @[lut_35.scala 369:34]
      dispatch_reg_29 <= 1'h0; // @[lut_35.scala 369:34]
    end else begin
      dispatch_reg_29 <= io_dispatch_29; // @[lut_35.scala 406:26]
    end
    if (reset) begin // @[lut_35.scala 370:34]
      dispatch_reg_30 <= 1'h0; // @[lut_35.scala 370:34]
    end else begin
      dispatch_reg_30 <= io_dispatch_30; // @[lut_35.scala 407:26]
    end
    if (reset) begin // @[lut_35.scala 371:34]
      dispatch_reg_31 <= 1'h0; // @[lut_35.scala 371:34]
    end else begin
      dispatch_reg_31 <= io_dispatch_31; // @[lut_35.scala 408:26]
    end
    if (reset) begin // @[lut_35.scala 372:34]
      dispatch_reg_32 <= 1'h0; // @[lut_35.scala 372:34]
    end else begin
      dispatch_reg_32 <= io_dispatch_32; // @[lut_35.scala 409:26]
    end
    if (reset) begin // @[lut_35.scala 373:34]
      dispatch_reg_33 <= 1'h0; // @[lut_35.scala 373:34]
    end else begin
      dispatch_reg_33 <= io_dispatch_33; // @[lut_35.scala 410:26]
    end
    if (reset) begin // @[lut_35.scala 374:34]
      dispatch_reg_34 <= 1'h0; // @[lut_35.scala 374:34]
    end else begin
      dispatch_reg_34 <= io_dispatch_34; // @[lut_35.scala 411:26]
    end
    if (reset) begin // @[lut_35.scala 521:39]
      push_mem_temp <= 6'h23; // @[lut_35.scala 521:39]
    end else if (push_1 & push_valid) begin // @[lut_35.scala 524:46]
      if (!(LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid)) begin // @[lut_35.scala 525:68]
        if (!(LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid)) begin // @[lut_35.scala 563:74]
          push_mem_temp <= _GEN_8968;
        end
      end
    end else begin
      push_mem_temp <= 6'h23; // @[lut_35.scala 3413:42]
    end
    if (reset) begin // @[lut_35.scala 522:39]
      push_id_temp <= 32'h0; // @[lut_35.scala 522:39]
    end else if (push_1 & push_valid) begin // @[lut_35.scala 524:46]
      if (!(LUT_mem_MPORT_35_data[31:0] == push_ray_id & push_valid)) begin // @[lut_35.scala 525:68]
        if (!(LUT_mem_MPORT_36_data[31:0] == push_ray_id & push_valid)) begin // @[lut_35.scala 563:74]
          push_id_temp <= _GEN_8969;
        end
      end
    end else begin
      push_id_temp <= 32'h0; // @[lut_35.scala 3414:42]
    end
    if (reset) begin // @[lut_35.scala 3494:50]
      pop_1 <= 1'h0; // @[lut_35.scala 3494:50]
    end else begin
      pop_1 <= _T_567;
    end
    if (reset) begin // @[lut_35.scala 3495:38]
      read_stack0_pop <= 32'h0; // @[lut_35.scala 3495:38]
    end else begin
      read_stack0_pop <= LUT_mem_MPORT_105_data[31:0]; // @[lut_35.scala 3580:30]
    end
    if (reset) begin // @[lut_35.scala 3496:38]
      read_stack1_pop <= 32'h0; // @[lut_35.scala 3496:38]
    end else begin
      read_stack1_pop <= LUT_mem_MPORT_106_data[31:0]; // @[lut_35.scala 3581:30]
    end
    if (reset) begin // @[lut_35.scala 3497:38]
      read_stack2_pop <= 32'h0; // @[lut_35.scala 3497:38]
    end else begin
      read_stack2_pop <= LUT_mem_MPORT_107_data[31:0]; // @[lut_35.scala 3582:30]
    end
    if (reset) begin // @[lut_35.scala 3498:38]
      read_stack3_pop <= 32'h0; // @[lut_35.scala 3498:38]
    end else begin
      read_stack3_pop <= LUT_mem_MPORT_108_data[31:0]; // @[lut_35.scala 3583:30]
    end
    if (reset) begin // @[lut_35.scala 3499:38]
      read_stack4_pop <= 32'h0; // @[lut_35.scala 3499:38]
    end else begin
      read_stack4_pop <= LUT_mem_MPORT_109_data[31:0]; // @[lut_35.scala 3584:30]
    end
    if (reset) begin // @[lut_35.scala 3500:38]
      read_stack5_pop <= 32'h0; // @[lut_35.scala 3500:38]
    end else begin
      read_stack5_pop <= LUT_mem_MPORT_110_data[31:0]; // @[lut_35.scala 3585:30]
    end
    if (reset) begin // @[lut_35.scala 3501:38]
      read_stack6_pop <= 32'h0; // @[lut_35.scala 3501:38]
    end else begin
      read_stack6_pop <= LUT_mem_MPORT_111_data[31:0]; // @[lut_35.scala 3586:30]
    end
    if (reset) begin // @[lut_35.scala 3502:38]
      read_stack7_pop <= 32'h0; // @[lut_35.scala 3502:38]
    end else begin
      read_stack7_pop <= LUT_mem_MPORT_112_data[31:0]; // @[lut_35.scala 3587:30]
    end
    if (reset) begin // @[lut_35.scala 3503:38]
      read_stack8_pop <= 32'h0; // @[lut_35.scala 3503:38]
    end else begin
      read_stack8_pop <= LUT_mem_MPORT_113_data[31:0]; // @[lut_35.scala 3588:30]
    end
    if (reset) begin // @[lut_35.scala 3504:38]
      read_stack9_pop <= 32'h0; // @[lut_35.scala 3504:38]
    end else begin
      read_stack9_pop <= LUT_mem_MPORT_114_data[31:0]; // @[lut_35.scala 3589:30]
    end
    if (reset) begin // @[lut_35.scala 3505:39]
      read_stack10_pop <= 32'h0; // @[lut_35.scala 3505:39]
    end else begin
      read_stack10_pop <= LUT_mem_MPORT_115_data[31:0]; // @[lut_35.scala 3591:31]
    end
    if (reset) begin // @[lut_35.scala 3506:39]
      read_stack11_pop <= 32'h0; // @[lut_35.scala 3506:39]
    end else begin
      read_stack11_pop <= LUT_mem_MPORT_116_data[31:0]; // @[lut_35.scala 3592:31]
    end
    if (reset) begin // @[lut_35.scala 3507:39]
      read_stack12_pop <= 32'h0; // @[lut_35.scala 3507:39]
    end else begin
      read_stack12_pop <= LUT_mem_MPORT_117_data[31:0]; // @[lut_35.scala 3593:31]
    end
    if (reset) begin // @[lut_35.scala 3508:39]
      read_stack13_pop <= 32'h0; // @[lut_35.scala 3508:39]
    end else begin
      read_stack13_pop <= LUT_mem_MPORT_118_data[31:0]; // @[lut_35.scala 3594:31]
    end
    if (reset) begin // @[lut_35.scala 3509:39]
      read_stack14_pop <= 32'h0; // @[lut_35.scala 3509:39]
    end else begin
      read_stack14_pop <= LUT_mem_MPORT_119_data[31:0]; // @[lut_35.scala 3595:31]
    end
    if (reset) begin // @[lut_35.scala 3510:39]
      read_stack15_pop <= 32'h0; // @[lut_35.scala 3510:39]
    end else begin
      read_stack15_pop <= LUT_mem_MPORT_120_data[31:0]; // @[lut_35.scala 3596:31]
    end
    if (reset) begin // @[lut_35.scala 3511:39]
      read_stack16_pop <= 32'h0; // @[lut_35.scala 3511:39]
    end else begin
      read_stack16_pop <= LUT_mem_MPORT_121_data[31:0]; // @[lut_35.scala 3597:31]
    end
    if (reset) begin // @[lut_35.scala 3512:39]
      read_stack17_pop <= 32'h0; // @[lut_35.scala 3512:39]
    end else begin
      read_stack17_pop <= LUT_mem_MPORT_122_data[31:0]; // @[lut_35.scala 3598:31]
    end
    if (reset) begin // @[lut_35.scala 3513:39]
      read_stack18_pop <= 32'h0; // @[lut_35.scala 3513:39]
    end else begin
      read_stack18_pop <= LUT_mem_MPORT_123_data[31:0]; // @[lut_35.scala 3599:31]
    end
    if (reset) begin // @[lut_35.scala 3514:39]
      read_stack19_pop <= 32'h0; // @[lut_35.scala 3514:39]
    end else begin
      read_stack19_pop <= LUT_mem_MPORT_124_data[31:0]; // @[lut_35.scala 3600:31]
    end
    if (reset) begin // @[lut_35.scala 3515:39]
      read_stack20_pop <= 32'h0; // @[lut_35.scala 3515:39]
    end else begin
      read_stack20_pop <= LUT_mem_MPORT_125_data[31:0]; // @[lut_35.scala 3602:31]
    end
    if (reset) begin // @[lut_35.scala 3516:39]
      read_stack21_pop <= 32'h0; // @[lut_35.scala 3516:39]
    end else begin
      read_stack21_pop <= LUT_mem_MPORT_126_data[31:0]; // @[lut_35.scala 3603:31]
    end
    if (reset) begin // @[lut_35.scala 3517:39]
      read_stack22_pop <= 32'h0; // @[lut_35.scala 3517:39]
    end else begin
      read_stack22_pop <= LUT_mem_MPORT_127_data[31:0]; // @[lut_35.scala 3604:31]
    end
    if (reset) begin // @[lut_35.scala 3518:39]
      read_stack23_pop <= 32'h0; // @[lut_35.scala 3518:39]
    end else begin
      read_stack23_pop <= LUT_mem_MPORT_128_data[31:0]; // @[lut_35.scala 3605:31]
    end
    if (reset) begin // @[lut_35.scala 3519:39]
      read_stack24_pop <= 32'h0; // @[lut_35.scala 3519:39]
    end else begin
      read_stack24_pop <= LUT_mem_MPORT_129_data[31:0]; // @[lut_35.scala 3606:31]
    end
    if (reset) begin // @[lut_35.scala 3520:39]
      read_stack25_pop <= 32'h0; // @[lut_35.scala 3520:39]
    end else begin
      read_stack25_pop <= LUT_mem_MPORT_130_data[31:0]; // @[lut_35.scala 3607:31]
    end
    if (reset) begin // @[lut_35.scala 3521:39]
      read_stack26_pop <= 32'h0; // @[lut_35.scala 3521:39]
    end else begin
      read_stack26_pop <= LUT_mem_MPORT_131_data[31:0]; // @[lut_35.scala 3608:31]
    end
    if (reset) begin // @[lut_35.scala 3522:39]
      read_stack27_pop <= 32'h0; // @[lut_35.scala 3522:39]
    end else begin
      read_stack27_pop <= LUT_mem_MPORT_132_data[31:0]; // @[lut_35.scala 3609:31]
    end
    if (reset) begin // @[lut_35.scala 3523:39]
      read_stack28_pop <= 32'h0; // @[lut_35.scala 3523:39]
    end else begin
      read_stack28_pop <= LUT_mem_MPORT_133_data[31:0]; // @[lut_35.scala 3610:31]
    end
    if (reset) begin // @[lut_35.scala 3524:39]
      read_stack29_pop <= 32'h0; // @[lut_35.scala 3524:39]
    end else begin
      read_stack29_pop <= LUT_mem_MPORT_134_data[31:0]; // @[lut_35.scala 3611:31]
    end
    if (reset) begin // @[lut_35.scala 3525:39]
      read_stack30_pop <= 32'h0; // @[lut_35.scala 3525:39]
    end else begin
      read_stack30_pop <= LUT_mem_MPORT_135_data[31:0]; // @[lut_35.scala 3613:31]
    end
    if (reset) begin // @[lut_35.scala 3526:39]
      read_stack31_pop <= 32'h0; // @[lut_35.scala 3526:39]
    end else begin
      read_stack31_pop <= LUT_mem_MPORT_136_data[31:0]; // @[lut_35.scala 3614:31]
    end
    if (reset) begin // @[lut_35.scala 3527:39]
      read_stack32_pop <= 32'h0; // @[lut_35.scala 3527:39]
    end else begin
      read_stack32_pop <= LUT_mem_MPORT_137_data[31:0]; // @[lut_35.scala 3615:31]
    end
    if (reset) begin // @[lut_35.scala 3528:39]
      read_stack33_pop <= 32'h0; // @[lut_35.scala 3528:39]
    end else begin
      read_stack33_pop <= LUT_mem_MPORT_138_data[31:0]; // @[lut_35.scala 3616:31]
    end
    if (reset) begin // @[lut_35.scala 3529:39]
      read_stack34_pop <= 32'h0; // @[lut_35.scala 3529:39]
    end else begin
      read_stack34_pop <= LUT_mem_MPORT_139_data[31:0]; // @[lut_35.scala 3617:31]
    end
    if (reset) begin // @[lut_35.scala 3532:37]
      pop_ray_id <= 32'h0; // @[lut_35.scala 3532:37]
    end else if (io_pop & io_pop_valid) begin // @[lut_35.scala 3619:44]
      pop_ray_id <= io_ray_id_pop; // @[lut_35.scala 3624:26]
    end
    if (reset) begin // @[lut_35.scala 3533:37]
      pop_hitT_1 <= 32'h0; // @[lut_35.scala 3533:37]
    end else if (io_pop & io_pop_valid) begin // @[lut_35.scala 3619:44]
      pop_hitT_1 <= io_hitT_in; // @[lut_35.scala 3625:26]
    end
    if (reset) begin // @[lut_35.scala 3534:36]
      pop_valid <= 1'h0; // @[lut_35.scala 3534:36]
    end else begin
      pop_valid <= _T_567;
    end
    if (reset) begin // @[lut_35.scala 3537:46]
      pop_0_1 <= 1'h0; // @[lut_35.scala 3537:46]
    end else begin
      pop_0_1 <= _GEN_10618;
    end
    if (reset) begin // @[lut_35.scala 3538:46]
      pop_1_1 <= 1'h0; // @[lut_35.scala 3538:46]
    end else begin
      pop_1_1 <= _GEN_10619;
    end
    if (reset) begin // @[lut_35.scala 3539:46]
      pop_2_1 <= 1'h0; // @[lut_35.scala 3539:46]
    end else begin
      pop_2_1 <= _GEN_10620;
    end
    if (reset) begin // @[lut_35.scala 3540:46]
      pop_3_1 <= 1'h0; // @[lut_35.scala 3540:46]
    end else begin
      pop_3_1 <= _GEN_10621;
    end
    if (reset) begin // @[lut_35.scala 3541:46]
      pop_4_1 <= 1'h0; // @[lut_35.scala 3541:46]
    end else begin
      pop_4_1 <= _GEN_10622;
    end
    if (reset) begin // @[lut_35.scala 3542:46]
      pop_5_1 <= 1'h0; // @[lut_35.scala 3542:46]
    end else begin
      pop_5_1 <= _GEN_10623;
    end
    if (reset) begin // @[lut_35.scala 3543:46]
      pop_6_1 <= 1'h0; // @[lut_35.scala 3543:46]
    end else begin
      pop_6_1 <= _GEN_10624;
    end
    if (reset) begin // @[lut_35.scala 3544:46]
      pop_7_1 <= 1'h0; // @[lut_35.scala 3544:46]
    end else begin
      pop_7_1 <= _GEN_10625;
    end
    if (reset) begin // @[lut_35.scala 3545:46]
      pop_8_1 <= 1'h0; // @[lut_35.scala 3545:46]
    end else begin
      pop_8_1 <= _GEN_10626;
    end
    if (reset) begin // @[lut_35.scala 3546:46]
      pop_9_1 <= 1'h0; // @[lut_35.scala 3546:46]
    end else begin
      pop_9_1 <= _GEN_10627;
    end
    if (reset) begin // @[lut_35.scala 3547:47]
      pop_10_1 <= 1'h0; // @[lut_35.scala 3547:47]
    end else begin
      pop_10_1 <= _GEN_10628;
    end
    if (reset) begin // @[lut_35.scala 3548:47]
      pop_11_1 <= 1'h0; // @[lut_35.scala 3548:47]
    end else begin
      pop_11_1 <= _GEN_10629;
    end
    if (reset) begin // @[lut_35.scala 3549:47]
      pop_12_1 <= 1'h0; // @[lut_35.scala 3549:47]
    end else begin
      pop_12_1 <= _GEN_10630;
    end
    if (reset) begin // @[lut_35.scala 3550:47]
      pop_13_1 <= 1'h0; // @[lut_35.scala 3550:47]
    end else begin
      pop_13_1 <= _GEN_10631;
    end
    if (reset) begin // @[lut_35.scala 3551:47]
      pop_14_1 <= 1'h0; // @[lut_35.scala 3551:47]
    end else begin
      pop_14_1 <= _GEN_10632;
    end
    if (reset) begin // @[lut_35.scala 3552:47]
      pop_15_1 <= 1'h0; // @[lut_35.scala 3552:47]
    end else begin
      pop_15_1 <= _GEN_10633;
    end
    if (reset) begin // @[lut_35.scala 3553:47]
      pop_16_1 <= 1'h0; // @[lut_35.scala 3553:47]
    end else begin
      pop_16_1 <= _GEN_10634;
    end
    if (reset) begin // @[lut_35.scala 3554:47]
      pop_17_1 <= 1'h0; // @[lut_35.scala 3554:47]
    end else begin
      pop_17_1 <= _GEN_10635;
    end
    if (reset) begin // @[lut_35.scala 3555:47]
      pop_18_1 <= 1'h0; // @[lut_35.scala 3555:47]
    end else begin
      pop_18_1 <= _GEN_10636;
    end
    if (reset) begin // @[lut_35.scala 3556:47]
      pop_19_1 <= 1'h0; // @[lut_35.scala 3556:47]
    end else begin
      pop_19_1 <= _GEN_10637;
    end
    if (reset) begin // @[lut_35.scala 3557:47]
      pop_20_1 <= 1'h0; // @[lut_35.scala 3557:47]
    end else begin
      pop_20_1 <= _GEN_10638;
    end
    if (reset) begin // @[lut_35.scala 3558:47]
      pop_21_1 <= 1'h0; // @[lut_35.scala 3558:47]
    end else begin
      pop_21_1 <= _GEN_10639;
    end
    if (reset) begin // @[lut_35.scala 3559:47]
      pop_22_1 <= 1'h0; // @[lut_35.scala 3559:47]
    end else begin
      pop_22_1 <= _GEN_10640;
    end
    if (reset) begin // @[lut_35.scala 3560:47]
      pop_23_1 <= 1'h0; // @[lut_35.scala 3560:47]
    end else begin
      pop_23_1 <= _GEN_10641;
    end
    if (reset) begin // @[lut_35.scala 3561:47]
      pop_24_1 <= 1'h0; // @[lut_35.scala 3561:47]
    end else begin
      pop_24_1 <= _GEN_10642;
    end
    if (reset) begin // @[lut_35.scala 3562:47]
      pop_25_1 <= 1'h0; // @[lut_35.scala 3562:47]
    end else begin
      pop_25_1 <= _GEN_10643;
    end
    if (reset) begin // @[lut_35.scala 3563:47]
      pop_26_1 <= 1'h0; // @[lut_35.scala 3563:47]
    end else begin
      pop_26_1 <= _GEN_10644;
    end
    if (reset) begin // @[lut_35.scala 3564:47]
      pop_27_1 <= 1'h0; // @[lut_35.scala 3564:47]
    end else begin
      pop_27_1 <= _GEN_10645;
    end
    if (reset) begin // @[lut_35.scala 3565:47]
      pop_28_1 <= 1'h0; // @[lut_35.scala 3565:47]
    end else begin
      pop_28_1 <= _GEN_10646;
    end
    if (reset) begin // @[lut_35.scala 3566:47]
      pop_29_1 <= 1'h0; // @[lut_35.scala 3566:47]
    end else begin
      pop_29_1 <= _GEN_10647;
    end
    if (reset) begin // @[lut_35.scala 3567:47]
      pop_30_1 <= 1'h0; // @[lut_35.scala 3567:47]
    end else begin
      pop_30_1 <= _GEN_10648;
    end
    if (reset) begin // @[lut_35.scala 3568:47]
      pop_31_1 <= 1'h0; // @[lut_35.scala 3568:47]
    end else begin
      pop_31_1 <= _GEN_10649;
    end
    if (reset) begin // @[lut_35.scala 3569:47]
      pop_32_1 <= 1'h0; // @[lut_35.scala 3569:47]
    end else begin
      pop_32_1 <= _GEN_10650;
    end
    if (reset) begin // @[lut_35.scala 3570:47]
      pop_33_1 <= 1'h0; // @[lut_35.scala 3570:47]
    end else begin
      pop_33_1 <= _GEN_10651;
    end
    if (reset) begin // @[lut_35.scala 3571:47]
      pop_34_1 <= 1'h0; // @[lut_35.scala 3571:47]
    end else begin
      pop_34_1 <= _GEN_10652;
    end
    if (reset) begin // @[lut_35.scala 3573:47]
      pop_valid_2 <= 1'h0; // @[lut_35.scala 3573:47]
    end else begin
      pop_valid_2 <= _GEN_10653;
    end
    if (reset) begin // @[lut_35.scala 3575:47]
      pop_ray_id_2 <= 32'h0; // @[lut_35.scala 3575:47]
    end else if (pop_1 & pop_valid) begin // @[lut_35.scala 3649:46]
      if (read_stack0_pop == pop_ray_id & pop_valid) begin // @[lut_35.scala 3650:67]
        pop_ray_id_2 <= pop_ray_id; // @[lut_35.scala 3688:34]
      end else if (read_stack1_pop == pop_ray_id & pop_valid) begin // @[lut_35.scala 3690:77]
        pop_ray_id_2 <= pop_ray_id; // @[lut_35.scala 3728:38]
      end else begin
        pop_ray_id_2 <= _GEN_10538;
      end
    end
    if (reset) begin // @[lut_35.scala 3576:47]
      pop_hitT_2 <= 32'h0; // @[lut_35.scala 3576:47]
    end else if (pop_1 & pop_valid) begin // @[lut_35.scala 3649:46]
      if (read_stack0_pop == pop_ray_id & pop_valid) begin // @[lut_35.scala 3650:67]
        pop_hitT_2 <= pop_hitT_1; // @[lut_35.scala 3689:37]
      end else if (read_stack1_pop == pop_ray_id & pop_valid) begin // @[lut_35.scala 3690:77]
        pop_hitT_2 <= pop_hitT_1; // @[lut_35.scala 3729:41]
      end else begin
        pop_hitT_2 <= _GEN_10539;
      end
    end
    if (reset) begin // @[lut_35.scala 3578:47]
      no_match <= 1'h0; // @[lut_35.scala 3578:47]
    end else begin
      no_match <= _T_640;
    end
    if (reset) begin // @[lut_35.scala 3644:51]
      no_match_1 <= 1'h0; // @[lut_35.scala 3644:51]
    end else begin
      no_match_1 <= no_match; // @[lut_35.scala 3646:41]
    end
    if (reset) begin // @[lut_35.scala 3645:51]
      no_match_2 <= 1'h0; // @[lut_35.scala 3645:51]
    end else begin
      no_match_2 <= no_match_1; // @[lut_35.scala 3647:41]
    end
    if (reset) begin // @[lut_35.scala 5175:38]
      clear_1 <= 1'h0; // @[lut_35.scala 5175:38]
    end else begin
      clear_1 <= io_clear;
    end
    if (reset) begin // @[lut_35.scala 5176:40]
      read_stack0_clear <= 32'h0; // @[lut_35.scala 5176:40]
    end else begin
      read_stack0_clear <= LUT_mem_MPORT_140_data[31:0]; // @[lut_35.scala 5255:32]
    end
    if (reset) begin // @[lut_35.scala 5177:40]
      read_stack1_clear <= 32'h0; // @[lut_35.scala 5177:40]
    end else begin
      read_stack1_clear <= LUT_mem_MPORT_141_data[31:0]; // @[lut_35.scala 5256:32]
    end
    if (reset) begin // @[lut_35.scala 5179:40]
      read_stack3_clear <= 32'h0; // @[lut_35.scala 5179:40]
    end else begin
      read_stack3_clear <= LUT_mem_MPORT_143_data[31:0]; // @[lut_35.scala 5258:32]
    end
    if (reset) begin // @[lut_35.scala 5180:40]
      read_stack4_clear <= 32'h0; // @[lut_35.scala 5180:40]
    end else begin
      read_stack4_clear <= LUT_mem_MPORT_144_data[31:0]; // @[lut_35.scala 5259:32]
    end
    if (reset) begin // @[lut_35.scala 5181:40]
      read_stack5_clear <= 32'h0; // @[lut_35.scala 5181:40]
    end else begin
      read_stack5_clear <= LUT_mem_MPORT_145_data[31:0]; // @[lut_35.scala 5260:32]
    end
    if (reset) begin // @[lut_35.scala 5182:40]
      read_stack6_clear <= 32'h0; // @[lut_35.scala 5182:40]
    end else begin
      read_stack6_clear <= LUT_mem_MPORT_146_data[31:0]; // @[lut_35.scala 5261:32]
    end
    if (reset) begin // @[lut_35.scala 5183:40]
      read_stack7_clear <= 32'h0; // @[lut_35.scala 5183:40]
    end else begin
      read_stack7_clear <= LUT_mem_MPORT_147_data[31:0]; // @[lut_35.scala 5262:32]
    end
    if (reset) begin // @[lut_35.scala 5184:40]
      read_stack8_clear <= 32'h0; // @[lut_35.scala 5184:40]
    end else begin
      read_stack8_clear <= LUT_mem_MPORT_148_data[31:0]; // @[lut_35.scala 5263:32]
    end
    if (reset) begin // @[lut_35.scala 5185:40]
      read_stack9_clear <= 32'h0; // @[lut_35.scala 5185:40]
    end else begin
      read_stack9_clear <= LUT_mem_MPORT_149_data[31:0]; // @[lut_35.scala 5264:32]
    end
    if (reset) begin // @[lut_35.scala 5186:41]
      read_stack10_clear <= 32'h0; // @[lut_35.scala 5186:41]
    end else begin
      read_stack10_clear <= LUT_mem_MPORT_150_data[31:0]; // @[lut_35.scala 5266:33]
    end
    if (reset) begin // @[lut_35.scala 5187:41]
      read_stack11_clear <= 32'h0; // @[lut_35.scala 5187:41]
    end else begin
      read_stack11_clear <= LUT_mem_MPORT_151_data[31:0]; // @[lut_35.scala 5267:33]
    end
    if (reset) begin // @[lut_35.scala 5188:41]
      read_stack12_clear <= 32'h0; // @[lut_35.scala 5188:41]
    end else begin
      read_stack12_clear <= LUT_mem_MPORT_152_data[31:0]; // @[lut_35.scala 5268:33]
    end
    if (reset) begin // @[lut_35.scala 5189:41]
      read_stack13_clear <= 32'h0; // @[lut_35.scala 5189:41]
    end else begin
      read_stack13_clear <= LUT_mem_MPORT_153_data[31:0]; // @[lut_35.scala 5269:33]
    end
    if (reset) begin // @[lut_35.scala 5190:41]
      read_stack14_clear <= 32'h0; // @[lut_35.scala 5190:41]
    end else begin
      read_stack14_clear <= LUT_mem_MPORT_154_data[31:0]; // @[lut_35.scala 5270:33]
    end
    if (reset) begin // @[lut_35.scala 5191:41]
      read_stack15_clear <= 32'h0; // @[lut_35.scala 5191:41]
    end else begin
      read_stack15_clear <= LUT_mem_MPORT_155_data[31:0]; // @[lut_35.scala 5271:33]
    end
    if (reset) begin // @[lut_35.scala 5192:41]
      read_stack16_clear <= 32'h0; // @[lut_35.scala 5192:41]
    end else begin
      read_stack16_clear <= LUT_mem_MPORT_156_data[31:0]; // @[lut_35.scala 5272:33]
    end
    if (reset) begin // @[lut_35.scala 5193:41]
      read_stack17_clear <= 32'h0; // @[lut_35.scala 5193:41]
    end else begin
      read_stack17_clear <= LUT_mem_MPORT_157_data[31:0]; // @[lut_35.scala 5273:33]
    end
    if (reset) begin // @[lut_35.scala 5194:41]
      read_stack18_clear <= 32'h0; // @[lut_35.scala 5194:41]
    end else begin
      read_stack18_clear <= LUT_mem_MPORT_158_data[31:0]; // @[lut_35.scala 5274:33]
    end
    if (reset) begin // @[lut_35.scala 5195:41]
      read_stack19_clear <= 32'h0; // @[lut_35.scala 5195:41]
    end else begin
      read_stack19_clear <= LUT_mem_MPORT_159_data[31:0]; // @[lut_35.scala 5275:33]
    end
    if (reset) begin // @[lut_35.scala 5196:41]
      read_stack20_clear <= 32'h0; // @[lut_35.scala 5196:41]
    end else begin
      read_stack20_clear <= LUT_mem_MPORT_160_data[31:0]; // @[lut_35.scala 5277:33]
    end
    if (reset) begin // @[lut_35.scala 5197:41]
      read_stack21_clear <= 32'h0; // @[lut_35.scala 5197:41]
    end else begin
      read_stack21_clear <= LUT_mem_MPORT_161_data[31:0]; // @[lut_35.scala 5278:33]
    end
    if (reset) begin // @[lut_35.scala 5198:41]
      read_stack22_clear <= 32'h0; // @[lut_35.scala 5198:41]
    end else begin
      read_stack22_clear <= LUT_mem_MPORT_162_data[31:0]; // @[lut_35.scala 5279:33]
    end
    if (reset) begin // @[lut_35.scala 5199:41]
      read_stack23_clear <= 32'h0; // @[lut_35.scala 5199:41]
    end else begin
      read_stack23_clear <= LUT_mem_MPORT_163_data[31:0]; // @[lut_35.scala 5280:33]
    end
    if (reset) begin // @[lut_35.scala 5200:41]
      read_stack24_clear <= 32'h0; // @[lut_35.scala 5200:41]
    end else begin
      read_stack24_clear <= LUT_mem_MPORT_164_data[31:0]; // @[lut_35.scala 5281:33]
    end
    if (reset) begin // @[lut_35.scala 5201:41]
      read_stack25_clear <= 32'h0; // @[lut_35.scala 5201:41]
    end else begin
      read_stack25_clear <= LUT_mem_MPORT_165_data[31:0]; // @[lut_35.scala 5282:33]
    end
    if (reset) begin // @[lut_35.scala 5202:41]
      read_stack26_clear <= 32'h0; // @[lut_35.scala 5202:41]
    end else begin
      read_stack26_clear <= LUT_mem_MPORT_166_data[31:0]; // @[lut_35.scala 5283:33]
    end
    if (reset) begin // @[lut_35.scala 5203:41]
      read_stack27_clear <= 32'h0; // @[lut_35.scala 5203:41]
    end else begin
      read_stack27_clear <= LUT_mem_MPORT_167_data[31:0]; // @[lut_35.scala 5284:33]
    end
    if (reset) begin // @[lut_35.scala 5204:41]
      read_stack28_clear <= 32'h0; // @[lut_35.scala 5204:41]
    end else begin
      read_stack28_clear <= LUT_mem_MPORT_168_data[31:0]; // @[lut_35.scala 5285:33]
    end
    if (reset) begin // @[lut_35.scala 5205:41]
      read_stack29_clear <= 32'h0; // @[lut_35.scala 5205:41]
    end else begin
      read_stack29_clear <= LUT_mem_MPORT_169_data[31:0]; // @[lut_35.scala 5286:33]
    end
    if (reset) begin // @[lut_35.scala 5206:41]
      read_stack30_clear <= 32'h0; // @[lut_35.scala 5206:41]
    end else begin
      read_stack30_clear <= LUT_mem_MPORT_170_data[31:0]; // @[lut_35.scala 5288:33]
    end
    if (reset) begin // @[lut_35.scala 5207:41]
      read_stack31_clear <= 32'h0; // @[lut_35.scala 5207:41]
    end else begin
      read_stack31_clear <= LUT_mem_MPORT_171_data[31:0]; // @[lut_35.scala 5289:33]
    end
    if (reset) begin // @[lut_35.scala 5208:41]
      read_stack32_clear <= 32'h0; // @[lut_35.scala 5208:41]
    end else begin
      read_stack32_clear <= LUT_mem_MPORT_172_data[31:0]; // @[lut_35.scala 5290:33]
    end
    if (reset) begin // @[lut_35.scala 5209:41]
      read_stack33_clear <= 32'h0; // @[lut_35.scala 5209:41]
    end else begin
      read_stack33_clear <= LUT_mem_MPORT_173_data[31:0]; // @[lut_35.scala 5291:33]
    end
    if (reset) begin // @[lut_35.scala 5210:41]
      read_stack34_clear <= 32'h0; // @[lut_35.scala 5210:41]
    end else begin
      read_stack34_clear <= LUT_mem_MPORT_174_data[31:0]; // @[lut_35.scala 5292:33]
    end
    if (reset) begin // @[lut_35.scala 5212:39]
      clear_ray_id <= 32'h0; // @[lut_35.scala 5212:39]
    end else if (io_clear) begin // @[lut_35.scala 5295:31]
      clear_ray_id <= io_ray_id_pop; // @[lut_35.scala 5299:34]
    end
    if (reset) begin // @[lut_35.scala 5213:38]
      clear_valid <= 1'h0; // @[lut_35.scala 5213:38]
    end else begin
      clear_valid <= io_clear;
    end
    if (reset) begin // @[lut_35.scala 5216:48]
      clear_0_1 <= 1'h0; // @[lut_35.scala 5216:48]
    end else begin
      clear_0_1 <= _GEN_11392;
    end
    if (reset) begin // @[lut_35.scala 5217:48]
      clear_1_1 <= 1'h0; // @[lut_35.scala 5217:48]
    end else begin
      clear_1_1 <= _GEN_11393;
    end
    if (reset) begin // @[lut_35.scala 5218:48]
      clear_2_1 <= 1'h0; // @[lut_35.scala 5218:48]
    end else begin
      clear_2_1 <= _GEN_11394;
    end
    if (reset) begin // @[lut_35.scala 5219:48]
      clear_3_1 <= 1'h0; // @[lut_35.scala 5219:48]
    end else begin
      clear_3_1 <= _GEN_11395;
    end
    if (reset) begin // @[lut_35.scala 5220:48]
      clear_4_1 <= 1'h0; // @[lut_35.scala 5220:48]
    end else begin
      clear_4_1 <= _GEN_11396;
    end
    if (reset) begin // @[lut_35.scala 5221:48]
      clear_5_1 <= 1'h0; // @[lut_35.scala 5221:48]
    end else begin
      clear_5_1 <= _GEN_11397;
    end
    if (reset) begin // @[lut_35.scala 5222:48]
      clear_6_1 <= 1'h0; // @[lut_35.scala 5222:48]
    end else begin
      clear_6_1 <= _GEN_11398;
    end
    if (reset) begin // @[lut_35.scala 5223:48]
      clear_7_1 <= 1'h0; // @[lut_35.scala 5223:48]
    end else begin
      clear_7_1 <= _GEN_11399;
    end
    if (reset) begin // @[lut_35.scala 5224:48]
      clear_8_1 <= 1'h0; // @[lut_35.scala 5224:48]
    end else begin
      clear_8_1 <= _GEN_11400;
    end
    if (reset) begin // @[lut_35.scala 5225:48]
      clear_9_1 <= 1'h0; // @[lut_35.scala 5225:48]
    end else begin
      clear_9_1 <= _GEN_11401;
    end
    if (reset) begin // @[lut_35.scala 5226:49]
      clear_10_1 <= 1'h0; // @[lut_35.scala 5226:49]
    end else begin
      clear_10_1 <= _GEN_11402;
    end
    if (reset) begin // @[lut_35.scala 5227:49]
      clear_11_1 <= 1'h0; // @[lut_35.scala 5227:49]
    end else begin
      clear_11_1 <= _GEN_11403;
    end
    if (reset) begin // @[lut_35.scala 5228:49]
      clear_12_1 <= 1'h0; // @[lut_35.scala 5228:49]
    end else begin
      clear_12_1 <= _GEN_11404;
    end
    if (reset) begin // @[lut_35.scala 5229:49]
      clear_13_1 <= 1'h0; // @[lut_35.scala 5229:49]
    end else begin
      clear_13_1 <= _GEN_11405;
    end
    if (reset) begin // @[lut_35.scala 5230:49]
      clear_14_1 <= 1'h0; // @[lut_35.scala 5230:49]
    end else begin
      clear_14_1 <= _GEN_11406;
    end
    if (reset) begin // @[lut_35.scala 5231:49]
      clear_15_1 <= 1'h0; // @[lut_35.scala 5231:49]
    end else begin
      clear_15_1 <= _GEN_11407;
    end
    if (reset) begin // @[lut_35.scala 5232:49]
      clear_16_1 <= 1'h0; // @[lut_35.scala 5232:49]
    end else begin
      clear_16_1 <= _GEN_11408;
    end
    if (reset) begin // @[lut_35.scala 5233:49]
      clear_17_1 <= 1'h0; // @[lut_35.scala 5233:49]
    end else begin
      clear_17_1 <= _GEN_11409;
    end
    if (reset) begin // @[lut_35.scala 5234:49]
      clear_18_1 <= 1'h0; // @[lut_35.scala 5234:49]
    end else begin
      clear_18_1 <= _GEN_11410;
    end
    if (reset) begin // @[lut_35.scala 5235:49]
      clear_19_1 <= 1'h0; // @[lut_35.scala 5235:49]
    end else begin
      clear_19_1 <= _GEN_11411;
    end
    if (reset) begin // @[lut_35.scala 5236:49]
      clear_20_1 <= 1'h0; // @[lut_35.scala 5236:49]
    end else begin
      clear_20_1 <= _GEN_11412;
    end
    if (reset) begin // @[lut_35.scala 5237:49]
      clear_21_1 <= 1'h0; // @[lut_35.scala 5237:49]
    end else begin
      clear_21_1 <= _GEN_11413;
    end
    if (reset) begin // @[lut_35.scala 5238:49]
      clear_22_1 <= 1'h0; // @[lut_35.scala 5238:49]
    end else begin
      clear_22_1 <= _GEN_11414;
    end
    if (reset) begin // @[lut_35.scala 5239:49]
      clear_23_1 <= 1'h0; // @[lut_35.scala 5239:49]
    end else begin
      clear_23_1 <= _GEN_11415;
    end
    if (reset) begin // @[lut_35.scala 5240:49]
      clear_24_1 <= 1'h0; // @[lut_35.scala 5240:49]
    end else begin
      clear_24_1 <= _GEN_11416;
    end
    if (reset) begin // @[lut_35.scala 5241:49]
      clear_25_1 <= 1'h0; // @[lut_35.scala 5241:49]
    end else begin
      clear_25_1 <= _GEN_11417;
    end
    if (reset) begin // @[lut_35.scala 5242:49]
      clear_26_1 <= 1'h0; // @[lut_35.scala 5242:49]
    end else begin
      clear_26_1 <= _GEN_11418;
    end
    if (reset) begin // @[lut_35.scala 5243:49]
      clear_27_1 <= 1'h0; // @[lut_35.scala 5243:49]
    end else begin
      clear_27_1 <= _GEN_11419;
    end
    if (reset) begin // @[lut_35.scala 5244:49]
      clear_28_1 <= 1'h0; // @[lut_35.scala 5244:49]
    end else begin
      clear_28_1 <= _GEN_11420;
    end
    if (reset) begin // @[lut_35.scala 5245:49]
      clear_29_1 <= 1'h0; // @[lut_35.scala 5245:49]
    end else begin
      clear_29_1 <= _GEN_11421;
    end
    if (reset) begin // @[lut_35.scala 5246:49]
      clear_30_1 <= 1'h0; // @[lut_35.scala 5246:49]
    end else begin
      clear_30_1 <= _GEN_11422;
    end
    if (reset) begin // @[lut_35.scala 5247:49]
      clear_31_1 <= 1'h0; // @[lut_35.scala 5247:49]
    end else begin
      clear_31_1 <= _GEN_11423;
    end
    if (reset) begin // @[lut_35.scala 5248:49]
      clear_32_1 <= 1'h0; // @[lut_35.scala 5248:49]
    end else begin
      clear_32_1 <= _GEN_11424;
    end
    if (reset) begin // @[lut_35.scala 5249:49]
      clear_33_1 <= 1'h0; // @[lut_35.scala 5249:49]
    end else begin
      clear_33_1 <= _GEN_11425;
    end
    if (reset) begin // @[lut_35.scala 5250:49]
      clear_34_1 <= 1'h0; // @[lut_35.scala 5250:49]
    end else begin
      clear_34_1 <= _GEN_11426;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {2{`RANDOM}};
  _RAND_2 = {2{`RANDOM}};
  _RAND_3 = {2{`RANDOM}};
  _RAND_4 = {2{`RANDOM}};
  _RAND_5 = {2{`RANDOM}};
  _RAND_6 = {2{`RANDOM}};
  _RAND_7 = {2{`RANDOM}};
  _RAND_8 = {2{`RANDOM}};
  _RAND_9 = {2{`RANDOM}};
  _RAND_10 = {2{`RANDOM}};
  _RAND_11 = {2{`RANDOM}};
  _RAND_12 = {2{`RANDOM}};
  _RAND_13 = {2{`RANDOM}};
  _RAND_14 = {2{`RANDOM}};
  _RAND_15 = {2{`RANDOM}};
  _RAND_16 = {2{`RANDOM}};
  _RAND_17 = {2{`RANDOM}};
  _RAND_18 = {2{`RANDOM}};
  _RAND_19 = {2{`RANDOM}};
  _RAND_20 = {2{`RANDOM}};
  _RAND_21 = {2{`RANDOM}};
  _RAND_22 = {2{`RANDOM}};
  _RAND_23 = {2{`RANDOM}};
  _RAND_24 = {2{`RANDOM}};
  _RAND_25 = {2{`RANDOM}};
  _RAND_26 = {2{`RANDOM}};
  _RAND_27 = {2{`RANDOM}};
  _RAND_28 = {2{`RANDOM}};
  _RAND_29 = {2{`RANDOM}};
  _RAND_30 = {2{`RANDOM}};
  _RAND_31 = {2{`RANDOM}};
  _RAND_32 = {2{`RANDOM}};
  _RAND_33 = {2{`RANDOM}};
  _RAND_34 = {2{`RANDOM}};
  _RAND_35 = {2{`RANDOM}};
  _RAND_36 = {2{`RANDOM}};
  _RAND_37 = {2{`RANDOM}};
  _RAND_38 = {2{`RANDOM}};
  _RAND_39 = {2{`RANDOM}};
  _RAND_40 = {2{`RANDOM}};
  _RAND_41 = {2{`RANDOM}};
  _RAND_42 = {2{`RANDOM}};
  _RAND_43 = {2{`RANDOM}};
  _RAND_44 = {2{`RANDOM}};
  _RAND_45 = {2{`RANDOM}};
  _RAND_46 = {2{`RANDOM}};
  _RAND_47 = {2{`RANDOM}};
  _RAND_48 = {2{`RANDOM}};
  _RAND_49 = {2{`RANDOM}};
  _RAND_50 = {2{`RANDOM}};
  _RAND_51 = {2{`RANDOM}};
  _RAND_52 = {2{`RANDOM}};
  _RAND_53 = {2{`RANDOM}};
  _RAND_54 = {2{`RANDOM}};
  _RAND_55 = {2{`RANDOM}};
  _RAND_56 = {2{`RANDOM}};
  _RAND_57 = {2{`RANDOM}};
  _RAND_58 = {2{`RANDOM}};
  _RAND_59 = {2{`RANDOM}};
  _RAND_60 = {2{`RANDOM}};
  _RAND_61 = {2{`RANDOM}};
  _RAND_62 = {2{`RANDOM}};
  _RAND_63 = {2{`RANDOM}};
  _RAND_64 = {2{`RANDOM}};
  _RAND_65 = {2{`RANDOM}};
  _RAND_66 = {2{`RANDOM}};
  _RAND_67 = {2{`RANDOM}};
  _RAND_68 = {2{`RANDOM}};
  _RAND_69 = {2{`RANDOM}};
  _RAND_70 = {2{`RANDOM}};
  _RAND_71 = {2{`RANDOM}};
  _RAND_72 = {2{`RANDOM}};
  _RAND_73 = {2{`RANDOM}};
  _RAND_74 = {2{`RANDOM}};
  _RAND_75 = {2{`RANDOM}};
  _RAND_76 = {2{`RANDOM}};
  _RAND_77 = {2{`RANDOM}};
  _RAND_78 = {2{`RANDOM}};
  _RAND_79 = {2{`RANDOM}};
  _RAND_80 = {2{`RANDOM}};
  _RAND_81 = {2{`RANDOM}};
  _RAND_82 = {2{`RANDOM}};
  _RAND_83 = {2{`RANDOM}};
  _RAND_84 = {2{`RANDOM}};
  _RAND_85 = {2{`RANDOM}};
  _RAND_86 = {2{`RANDOM}};
  _RAND_87 = {2{`RANDOM}};
  _RAND_88 = {2{`RANDOM}};
  _RAND_89 = {2{`RANDOM}};
  _RAND_90 = {2{`RANDOM}};
  _RAND_91 = {2{`RANDOM}};
  _RAND_92 = {2{`RANDOM}};
  _RAND_93 = {2{`RANDOM}};
  _RAND_94 = {2{`RANDOM}};
  _RAND_95 = {2{`RANDOM}};
  _RAND_96 = {2{`RANDOM}};
  _RAND_97 = {2{`RANDOM}};
  _RAND_98 = {2{`RANDOM}};
  _RAND_99 = {2{`RANDOM}};
  _RAND_100 = {2{`RANDOM}};
  _RAND_101 = {2{`RANDOM}};
  _RAND_102 = {2{`RANDOM}};
  _RAND_103 = {2{`RANDOM}};
  _RAND_104 = {2{`RANDOM}};
  _RAND_105 = {2{`RANDOM}};
  _RAND_106 = {2{`RANDOM}};
  _RAND_107 = {2{`RANDOM}};
  _RAND_108 = {2{`RANDOM}};
  _RAND_109 = {2{`RANDOM}};
  _RAND_110 = {2{`RANDOM}};
  _RAND_111 = {2{`RANDOM}};
  _RAND_112 = {2{`RANDOM}};
  _RAND_113 = {2{`RANDOM}};
  _RAND_114 = {2{`RANDOM}};
  _RAND_115 = {2{`RANDOM}};
  _RAND_116 = {2{`RANDOM}};
  _RAND_117 = {2{`RANDOM}};
  _RAND_118 = {2{`RANDOM}};
  _RAND_119 = {2{`RANDOM}};
  _RAND_120 = {2{`RANDOM}};
  _RAND_121 = {2{`RANDOM}};
  _RAND_122 = {2{`RANDOM}};
  _RAND_123 = {2{`RANDOM}};
  _RAND_124 = {2{`RANDOM}};
  _RAND_125 = {2{`RANDOM}};
  _RAND_126 = {2{`RANDOM}};
  _RAND_127 = {2{`RANDOM}};
  _RAND_128 = {2{`RANDOM}};
  _RAND_129 = {2{`RANDOM}};
  _RAND_130 = {2{`RANDOM}};
  _RAND_131 = {2{`RANDOM}};
  _RAND_132 = {2{`RANDOM}};
  _RAND_133 = {2{`RANDOM}};
  _RAND_134 = {2{`RANDOM}};
  _RAND_135 = {2{`RANDOM}};
  _RAND_136 = {2{`RANDOM}};
  _RAND_137 = {2{`RANDOM}};
  _RAND_138 = {2{`RANDOM}};
  _RAND_139 = {2{`RANDOM}};
  _RAND_140 = {2{`RANDOM}};
  _RAND_141 = {2{`RANDOM}};
  _RAND_142 = {2{`RANDOM}};
  _RAND_143 = {2{`RANDOM}};
  _RAND_144 = {2{`RANDOM}};
  _RAND_145 = {2{`RANDOM}};
  _RAND_146 = {2{`RANDOM}};
  _RAND_147 = {2{`RANDOM}};
  _RAND_148 = {2{`RANDOM}};
  _RAND_149 = {2{`RANDOM}};
  _RAND_150 = {2{`RANDOM}};
  _RAND_151 = {2{`RANDOM}};
  _RAND_152 = {2{`RANDOM}};
  _RAND_153 = {2{`RANDOM}};
  _RAND_154 = {2{`RANDOM}};
  _RAND_155 = {2{`RANDOM}};
  _RAND_156 = {2{`RANDOM}};
  _RAND_157 = {2{`RANDOM}};
  _RAND_158 = {2{`RANDOM}};
  _RAND_159 = {2{`RANDOM}};
  _RAND_160 = {2{`RANDOM}};
  _RAND_161 = {2{`RANDOM}};
  _RAND_162 = {2{`RANDOM}};
  _RAND_163 = {2{`RANDOM}};
  _RAND_164 = {2{`RANDOM}};
  _RAND_165 = {2{`RANDOM}};
  _RAND_166 = {2{`RANDOM}};
  _RAND_167 = {2{`RANDOM}};
  _RAND_168 = {2{`RANDOM}};
  _RAND_169 = {2{`RANDOM}};
  _RAND_170 = {2{`RANDOM}};
  _RAND_171 = {2{`RANDOM}};
  _RAND_172 = {2{`RANDOM}};
  _RAND_173 = {2{`RANDOM}};
  _RAND_174 = {2{`RANDOM}};
  _RAND_175 = {2{`RANDOM}};
  _RAND_176 = {2{`RANDOM}};
  _RAND_177 = {2{`RANDOM}};
  _RAND_178 = {2{`RANDOM}};
  _RAND_179 = {2{`RANDOM}};
  _RAND_180 = {2{`RANDOM}};
  _RAND_181 = {2{`RANDOM}};
  _RAND_182 = {2{`RANDOM}};
  _RAND_183 = {2{`RANDOM}};
  _RAND_184 = {2{`RANDOM}};
  _RAND_185 = {2{`RANDOM}};
  _RAND_186 = {2{`RANDOM}};
  _RAND_187 = {2{`RANDOM}};
  _RAND_188 = {2{`RANDOM}};
  _RAND_189 = {2{`RANDOM}};
  _RAND_190 = {2{`RANDOM}};
  _RAND_191 = {2{`RANDOM}};
  _RAND_192 = {2{`RANDOM}};
  _RAND_193 = {2{`RANDOM}};
  _RAND_194 = {2{`RANDOM}};
  _RAND_195 = {2{`RANDOM}};
  _RAND_196 = {2{`RANDOM}};
  _RAND_197 = {2{`RANDOM}};
  _RAND_198 = {2{`RANDOM}};
  _RAND_199 = {2{`RANDOM}};
  _RAND_200 = {2{`RANDOM}};
  _RAND_201 = {2{`RANDOM}};
  _RAND_202 = {2{`RANDOM}};
  _RAND_203 = {2{`RANDOM}};
  _RAND_204 = {2{`RANDOM}};
  _RAND_205 = {2{`RANDOM}};
  _RAND_206 = {2{`RANDOM}};
  _RAND_207 = {2{`RANDOM}};
  _RAND_208 = {2{`RANDOM}};
  _RAND_209 = {2{`RANDOM}};
  _RAND_210 = {2{`RANDOM}};
  _RAND_211 = {2{`RANDOM}};
  _RAND_212 = {2{`RANDOM}};
  _RAND_213 = {2{`RANDOM}};
  _RAND_214 = {2{`RANDOM}};
  _RAND_215 = {2{`RANDOM}};
  _RAND_216 = {2{`RANDOM}};
  _RAND_217 = {2{`RANDOM}};
  _RAND_218 = {2{`RANDOM}};
  _RAND_219 = {2{`RANDOM}};
  _RAND_220 = {2{`RANDOM}};
  _RAND_221 = {2{`RANDOM}};
  _RAND_222 = {2{`RANDOM}};
  _RAND_223 = {2{`RANDOM}};
  _RAND_224 = {2{`RANDOM}};
  _RAND_225 = {2{`RANDOM}};
  _RAND_226 = {2{`RANDOM}};
  _RAND_227 = {2{`RANDOM}};
  _RAND_228 = {2{`RANDOM}};
  _RAND_229 = {2{`RANDOM}};
  _RAND_230 = {2{`RANDOM}};
  _RAND_231 = {2{`RANDOM}};
  _RAND_232 = {2{`RANDOM}};
  _RAND_233 = {2{`RANDOM}};
  _RAND_234 = {2{`RANDOM}};
  _RAND_235 = {2{`RANDOM}};
  _RAND_236 = {2{`RANDOM}};
  _RAND_237 = {2{`RANDOM}};
  _RAND_238 = {2{`RANDOM}};
  _RAND_239 = {2{`RANDOM}};
  _RAND_240 = {2{`RANDOM}};
  _RAND_241 = {2{`RANDOM}};
  _RAND_242 = {2{`RANDOM}};
  _RAND_243 = {2{`RANDOM}};
  _RAND_244 = {2{`RANDOM}};
  _RAND_245 = {2{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 35; initvar = initvar+1)
    LUT_mem[initvar] = _RAND_0[32:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  read_stack0 = _RAND_246[31:0];
  _RAND_247 = {1{`RANDOM}};
  read_stack1 = _RAND_247[31:0];
  _RAND_248 = {1{`RANDOM}};
  read_stack2 = _RAND_248[31:0];
  _RAND_249 = {1{`RANDOM}};
  read_stack3 = _RAND_249[31:0];
  _RAND_250 = {1{`RANDOM}};
  read_stack4 = _RAND_250[31:0];
  _RAND_251 = {1{`RANDOM}};
  read_stack5 = _RAND_251[31:0];
  _RAND_252 = {1{`RANDOM}};
  read_stack6 = _RAND_252[31:0];
  _RAND_253 = {1{`RANDOM}};
  read_stack7 = _RAND_253[31:0];
  _RAND_254 = {1{`RANDOM}};
  read_stack8 = _RAND_254[31:0];
  _RAND_255 = {1{`RANDOM}};
  read_stack9 = _RAND_255[31:0];
  _RAND_256 = {1{`RANDOM}};
  read_stack10 = _RAND_256[31:0];
  _RAND_257 = {1{`RANDOM}};
  read_stack11 = _RAND_257[31:0];
  _RAND_258 = {1{`RANDOM}};
  read_stack12 = _RAND_258[31:0];
  _RAND_259 = {1{`RANDOM}};
  read_stack13 = _RAND_259[31:0];
  _RAND_260 = {1{`RANDOM}};
  read_stack14 = _RAND_260[31:0];
  _RAND_261 = {1{`RANDOM}};
  read_stack15 = _RAND_261[31:0];
  _RAND_262 = {1{`RANDOM}};
  read_stack16 = _RAND_262[31:0];
  _RAND_263 = {1{`RANDOM}};
  read_stack17 = _RAND_263[31:0];
  _RAND_264 = {1{`RANDOM}};
  read_stack18 = _RAND_264[31:0];
  _RAND_265 = {1{`RANDOM}};
  read_stack19 = _RAND_265[31:0];
  _RAND_266 = {1{`RANDOM}};
  read_stack20 = _RAND_266[31:0];
  _RAND_267 = {1{`RANDOM}};
  read_stack21 = _RAND_267[31:0];
  _RAND_268 = {1{`RANDOM}};
  read_stack22 = _RAND_268[31:0];
  _RAND_269 = {1{`RANDOM}};
  read_stack23 = _RAND_269[31:0];
  _RAND_270 = {1{`RANDOM}};
  read_stack24 = _RAND_270[31:0];
  _RAND_271 = {1{`RANDOM}};
  read_stack25 = _RAND_271[31:0];
  _RAND_272 = {1{`RANDOM}};
  read_stack26 = _RAND_272[31:0];
  _RAND_273 = {1{`RANDOM}};
  read_stack27 = _RAND_273[31:0];
  _RAND_274 = {1{`RANDOM}};
  read_stack28 = _RAND_274[31:0];
  _RAND_275 = {1{`RANDOM}};
  read_stack29 = _RAND_275[31:0];
  _RAND_276 = {1{`RANDOM}};
  read_stack30 = _RAND_276[31:0];
  _RAND_277 = {1{`RANDOM}};
  read_stack31 = _RAND_277[31:0];
  _RAND_278 = {1{`RANDOM}};
  read_stack32 = _RAND_278[31:0];
  _RAND_279 = {1{`RANDOM}};
  read_stack33 = _RAND_279[31:0];
  _RAND_280 = {1{`RANDOM}};
  read_stack34 = _RAND_280[31:0];
  _RAND_281 = {1{`RANDOM}};
  push_0_1 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  push_1_1 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  push_2_1 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  push_3_1 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  push_4_1 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  push_5_1 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  push_6_1 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  push_7_1 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  push_8_1 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  push_9_1 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  push_10_1 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  push_11_1 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  push_12_1 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  push_13_1 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  push_14_1 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  push_15_1 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  push_16_1 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  push_17_1 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  push_18_1 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  push_19_1 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  push_20_1 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  push_21_1 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  push_22_1 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  push_23_1 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  push_24_1 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  push_25_1 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  push_26_1 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  push_27_1 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  push_28_1 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  push_29_1 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  push_30_1 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  push_31_1 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  push_32_1 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  push_33_1 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  push_34_1 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  push_1 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  push_valid = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  push_ray_id = _RAND_318[31:0];
  _RAND_319 = {1{`RANDOM}};
  push_valid_2 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  dispatch_reg_0 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  dispatch_reg_1 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  dispatch_reg_2 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  dispatch_reg_3 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  dispatch_reg_4 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  dispatch_reg_5 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  dispatch_reg_6 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  dispatch_reg_7 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  dispatch_reg_8 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  dispatch_reg_9 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  dispatch_reg_10 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  dispatch_reg_11 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  dispatch_reg_12 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  dispatch_reg_13 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  dispatch_reg_14 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  dispatch_reg_15 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  dispatch_reg_16 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  dispatch_reg_17 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  dispatch_reg_18 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  dispatch_reg_19 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  dispatch_reg_20 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  dispatch_reg_21 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  dispatch_reg_22 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  dispatch_reg_23 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  dispatch_reg_24 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  dispatch_reg_25 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  dispatch_reg_26 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  dispatch_reg_27 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  dispatch_reg_28 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  dispatch_reg_29 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  dispatch_reg_30 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  dispatch_reg_31 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  dispatch_reg_32 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  dispatch_reg_33 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  dispatch_reg_34 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  push_mem_temp = _RAND_355[5:0];
  _RAND_356 = {1{`RANDOM}};
  push_id_temp = _RAND_356[31:0];
  _RAND_357 = {1{`RANDOM}};
  pop_1 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  read_stack0_pop = _RAND_358[31:0];
  _RAND_359 = {1{`RANDOM}};
  read_stack1_pop = _RAND_359[31:0];
  _RAND_360 = {1{`RANDOM}};
  read_stack2_pop = _RAND_360[31:0];
  _RAND_361 = {1{`RANDOM}};
  read_stack3_pop = _RAND_361[31:0];
  _RAND_362 = {1{`RANDOM}};
  read_stack4_pop = _RAND_362[31:0];
  _RAND_363 = {1{`RANDOM}};
  read_stack5_pop = _RAND_363[31:0];
  _RAND_364 = {1{`RANDOM}};
  read_stack6_pop = _RAND_364[31:0];
  _RAND_365 = {1{`RANDOM}};
  read_stack7_pop = _RAND_365[31:0];
  _RAND_366 = {1{`RANDOM}};
  read_stack8_pop = _RAND_366[31:0];
  _RAND_367 = {1{`RANDOM}};
  read_stack9_pop = _RAND_367[31:0];
  _RAND_368 = {1{`RANDOM}};
  read_stack10_pop = _RAND_368[31:0];
  _RAND_369 = {1{`RANDOM}};
  read_stack11_pop = _RAND_369[31:0];
  _RAND_370 = {1{`RANDOM}};
  read_stack12_pop = _RAND_370[31:0];
  _RAND_371 = {1{`RANDOM}};
  read_stack13_pop = _RAND_371[31:0];
  _RAND_372 = {1{`RANDOM}};
  read_stack14_pop = _RAND_372[31:0];
  _RAND_373 = {1{`RANDOM}};
  read_stack15_pop = _RAND_373[31:0];
  _RAND_374 = {1{`RANDOM}};
  read_stack16_pop = _RAND_374[31:0];
  _RAND_375 = {1{`RANDOM}};
  read_stack17_pop = _RAND_375[31:0];
  _RAND_376 = {1{`RANDOM}};
  read_stack18_pop = _RAND_376[31:0];
  _RAND_377 = {1{`RANDOM}};
  read_stack19_pop = _RAND_377[31:0];
  _RAND_378 = {1{`RANDOM}};
  read_stack20_pop = _RAND_378[31:0];
  _RAND_379 = {1{`RANDOM}};
  read_stack21_pop = _RAND_379[31:0];
  _RAND_380 = {1{`RANDOM}};
  read_stack22_pop = _RAND_380[31:0];
  _RAND_381 = {1{`RANDOM}};
  read_stack23_pop = _RAND_381[31:0];
  _RAND_382 = {1{`RANDOM}};
  read_stack24_pop = _RAND_382[31:0];
  _RAND_383 = {1{`RANDOM}};
  read_stack25_pop = _RAND_383[31:0];
  _RAND_384 = {1{`RANDOM}};
  read_stack26_pop = _RAND_384[31:0];
  _RAND_385 = {1{`RANDOM}};
  read_stack27_pop = _RAND_385[31:0];
  _RAND_386 = {1{`RANDOM}};
  read_stack28_pop = _RAND_386[31:0];
  _RAND_387 = {1{`RANDOM}};
  read_stack29_pop = _RAND_387[31:0];
  _RAND_388 = {1{`RANDOM}};
  read_stack30_pop = _RAND_388[31:0];
  _RAND_389 = {1{`RANDOM}};
  read_stack31_pop = _RAND_389[31:0];
  _RAND_390 = {1{`RANDOM}};
  read_stack32_pop = _RAND_390[31:0];
  _RAND_391 = {1{`RANDOM}};
  read_stack33_pop = _RAND_391[31:0];
  _RAND_392 = {1{`RANDOM}};
  read_stack34_pop = _RAND_392[31:0];
  _RAND_393 = {1{`RANDOM}};
  pop_ray_id = _RAND_393[31:0];
  _RAND_394 = {1{`RANDOM}};
  pop_hitT_1 = _RAND_394[31:0];
  _RAND_395 = {1{`RANDOM}};
  pop_valid = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  pop_0_1 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  pop_1_1 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  pop_2_1 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  pop_3_1 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  pop_4_1 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  pop_5_1 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  pop_6_1 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  pop_7_1 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  pop_8_1 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  pop_9_1 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  pop_10_1 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  pop_11_1 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  pop_12_1 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  pop_13_1 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  pop_14_1 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  pop_15_1 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  pop_16_1 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  pop_17_1 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  pop_18_1 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  pop_19_1 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  pop_20_1 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  pop_21_1 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  pop_22_1 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  pop_23_1 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  pop_24_1 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  pop_25_1 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  pop_26_1 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  pop_27_1 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  pop_28_1 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  pop_29_1 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  pop_30_1 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  pop_31_1 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  pop_32_1 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  pop_33_1 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  pop_34_1 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  pop_valid_2 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  pop_ray_id_2 = _RAND_432[31:0];
  _RAND_433 = {1{`RANDOM}};
  pop_hitT_2 = _RAND_433[31:0];
  _RAND_434 = {1{`RANDOM}};
  no_match = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  no_match_1 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  no_match_2 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  clear_1 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  read_stack0_clear = _RAND_438[31:0];
  _RAND_439 = {1{`RANDOM}};
  read_stack1_clear = _RAND_439[31:0];
  _RAND_440 = {1{`RANDOM}};
  read_stack3_clear = _RAND_440[31:0];
  _RAND_441 = {1{`RANDOM}};
  read_stack4_clear = _RAND_441[31:0];
  _RAND_442 = {1{`RANDOM}};
  read_stack5_clear = _RAND_442[31:0];
  _RAND_443 = {1{`RANDOM}};
  read_stack6_clear = _RAND_443[31:0];
  _RAND_444 = {1{`RANDOM}};
  read_stack7_clear = _RAND_444[31:0];
  _RAND_445 = {1{`RANDOM}};
  read_stack8_clear = _RAND_445[31:0];
  _RAND_446 = {1{`RANDOM}};
  read_stack9_clear = _RAND_446[31:0];
  _RAND_447 = {1{`RANDOM}};
  read_stack10_clear = _RAND_447[31:0];
  _RAND_448 = {1{`RANDOM}};
  read_stack11_clear = _RAND_448[31:0];
  _RAND_449 = {1{`RANDOM}};
  read_stack12_clear = _RAND_449[31:0];
  _RAND_450 = {1{`RANDOM}};
  read_stack13_clear = _RAND_450[31:0];
  _RAND_451 = {1{`RANDOM}};
  read_stack14_clear = _RAND_451[31:0];
  _RAND_452 = {1{`RANDOM}};
  read_stack15_clear = _RAND_452[31:0];
  _RAND_453 = {1{`RANDOM}};
  read_stack16_clear = _RAND_453[31:0];
  _RAND_454 = {1{`RANDOM}};
  read_stack17_clear = _RAND_454[31:0];
  _RAND_455 = {1{`RANDOM}};
  read_stack18_clear = _RAND_455[31:0];
  _RAND_456 = {1{`RANDOM}};
  read_stack19_clear = _RAND_456[31:0];
  _RAND_457 = {1{`RANDOM}};
  read_stack20_clear = _RAND_457[31:0];
  _RAND_458 = {1{`RANDOM}};
  read_stack21_clear = _RAND_458[31:0];
  _RAND_459 = {1{`RANDOM}};
  read_stack22_clear = _RAND_459[31:0];
  _RAND_460 = {1{`RANDOM}};
  read_stack23_clear = _RAND_460[31:0];
  _RAND_461 = {1{`RANDOM}};
  read_stack24_clear = _RAND_461[31:0];
  _RAND_462 = {1{`RANDOM}};
  read_stack25_clear = _RAND_462[31:0];
  _RAND_463 = {1{`RANDOM}};
  read_stack26_clear = _RAND_463[31:0];
  _RAND_464 = {1{`RANDOM}};
  read_stack27_clear = _RAND_464[31:0];
  _RAND_465 = {1{`RANDOM}};
  read_stack28_clear = _RAND_465[31:0];
  _RAND_466 = {1{`RANDOM}};
  read_stack29_clear = _RAND_466[31:0];
  _RAND_467 = {1{`RANDOM}};
  read_stack30_clear = _RAND_467[31:0];
  _RAND_468 = {1{`RANDOM}};
  read_stack31_clear = _RAND_468[31:0];
  _RAND_469 = {1{`RANDOM}};
  read_stack32_clear = _RAND_469[31:0];
  _RAND_470 = {1{`RANDOM}};
  read_stack33_clear = _RAND_470[31:0];
  _RAND_471 = {1{`RANDOM}};
  read_stack34_clear = _RAND_471[31:0];
  _RAND_472 = {1{`RANDOM}};
  clear_ray_id = _RAND_472[31:0];
  _RAND_473 = {1{`RANDOM}};
  clear_valid = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  clear_0_1 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  clear_1_1 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  clear_2_1 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  clear_3_1 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  clear_4_1 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  clear_5_1 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  clear_6_1 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  clear_7_1 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  clear_8_1 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  clear_9_1 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  clear_10_1 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  clear_11_1 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  clear_12_1 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  clear_13_1 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  clear_14_1 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  clear_15_1 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  clear_16_1 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  clear_17_1 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  clear_18_1 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  clear_19_1 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  clear_20_1 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  clear_21_1 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  clear_22_1 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  clear_23_1 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  clear_24_1 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  clear_25_1 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  clear_26_1 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  clear_27_1 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  clear_28_1 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  clear_29_1 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  clear_30_1 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  clear_31_1 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  clear_32_1 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  clear_33_1 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  clear_34_1 = _RAND_508[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Stack(
  input         clock,
  input         reset,
  input         io_push,
  input         io_pop,
  input  [31:0] io_dataIn,
  input         io_clear,
  input  [31:0] io_ray_id,
  output [31:0] io_dataOut,
  output        io_empty,
  input  [31:0] io_hit_in,
  output [31:0] io_hit_out,
  output [31:0] io_ray_out,
  output        io_enable
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] stack_mem [0:31]; // @[stack.scala 27:24]
  wire [31:0] stack_mem_MPORT_1_data; // @[stack.scala 27:24]
  wire [4:0] stack_mem_MPORT_1_addr; // @[stack.scala 27:24]
  wire [31:0] stack_mem_MPORT_data; // @[stack.scala 27:24]
  wire [4:0] stack_mem_MPORT_addr; // @[stack.scala 27:24]
  wire  stack_mem_MPORT_mask; // @[stack.scala 27:24]
  wire  stack_mem_MPORT_en; // @[stack.scala 27:24]
  reg [5:0] sp; // @[stack.scala 28:21]
  reg [31:0] out; // @[stack.scala 29:22]
  reg [31:0] hit_1; // @[stack.scala 30:23]
  reg [31:0] ray_1; // @[stack.scala 31:23]
  reg  enable; // @[stack.scala 32:25]
  wire  _T_1 = io_push & sp < 6'h20; // @[stack.scala 39:18]
  wire  _T_2 = ~io_clear; // @[stack.scala 39:45]
  wire  _T_3 = io_push & sp < 6'h20 & ~io_clear; // @[stack.scala 39:41]
  wire [5:0] _T_6 = sp + 6'h1; // @[stack.scala 41:18]
  wire  _T_10 = io_pop & sp >= 6'h1 & _T_2; // @[stack.scala 44:37]
  wire [5:0] _T_12 = sp - 6'h1; // @[stack.scala 45:28]
  wire  _GEN_1 = io_clear | enable; // @[stack.scala 50:25 stack.scala 52:16 stack.scala 57:15]
  wire  _GEN_11 = io_pop & sp >= 6'h1 & _T_2 | _GEN_1; // @[stack.scala 44:53 stack.scala 49:16]
  assign stack_mem_MPORT_1_addr = _T_12[4:0];
  assign stack_mem_MPORT_1_data = stack_mem[stack_mem_MPORT_1_addr]; // @[stack.scala 27:24]
  assign stack_mem_MPORT_data = io_dataIn;
  assign stack_mem_MPORT_addr = sp[4:0];
  assign stack_mem_MPORT_mask = 1'h1;
  assign stack_mem_MPORT_en = _T_1 & _T_2;
  assign io_dataOut = out; // @[stack.scala 67:16]
  assign io_empty = sp == 6'h0; // @[stack.scala 66:21]
  assign io_hit_out = hit_1; // @[stack.scala 68:18]
  assign io_ray_out = ray_1; // @[stack.scala 69:21]
  assign io_enable = enable; // @[stack.scala 70:18]
  always @(posedge clock) begin
    if(stack_mem_MPORT_en & stack_mem_MPORT_mask) begin
      stack_mem[stack_mem_MPORT_addr] <= stack_mem_MPORT_data; // @[stack.scala 27:24]
    end
    if (reset) begin // @[stack.scala 28:21]
      sp <= 6'h0; // @[stack.scala 28:21]
    end else if (io_push & sp < 6'h20 & ~io_clear) begin // @[stack.scala 39:57]
      sp <= _T_6; // @[stack.scala 41:12]
    end else if (io_pop & sp >= 6'h1 & _T_2) begin // @[stack.scala 44:53]
      sp <= _T_12; // @[stack.scala 46:12]
    end else if (io_clear) begin // @[stack.scala 50:25]
      sp <= 6'h0; // @[stack.scala 51:12]
    end
    if (reset) begin // @[stack.scala 29:22]
      out <= 32'sh0; // @[stack.scala 29:22]
    end else if (!(io_push & sp < 6'h20 & ~io_clear)) begin // @[stack.scala 39:57]
      if (io_pop & sp >= 6'h1 & _T_2) begin // @[stack.scala 44:53]
        out <= stack_mem_MPORT_1_data; // @[stack.scala 45:13]
      end
    end
    if (reset) begin // @[stack.scala 30:23]
      hit_1 <= 32'h0; // @[stack.scala 30:23]
    end else if (!(io_push & sp < 6'h20 & ~io_clear)) begin // @[stack.scala 39:57]
      if (io_pop & sp >= 6'h1 & _T_2) begin // @[stack.scala 44:53]
        hit_1 <= io_hit_in; // @[stack.scala 47:15]
      end else if (!(io_clear)) begin // @[stack.scala 50:25]
        hit_1 <= 32'h0; // @[stack.scala 55:16]
      end
    end
    if (reset) begin // @[stack.scala 31:23]
      ray_1 <= 32'h0; // @[stack.scala 31:23]
    end else if (!(io_push & sp < 6'h20 & ~io_clear)) begin // @[stack.scala 39:57]
      if (io_pop & sp >= 6'h1 & _T_2) begin // @[stack.scala 44:53]
        ray_1 <= io_ray_id; // @[stack.scala 48:15]
      end else if (!(io_clear)) begin // @[stack.scala 50:25]
        ray_1 <= 32'h0; // @[stack.scala 56:15]
      end
    end
    if (reset) begin // @[stack.scala 32:25]
      enable <= 1'h0; // @[stack.scala 32:25]
    end else if (io_push & sp < 6'h20 & ~io_clear) begin // @[stack.scala 39:57]
      enable <= 1'h0; // @[stack.scala 42:15]
    end else begin
      enable <= _GEN_11;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    stack_mem[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  sp = _RAND_1[5:0];
  _RAND_2 = {1{`RANDOM}};
  out = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  hit_1 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  ray_1 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  enable = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Stackmanage(
  input         clock,
  input         reset,
  input         io_push,
  input         io_push_en,
  input         io_pop,
  input         io_pop_en,
  input  [31:0] io_ray_id_push,
  input  [31:0] io_ray_id_pop,
  input  [31:0] io_node_id_push_in,
  input  [31:0] io_hitT_in,
  input         io_clear,
  output [31:0] io_hitT_out,
  output [31:0] io_node_id_out,
  output [31:0] io_ray_id_out,
  output        io_pop_valid,
  output        io_Dis_en,
  output        io_Finish
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
`endif // RANDOMIZE_REG_INIT
  wire  LUT_stack_clock; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_reset; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_push; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_push_valid; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_pop; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_pop_valid; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_clear; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_empty_0; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_empty_1; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_empty_2; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_empty_3; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_empty_4; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_empty_5; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_empty_6; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_empty_7; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_empty_8; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_empty_9; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_empty_10; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_empty_11; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_empty_12; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_empty_13; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_empty_14; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_empty_15; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_empty_16; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_empty_17; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_empty_18; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_empty_19; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_empty_20; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_empty_21; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_empty_22; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_empty_23; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_empty_24; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_empty_25; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_empty_26; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_empty_27; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_empty_28; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_empty_29; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_empty_30; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_empty_31; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_empty_32; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_empty_33; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_empty_34; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_dispatch_0; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_dispatch_1; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_dispatch_2; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_dispatch_3; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_dispatch_4; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_dispatch_5; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_dispatch_6; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_dispatch_7; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_dispatch_8; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_dispatch_9; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_dispatch_10; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_dispatch_11; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_dispatch_12; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_dispatch_13; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_dispatch_14; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_dispatch_15; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_dispatch_16; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_dispatch_17; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_dispatch_18; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_dispatch_19; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_dispatch_20; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_dispatch_21; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_dispatch_22; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_dispatch_23; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_dispatch_24; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_dispatch_25; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_dispatch_26; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_dispatch_27; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_dispatch_28; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_dispatch_29; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_dispatch_30; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_dispatch_31; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_dispatch_32; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_dispatch_33; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_dispatch_34; // @[stackmanage_35.scala 35:45]
  wire [31:0] LUT_stack_io_ray_id_push; // @[stackmanage_35.scala 35:45]
  wire [31:0] LUT_stack_io_ray_id_pop; // @[stackmanage_35.scala 35:45]
  wire [31:0] LUT_stack_io_node_id_push_in; // @[stackmanage_35.scala 35:45]
  wire [31:0] LUT_stack_io_hitT_in; // @[stackmanage_35.scala 35:45]
  wire [31:0] LUT_stack_io_ray_id_pop_out; // @[stackmanage_35.scala 35:45]
  wire [31:0] LUT_stack_io_hitT_out; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_pop_0; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_pop_1; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_pop_2; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_pop_3; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_pop_4; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_pop_5; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_pop_6; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_pop_7; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_pop_8; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_pop_9; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_pop_10; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_pop_11; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_pop_12; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_pop_13; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_pop_14; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_pop_15; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_pop_16; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_pop_17; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_pop_18; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_pop_19; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_pop_20; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_pop_21; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_pop_22; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_pop_23; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_pop_24; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_pop_25; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_pop_26; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_pop_27; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_pop_28; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_pop_29; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_pop_30; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_pop_31; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_pop_32; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_pop_33; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_pop_34; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_pop_en; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_push_0; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_push_1; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_push_2; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_push_3; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_push_4; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_push_5; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_push_6; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_push_7; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_push_8; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_push_9; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_push_10; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_push_11; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_push_12; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_push_13; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_push_14; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_push_15; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_push_16; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_push_17; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_push_18; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_push_19; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_push_20; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_push_21; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_push_22; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_push_23; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_push_24; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_push_25; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_push_26; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_push_27; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_push_28; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_push_29; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_push_30; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_push_31; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_push_32; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_push_33; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_push_34; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_clear_0; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_clear_1; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_clear_2; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_clear_3; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_clear_4; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_clear_5; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_clear_6; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_clear_7; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_clear_8; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_clear_9; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_clear_10; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_clear_11; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_clear_12; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_clear_13; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_clear_14; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_clear_15; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_clear_16; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_clear_17; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_clear_18; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_clear_19; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_clear_20; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_clear_21; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_clear_22; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_clear_23; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_clear_24; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_clear_25; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_clear_26; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_clear_27; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_clear_28; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_clear_29; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_clear_30; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_clear_31; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_clear_32; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_clear_33; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_clear_34; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_push_en; // @[stackmanage_35.scala 35:45]
  wire  LUT_stack_io_no_match; // @[stackmanage_35.scala 35:45]
  wire  Stack_0_clock; // @[stackmanage_35.scala 36:48]
  wire  Stack_0_reset; // @[stackmanage_35.scala 36:48]
  wire  Stack_0_io_push; // @[stackmanage_35.scala 36:48]
  wire  Stack_0_io_pop; // @[stackmanage_35.scala 36:48]
  wire [31:0] Stack_0_io_dataIn; // @[stackmanage_35.scala 36:48]
  wire  Stack_0_io_clear; // @[stackmanage_35.scala 36:48]
  wire [31:0] Stack_0_io_ray_id; // @[stackmanage_35.scala 36:48]
  wire [31:0] Stack_0_io_dataOut; // @[stackmanage_35.scala 36:48]
  wire  Stack_0_io_empty; // @[stackmanage_35.scala 36:48]
  wire [31:0] Stack_0_io_hit_in; // @[stackmanage_35.scala 36:48]
  wire [31:0] Stack_0_io_hit_out; // @[stackmanage_35.scala 36:48]
  wire [31:0] Stack_0_io_ray_out; // @[stackmanage_35.scala 36:48]
  wire  Stack_0_io_enable; // @[stackmanage_35.scala 36:48]
  wire  Stack_1_clock; // @[stackmanage_35.scala 37:48]
  wire  Stack_1_reset; // @[stackmanage_35.scala 37:48]
  wire  Stack_1_io_push; // @[stackmanage_35.scala 37:48]
  wire  Stack_1_io_pop; // @[stackmanage_35.scala 37:48]
  wire [31:0] Stack_1_io_dataIn; // @[stackmanage_35.scala 37:48]
  wire  Stack_1_io_clear; // @[stackmanage_35.scala 37:48]
  wire [31:0] Stack_1_io_ray_id; // @[stackmanage_35.scala 37:48]
  wire [31:0] Stack_1_io_dataOut; // @[stackmanage_35.scala 37:48]
  wire  Stack_1_io_empty; // @[stackmanage_35.scala 37:48]
  wire [31:0] Stack_1_io_hit_in; // @[stackmanage_35.scala 37:48]
  wire [31:0] Stack_1_io_hit_out; // @[stackmanage_35.scala 37:48]
  wire [31:0] Stack_1_io_ray_out; // @[stackmanage_35.scala 37:48]
  wire  Stack_1_io_enable; // @[stackmanage_35.scala 37:48]
  wire  Stack_2_clock; // @[stackmanage_35.scala 38:48]
  wire  Stack_2_reset; // @[stackmanage_35.scala 38:48]
  wire  Stack_2_io_push; // @[stackmanage_35.scala 38:48]
  wire  Stack_2_io_pop; // @[stackmanage_35.scala 38:48]
  wire [31:0] Stack_2_io_dataIn; // @[stackmanage_35.scala 38:48]
  wire  Stack_2_io_clear; // @[stackmanage_35.scala 38:48]
  wire [31:0] Stack_2_io_ray_id; // @[stackmanage_35.scala 38:48]
  wire [31:0] Stack_2_io_dataOut; // @[stackmanage_35.scala 38:48]
  wire  Stack_2_io_empty; // @[stackmanage_35.scala 38:48]
  wire [31:0] Stack_2_io_hit_in; // @[stackmanage_35.scala 38:48]
  wire [31:0] Stack_2_io_hit_out; // @[stackmanage_35.scala 38:48]
  wire [31:0] Stack_2_io_ray_out; // @[stackmanage_35.scala 38:48]
  wire  Stack_2_io_enable; // @[stackmanage_35.scala 38:48]
  wire  Stack_3_clock; // @[stackmanage_35.scala 39:48]
  wire  Stack_3_reset; // @[stackmanage_35.scala 39:48]
  wire  Stack_3_io_push; // @[stackmanage_35.scala 39:48]
  wire  Stack_3_io_pop; // @[stackmanage_35.scala 39:48]
  wire [31:0] Stack_3_io_dataIn; // @[stackmanage_35.scala 39:48]
  wire  Stack_3_io_clear; // @[stackmanage_35.scala 39:48]
  wire [31:0] Stack_3_io_ray_id; // @[stackmanage_35.scala 39:48]
  wire [31:0] Stack_3_io_dataOut; // @[stackmanage_35.scala 39:48]
  wire  Stack_3_io_empty; // @[stackmanage_35.scala 39:48]
  wire [31:0] Stack_3_io_hit_in; // @[stackmanage_35.scala 39:48]
  wire [31:0] Stack_3_io_hit_out; // @[stackmanage_35.scala 39:48]
  wire [31:0] Stack_3_io_ray_out; // @[stackmanage_35.scala 39:48]
  wire  Stack_3_io_enable; // @[stackmanage_35.scala 39:48]
  wire  Stack_4_clock; // @[stackmanage_35.scala 40:48]
  wire  Stack_4_reset; // @[stackmanage_35.scala 40:48]
  wire  Stack_4_io_push; // @[stackmanage_35.scala 40:48]
  wire  Stack_4_io_pop; // @[stackmanage_35.scala 40:48]
  wire [31:0] Stack_4_io_dataIn; // @[stackmanage_35.scala 40:48]
  wire  Stack_4_io_clear; // @[stackmanage_35.scala 40:48]
  wire [31:0] Stack_4_io_ray_id; // @[stackmanage_35.scala 40:48]
  wire [31:0] Stack_4_io_dataOut; // @[stackmanage_35.scala 40:48]
  wire  Stack_4_io_empty; // @[stackmanage_35.scala 40:48]
  wire [31:0] Stack_4_io_hit_in; // @[stackmanage_35.scala 40:48]
  wire [31:0] Stack_4_io_hit_out; // @[stackmanage_35.scala 40:48]
  wire [31:0] Stack_4_io_ray_out; // @[stackmanage_35.scala 40:48]
  wire  Stack_4_io_enable; // @[stackmanage_35.scala 40:48]
  wire  Stack_5_clock; // @[stackmanage_35.scala 41:48]
  wire  Stack_5_reset; // @[stackmanage_35.scala 41:48]
  wire  Stack_5_io_push; // @[stackmanage_35.scala 41:48]
  wire  Stack_5_io_pop; // @[stackmanage_35.scala 41:48]
  wire [31:0] Stack_5_io_dataIn; // @[stackmanage_35.scala 41:48]
  wire  Stack_5_io_clear; // @[stackmanage_35.scala 41:48]
  wire [31:0] Stack_5_io_ray_id; // @[stackmanage_35.scala 41:48]
  wire [31:0] Stack_5_io_dataOut; // @[stackmanage_35.scala 41:48]
  wire  Stack_5_io_empty; // @[stackmanage_35.scala 41:48]
  wire [31:0] Stack_5_io_hit_in; // @[stackmanage_35.scala 41:48]
  wire [31:0] Stack_5_io_hit_out; // @[stackmanage_35.scala 41:48]
  wire [31:0] Stack_5_io_ray_out; // @[stackmanage_35.scala 41:48]
  wire  Stack_5_io_enable; // @[stackmanage_35.scala 41:48]
  wire  Stack_6_clock; // @[stackmanage_35.scala 42:48]
  wire  Stack_6_reset; // @[stackmanage_35.scala 42:48]
  wire  Stack_6_io_push; // @[stackmanage_35.scala 42:48]
  wire  Stack_6_io_pop; // @[stackmanage_35.scala 42:48]
  wire [31:0] Stack_6_io_dataIn; // @[stackmanage_35.scala 42:48]
  wire  Stack_6_io_clear; // @[stackmanage_35.scala 42:48]
  wire [31:0] Stack_6_io_ray_id; // @[stackmanage_35.scala 42:48]
  wire [31:0] Stack_6_io_dataOut; // @[stackmanage_35.scala 42:48]
  wire  Stack_6_io_empty; // @[stackmanage_35.scala 42:48]
  wire [31:0] Stack_6_io_hit_in; // @[stackmanage_35.scala 42:48]
  wire [31:0] Stack_6_io_hit_out; // @[stackmanage_35.scala 42:48]
  wire [31:0] Stack_6_io_ray_out; // @[stackmanage_35.scala 42:48]
  wire  Stack_6_io_enable; // @[stackmanage_35.scala 42:48]
  wire  Stack_7_clock; // @[stackmanage_35.scala 43:48]
  wire  Stack_7_reset; // @[stackmanage_35.scala 43:48]
  wire  Stack_7_io_push; // @[stackmanage_35.scala 43:48]
  wire  Stack_7_io_pop; // @[stackmanage_35.scala 43:48]
  wire [31:0] Stack_7_io_dataIn; // @[stackmanage_35.scala 43:48]
  wire  Stack_7_io_clear; // @[stackmanage_35.scala 43:48]
  wire [31:0] Stack_7_io_ray_id; // @[stackmanage_35.scala 43:48]
  wire [31:0] Stack_7_io_dataOut; // @[stackmanage_35.scala 43:48]
  wire  Stack_7_io_empty; // @[stackmanage_35.scala 43:48]
  wire [31:0] Stack_7_io_hit_in; // @[stackmanage_35.scala 43:48]
  wire [31:0] Stack_7_io_hit_out; // @[stackmanage_35.scala 43:48]
  wire [31:0] Stack_7_io_ray_out; // @[stackmanage_35.scala 43:48]
  wire  Stack_7_io_enable; // @[stackmanage_35.scala 43:48]
  wire  Stack_8_clock; // @[stackmanage_35.scala 44:48]
  wire  Stack_8_reset; // @[stackmanage_35.scala 44:48]
  wire  Stack_8_io_push; // @[stackmanage_35.scala 44:48]
  wire  Stack_8_io_pop; // @[stackmanage_35.scala 44:48]
  wire [31:0] Stack_8_io_dataIn; // @[stackmanage_35.scala 44:48]
  wire  Stack_8_io_clear; // @[stackmanage_35.scala 44:48]
  wire [31:0] Stack_8_io_ray_id; // @[stackmanage_35.scala 44:48]
  wire [31:0] Stack_8_io_dataOut; // @[stackmanage_35.scala 44:48]
  wire  Stack_8_io_empty; // @[stackmanage_35.scala 44:48]
  wire [31:0] Stack_8_io_hit_in; // @[stackmanage_35.scala 44:48]
  wire [31:0] Stack_8_io_hit_out; // @[stackmanage_35.scala 44:48]
  wire [31:0] Stack_8_io_ray_out; // @[stackmanage_35.scala 44:48]
  wire  Stack_8_io_enable; // @[stackmanage_35.scala 44:48]
  wire  Stack_9_clock; // @[stackmanage_35.scala 45:48]
  wire  Stack_9_reset; // @[stackmanage_35.scala 45:48]
  wire  Stack_9_io_push; // @[stackmanage_35.scala 45:48]
  wire  Stack_9_io_pop; // @[stackmanage_35.scala 45:48]
  wire [31:0] Stack_9_io_dataIn; // @[stackmanage_35.scala 45:48]
  wire  Stack_9_io_clear; // @[stackmanage_35.scala 45:48]
  wire [31:0] Stack_9_io_ray_id; // @[stackmanage_35.scala 45:48]
  wire [31:0] Stack_9_io_dataOut; // @[stackmanage_35.scala 45:48]
  wire  Stack_9_io_empty; // @[stackmanage_35.scala 45:48]
  wire [31:0] Stack_9_io_hit_in; // @[stackmanage_35.scala 45:48]
  wire [31:0] Stack_9_io_hit_out; // @[stackmanage_35.scala 45:48]
  wire [31:0] Stack_9_io_ray_out; // @[stackmanage_35.scala 45:48]
  wire  Stack_9_io_enable; // @[stackmanage_35.scala 45:48]
  wire  Stack_10_clock; // @[stackmanage_35.scala 46:47]
  wire  Stack_10_reset; // @[stackmanage_35.scala 46:47]
  wire  Stack_10_io_push; // @[stackmanage_35.scala 46:47]
  wire  Stack_10_io_pop; // @[stackmanage_35.scala 46:47]
  wire [31:0] Stack_10_io_dataIn; // @[stackmanage_35.scala 46:47]
  wire  Stack_10_io_clear; // @[stackmanage_35.scala 46:47]
  wire [31:0] Stack_10_io_ray_id; // @[stackmanage_35.scala 46:47]
  wire [31:0] Stack_10_io_dataOut; // @[stackmanage_35.scala 46:47]
  wire  Stack_10_io_empty; // @[stackmanage_35.scala 46:47]
  wire [31:0] Stack_10_io_hit_in; // @[stackmanage_35.scala 46:47]
  wire [31:0] Stack_10_io_hit_out; // @[stackmanage_35.scala 46:47]
  wire [31:0] Stack_10_io_ray_out; // @[stackmanage_35.scala 46:47]
  wire  Stack_10_io_enable; // @[stackmanage_35.scala 46:47]
  wire  Stack_11_clock; // @[stackmanage_35.scala 47:47]
  wire  Stack_11_reset; // @[stackmanage_35.scala 47:47]
  wire  Stack_11_io_push; // @[stackmanage_35.scala 47:47]
  wire  Stack_11_io_pop; // @[stackmanage_35.scala 47:47]
  wire [31:0] Stack_11_io_dataIn; // @[stackmanage_35.scala 47:47]
  wire  Stack_11_io_clear; // @[stackmanage_35.scala 47:47]
  wire [31:0] Stack_11_io_ray_id; // @[stackmanage_35.scala 47:47]
  wire [31:0] Stack_11_io_dataOut; // @[stackmanage_35.scala 47:47]
  wire  Stack_11_io_empty; // @[stackmanage_35.scala 47:47]
  wire [31:0] Stack_11_io_hit_in; // @[stackmanage_35.scala 47:47]
  wire [31:0] Stack_11_io_hit_out; // @[stackmanage_35.scala 47:47]
  wire [31:0] Stack_11_io_ray_out; // @[stackmanage_35.scala 47:47]
  wire  Stack_11_io_enable; // @[stackmanage_35.scala 47:47]
  wire  Stack_12_clock; // @[stackmanage_35.scala 48:47]
  wire  Stack_12_reset; // @[stackmanage_35.scala 48:47]
  wire  Stack_12_io_push; // @[stackmanage_35.scala 48:47]
  wire  Stack_12_io_pop; // @[stackmanage_35.scala 48:47]
  wire [31:0] Stack_12_io_dataIn; // @[stackmanage_35.scala 48:47]
  wire  Stack_12_io_clear; // @[stackmanage_35.scala 48:47]
  wire [31:0] Stack_12_io_ray_id; // @[stackmanage_35.scala 48:47]
  wire [31:0] Stack_12_io_dataOut; // @[stackmanage_35.scala 48:47]
  wire  Stack_12_io_empty; // @[stackmanage_35.scala 48:47]
  wire [31:0] Stack_12_io_hit_in; // @[stackmanage_35.scala 48:47]
  wire [31:0] Stack_12_io_hit_out; // @[stackmanage_35.scala 48:47]
  wire [31:0] Stack_12_io_ray_out; // @[stackmanage_35.scala 48:47]
  wire  Stack_12_io_enable; // @[stackmanage_35.scala 48:47]
  wire  Stack_13_clock; // @[stackmanage_35.scala 49:47]
  wire  Stack_13_reset; // @[stackmanage_35.scala 49:47]
  wire  Stack_13_io_push; // @[stackmanage_35.scala 49:47]
  wire  Stack_13_io_pop; // @[stackmanage_35.scala 49:47]
  wire [31:0] Stack_13_io_dataIn; // @[stackmanage_35.scala 49:47]
  wire  Stack_13_io_clear; // @[stackmanage_35.scala 49:47]
  wire [31:0] Stack_13_io_ray_id; // @[stackmanage_35.scala 49:47]
  wire [31:0] Stack_13_io_dataOut; // @[stackmanage_35.scala 49:47]
  wire  Stack_13_io_empty; // @[stackmanage_35.scala 49:47]
  wire [31:0] Stack_13_io_hit_in; // @[stackmanage_35.scala 49:47]
  wire [31:0] Stack_13_io_hit_out; // @[stackmanage_35.scala 49:47]
  wire [31:0] Stack_13_io_ray_out; // @[stackmanage_35.scala 49:47]
  wire  Stack_13_io_enable; // @[stackmanage_35.scala 49:47]
  wire  Stack_14_clock; // @[stackmanage_35.scala 50:47]
  wire  Stack_14_reset; // @[stackmanage_35.scala 50:47]
  wire  Stack_14_io_push; // @[stackmanage_35.scala 50:47]
  wire  Stack_14_io_pop; // @[stackmanage_35.scala 50:47]
  wire [31:0] Stack_14_io_dataIn; // @[stackmanage_35.scala 50:47]
  wire  Stack_14_io_clear; // @[stackmanage_35.scala 50:47]
  wire [31:0] Stack_14_io_ray_id; // @[stackmanage_35.scala 50:47]
  wire [31:0] Stack_14_io_dataOut; // @[stackmanage_35.scala 50:47]
  wire  Stack_14_io_empty; // @[stackmanage_35.scala 50:47]
  wire [31:0] Stack_14_io_hit_in; // @[stackmanage_35.scala 50:47]
  wire [31:0] Stack_14_io_hit_out; // @[stackmanage_35.scala 50:47]
  wire [31:0] Stack_14_io_ray_out; // @[stackmanage_35.scala 50:47]
  wire  Stack_14_io_enable; // @[stackmanage_35.scala 50:47]
  wire  Stack_15_clock; // @[stackmanage_35.scala 51:47]
  wire  Stack_15_reset; // @[stackmanage_35.scala 51:47]
  wire  Stack_15_io_push; // @[stackmanage_35.scala 51:47]
  wire  Stack_15_io_pop; // @[stackmanage_35.scala 51:47]
  wire [31:0] Stack_15_io_dataIn; // @[stackmanage_35.scala 51:47]
  wire  Stack_15_io_clear; // @[stackmanage_35.scala 51:47]
  wire [31:0] Stack_15_io_ray_id; // @[stackmanage_35.scala 51:47]
  wire [31:0] Stack_15_io_dataOut; // @[stackmanage_35.scala 51:47]
  wire  Stack_15_io_empty; // @[stackmanage_35.scala 51:47]
  wire [31:0] Stack_15_io_hit_in; // @[stackmanage_35.scala 51:47]
  wire [31:0] Stack_15_io_hit_out; // @[stackmanage_35.scala 51:47]
  wire [31:0] Stack_15_io_ray_out; // @[stackmanage_35.scala 51:47]
  wire  Stack_15_io_enable; // @[stackmanage_35.scala 51:47]
  wire  Stack_16_clock; // @[stackmanage_35.scala 52:49]
  wire  Stack_16_reset; // @[stackmanage_35.scala 52:49]
  wire  Stack_16_io_push; // @[stackmanage_35.scala 52:49]
  wire  Stack_16_io_pop; // @[stackmanage_35.scala 52:49]
  wire [31:0] Stack_16_io_dataIn; // @[stackmanage_35.scala 52:49]
  wire  Stack_16_io_clear; // @[stackmanage_35.scala 52:49]
  wire [31:0] Stack_16_io_ray_id; // @[stackmanage_35.scala 52:49]
  wire [31:0] Stack_16_io_dataOut; // @[stackmanage_35.scala 52:49]
  wire  Stack_16_io_empty; // @[stackmanage_35.scala 52:49]
  wire [31:0] Stack_16_io_hit_in; // @[stackmanage_35.scala 52:49]
  wire [31:0] Stack_16_io_hit_out; // @[stackmanage_35.scala 52:49]
  wire [31:0] Stack_16_io_ray_out; // @[stackmanage_35.scala 52:49]
  wire  Stack_16_io_enable; // @[stackmanage_35.scala 52:49]
  wire  Stack_17_clock; // @[stackmanage_35.scala 53:49]
  wire  Stack_17_reset; // @[stackmanage_35.scala 53:49]
  wire  Stack_17_io_push; // @[stackmanage_35.scala 53:49]
  wire  Stack_17_io_pop; // @[stackmanage_35.scala 53:49]
  wire [31:0] Stack_17_io_dataIn; // @[stackmanage_35.scala 53:49]
  wire  Stack_17_io_clear; // @[stackmanage_35.scala 53:49]
  wire [31:0] Stack_17_io_ray_id; // @[stackmanage_35.scala 53:49]
  wire [31:0] Stack_17_io_dataOut; // @[stackmanage_35.scala 53:49]
  wire  Stack_17_io_empty; // @[stackmanage_35.scala 53:49]
  wire [31:0] Stack_17_io_hit_in; // @[stackmanage_35.scala 53:49]
  wire [31:0] Stack_17_io_hit_out; // @[stackmanage_35.scala 53:49]
  wire [31:0] Stack_17_io_ray_out; // @[stackmanage_35.scala 53:49]
  wire  Stack_17_io_enable; // @[stackmanage_35.scala 53:49]
  wire  Stack_18_clock; // @[stackmanage_35.scala 54:49]
  wire  Stack_18_reset; // @[stackmanage_35.scala 54:49]
  wire  Stack_18_io_push; // @[stackmanage_35.scala 54:49]
  wire  Stack_18_io_pop; // @[stackmanage_35.scala 54:49]
  wire [31:0] Stack_18_io_dataIn; // @[stackmanage_35.scala 54:49]
  wire  Stack_18_io_clear; // @[stackmanage_35.scala 54:49]
  wire [31:0] Stack_18_io_ray_id; // @[stackmanage_35.scala 54:49]
  wire [31:0] Stack_18_io_dataOut; // @[stackmanage_35.scala 54:49]
  wire  Stack_18_io_empty; // @[stackmanage_35.scala 54:49]
  wire [31:0] Stack_18_io_hit_in; // @[stackmanage_35.scala 54:49]
  wire [31:0] Stack_18_io_hit_out; // @[stackmanage_35.scala 54:49]
  wire [31:0] Stack_18_io_ray_out; // @[stackmanage_35.scala 54:49]
  wire  Stack_18_io_enable; // @[stackmanage_35.scala 54:49]
  wire  Stack_19_clock; // @[stackmanage_35.scala 55:49]
  wire  Stack_19_reset; // @[stackmanage_35.scala 55:49]
  wire  Stack_19_io_push; // @[stackmanage_35.scala 55:49]
  wire  Stack_19_io_pop; // @[stackmanage_35.scala 55:49]
  wire [31:0] Stack_19_io_dataIn; // @[stackmanage_35.scala 55:49]
  wire  Stack_19_io_clear; // @[stackmanage_35.scala 55:49]
  wire [31:0] Stack_19_io_ray_id; // @[stackmanage_35.scala 55:49]
  wire [31:0] Stack_19_io_dataOut; // @[stackmanage_35.scala 55:49]
  wire  Stack_19_io_empty; // @[stackmanage_35.scala 55:49]
  wire [31:0] Stack_19_io_hit_in; // @[stackmanage_35.scala 55:49]
  wire [31:0] Stack_19_io_hit_out; // @[stackmanage_35.scala 55:49]
  wire [31:0] Stack_19_io_ray_out; // @[stackmanage_35.scala 55:49]
  wire  Stack_19_io_enable; // @[stackmanage_35.scala 55:49]
  wire  Stack_20_clock; // @[stackmanage_35.scala 56:49]
  wire  Stack_20_reset; // @[stackmanage_35.scala 56:49]
  wire  Stack_20_io_push; // @[stackmanage_35.scala 56:49]
  wire  Stack_20_io_pop; // @[stackmanage_35.scala 56:49]
  wire [31:0] Stack_20_io_dataIn; // @[stackmanage_35.scala 56:49]
  wire  Stack_20_io_clear; // @[stackmanage_35.scala 56:49]
  wire [31:0] Stack_20_io_ray_id; // @[stackmanage_35.scala 56:49]
  wire [31:0] Stack_20_io_dataOut; // @[stackmanage_35.scala 56:49]
  wire  Stack_20_io_empty; // @[stackmanage_35.scala 56:49]
  wire [31:0] Stack_20_io_hit_in; // @[stackmanage_35.scala 56:49]
  wire [31:0] Stack_20_io_hit_out; // @[stackmanage_35.scala 56:49]
  wire [31:0] Stack_20_io_ray_out; // @[stackmanage_35.scala 56:49]
  wire  Stack_20_io_enable; // @[stackmanage_35.scala 56:49]
  wire  Stack_21_clock; // @[stackmanage_35.scala 57:49]
  wire  Stack_21_reset; // @[stackmanage_35.scala 57:49]
  wire  Stack_21_io_push; // @[stackmanage_35.scala 57:49]
  wire  Stack_21_io_pop; // @[stackmanage_35.scala 57:49]
  wire [31:0] Stack_21_io_dataIn; // @[stackmanage_35.scala 57:49]
  wire  Stack_21_io_clear; // @[stackmanage_35.scala 57:49]
  wire [31:0] Stack_21_io_ray_id; // @[stackmanage_35.scala 57:49]
  wire [31:0] Stack_21_io_dataOut; // @[stackmanage_35.scala 57:49]
  wire  Stack_21_io_empty; // @[stackmanage_35.scala 57:49]
  wire [31:0] Stack_21_io_hit_in; // @[stackmanage_35.scala 57:49]
  wire [31:0] Stack_21_io_hit_out; // @[stackmanage_35.scala 57:49]
  wire [31:0] Stack_21_io_ray_out; // @[stackmanage_35.scala 57:49]
  wire  Stack_21_io_enable; // @[stackmanage_35.scala 57:49]
  wire  Stack_22_clock; // @[stackmanage_35.scala 58:49]
  wire  Stack_22_reset; // @[stackmanage_35.scala 58:49]
  wire  Stack_22_io_push; // @[stackmanage_35.scala 58:49]
  wire  Stack_22_io_pop; // @[stackmanage_35.scala 58:49]
  wire [31:0] Stack_22_io_dataIn; // @[stackmanage_35.scala 58:49]
  wire  Stack_22_io_clear; // @[stackmanage_35.scala 58:49]
  wire [31:0] Stack_22_io_ray_id; // @[stackmanage_35.scala 58:49]
  wire [31:0] Stack_22_io_dataOut; // @[stackmanage_35.scala 58:49]
  wire  Stack_22_io_empty; // @[stackmanage_35.scala 58:49]
  wire [31:0] Stack_22_io_hit_in; // @[stackmanage_35.scala 58:49]
  wire [31:0] Stack_22_io_hit_out; // @[stackmanage_35.scala 58:49]
  wire [31:0] Stack_22_io_ray_out; // @[stackmanage_35.scala 58:49]
  wire  Stack_22_io_enable; // @[stackmanage_35.scala 58:49]
  wire  Stack_23_clock; // @[stackmanage_35.scala 59:48]
  wire  Stack_23_reset; // @[stackmanage_35.scala 59:48]
  wire  Stack_23_io_push; // @[stackmanage_35.scala 59:48]
  wire  Stack_23_io_pop; // @[stackmanage_35.scala 59:48]
  wire [31:0] Stack_23_io_dataIn; // @[stackmanage_35.scala 59:48]
  wire  Stack_23_io_clear; // @[stackmanage_35.scala 59:48]
  wire [31:0] Stack_23_io_ray_id; // @[stackmanage_35.scala 59:48]
  wire [31:0] Stack_23_io_dataOut; // @[stackmanage_35.scala 59:48]
  wire  Stack_23_io_empty; // @[stackmanage_35.scala 59:48]
  wire [31:0] Stack_23_io_hit_in; // @[stackmanage_35.scala 59:48]
  wire [31:0] Stack_23_io_hit_out; // @[stackmanage_35.scala 59:48]
  wire [31:0] Stack_23_io_ray_out; // @[stackmanage_35.scala 59:48]
  wire  Stack_23_io_enable; // @[stackmanage_35.scala 59:48]
  wire  Stack_24_clock; // @[stackmanage_35.scala 60:48]
  wire  Stack_24_reset; // @[stackmanage_35.scala 60:48]
  wire  Stack_24_io_push; // @[stackmanage_35.scala 60:48]
  wire  Stack_24_io_pop; // @[stackmanage_35.scala 60:48]
  wire [31:0] Stack_24_io_dataIn; // @[stackmanage_35.scala 60:48]
  wire  Stack_24_io_clear; // @[stackmanage_35.scala 60:48]
  wire [31:0] Stack_24_io_ray_id; // @[stackmanage_35.scala 60:48]
  wire [31:0] Stack_24_io_dataOut; // @[stackmanage_35.scala 60:48]
  wire  Stack_24_io_empty; // @[stackmanage_35.scala 60:48]
  wire [31:0] Stack_24_io_hit_in; // @[stackmanage_35.scala 60:48]
  wire [31:0] Stack_24_io_hit_out; // @[stackmanage_35.scala 60:48]
  wire [31:0] Stack_24_io_ray_out; // @[stackmanage_35.scala 60:48]
  wire  Stack_24_io_enable; // @[stackmanage_35.scala 60:48]
  wire  Stack_25_clock; // @[stackmanage_35.scala 61:49]
  wire  Stack_25_reset; // @[stackmanage_35.scala 61:49]
  wire  Stack_25_io_push; // @[stackmanage_35.scala 61:49]
  wire  Stack_25_io_pop; // @[stackmanage_35.scala 61:49]
  wire [31:0] Stack_25_io_dataIn; // @[stackmanage_35.scala 61:49]
  wire  Stack_25_io_clear; // @[stackmanage_35.scala 61:49]
  wire [31:0] Stack_25_io_ray_id; // @[stackmanage_35.scala 61:49]
  wire [31:0] Stack_25_io_dataOut; // @[stackmanage_35.scala 61:49]
  wire  Stack_25_io_empty; // @[stackmanage_35.scala 61:49]
  wire [31:0] Stack_25_io_hit_in; // @[stackmanage_35.scala 61:49]
  wire [31:0] Stack_25_io_hit_out; // @[stackmanage_35.scala 61:49]
  wire [31:0] Stack_25_io_ray_out; // @[stackmanage_35.scala 61:49]
  wire  Stack_25_io_enable; // @[stackmanage_35.scala 61:49]
  wire  Stack_26_clock; // @[stackmanage_35.scala 62:47]
  wire  Stack_26_reset; // @[stackmanage_35.scala 62:47]
  wire  Stack_26_io_push; // @[stackmanage_35.scala 62:47]
  wire  Stack_26_io_pop; // @[stackmanage_35.scala 62:47]
  wire [31:0] Stack_26_io_dataIn; // @[stackmanage_35.scala 62:47]
  wire  Stack_26_io_clear; // @[stackmanage_35.scala 62:47]
  wire [31:0] Stack_26_io_ray_id; // @[stackmanage_35.scala 62:47]
  wire [31:0] Stack_26_io_dataOut; // @[stackmanage_35.scala 62:47]
  wire  Stack_26_io_empty; // @[stackmanage_35.scala 62:47]
  wire [31:0] Stack_26_io_hit_in; // @[stackmanage_35.scala 62:47]
  wire [31:0] Stack_26_io_hit_out; // @[stackmanage_35.scala 62:47]
  wire [31:0] Stack_26_io_ray_out; // @[stackmanage_35.scala 62:47]
  wire  Stack_26_io_enable; // @[stackmanage_35.scala 62:47]
  wire  Stack_27_clock; // @[stackmanage_35.scala 63:47]
  wire  Stack_27_reset; // @[stackmanage_35.scala 63:47]
  wire  Stack_27_io_push; // @[stackmanage_35.scala 63:47]
  wire  Stack_27_io_pop; // @[stackmanage_35.scala 63:47]
  wire [31:0] Stack_27_io_dataIn; // @[stackmanage_35.scala 63:47]
  wire  Stack_27_io_clear; // @[stackmanage_35.scala 63:47]
  wire [31:0] Stack_27_io_ray_id; // @[stackmanage_35.scala 63:47]
  wire [31:0] Stack_27_io_dataOut; // @[stackmanage_35.scala 63:47]
  wire  Stack_27_io_empty; // @[stackmanage_35.scala 63:47]
  wire [31:0] Stack_27_io_hit_in; // @[stackmanage_35.scala 63:47]
  wire [31:0] Stack_27_io_hit_out; // @[stackmanage_35.scala 63:47]
  wire [31:0] Stack_27_io_ray_out; // @[stackmanage_35.scala 63:47]
  wire  Stack_27_io_enable; // @[stackmanage_35.scala 63:47]
  wire  Stack_28_clock; // @[stackmanage_35.scala 64:47]
  wire  Stack_28_reset; // @[stackmanage_35.scala 64:47]
  wire  Stack_28_io_push; // @[stackmanage_35.scala 64:47]
  wire  Stack_28_io_pop; // @[stackmanage_35.scala 64:47]
  wire [31:0] Stack_28_io_dataIn; // @[stackmanage_35.scala 64:47]
  wire  Stack_28_io_clear; // @[stackmanage_35.scala 64:47]
  wire [31:0] Stack_28_io_ray_id; // @[stackmanage_35.scala 64:47]
  wire [31:0] Stack_28_io_dataOut; // @[stackmanage_35.scala 64:47]
  wire  Stack_28_io_empty; // @[stackmanage_35.scala 64:47]
  wire [31:0] Stack_28_io_hit_in; // @[stackmanage_35.scala 64:47]
  wire [31:0] Stack_28_io_hit_out; // @[stackmanage_35.scala 64:47]
  wire [31:0] Stack_28_io_ray_out; // @[stackmanage_35.scala 64:47]
  wire  Stack_28_io_enable; // @[stackmanage_35.scala 64:47]
  wire  Stack_29_clock; // @[stackmanage_35.scala 65:47]
  wire  Stack_29_reset; // @[stackmanage_35.scala 65:47]
  wire  Stack_29_io_push; // @[stackmanage_35.scala 65:47]
  wire  Stack_29_io_pop; // @[stackmanage_35.scala 65:47]
  wire [31:0] Stack_29_io_dataIn; // @[stackmanage_35.scala 65:47]
  wire  Stack_29_io_clear; // @[stackmanage_35.scala 65:47]
  wire [31:0] Stack_29_io_ray_id; // @[stackmanage_35.scala 65:47]
  wire [31:0] Stack_29_io_dataOut; // @[stackmanage_35.scala 65:47]
  wire  Stack_29_io_empty; // @[stackmanage_35.scala 65:47]
  wire [31:0] Stack_29_io_hit_in; // @[stackmanage_35.scala 65:47]
  wire [31:0] Stack_29_io_hit_out; // @[stackmanage_35.scala 65:47]
  wire [31:0] Stack_29_io_ray_out; // @[stackmanage_35.scala 65:47]
  wire  Stack_29_io_enable; // @[stackmanage_35.scala 65:47]
  wire  Stack_30_clock; // @[stackmanage_35.scala 66:47]
  wire  Stack_30_reset; // @[stackmanage_35.scala 66:47]
  wire  Stack_30_io_push; // @[stackmanage_35.scala 66:47]
  wire  Stack_30_io_pop; // @[stackmanage_35.scala 66:47]
  wire [31:0] Stack_30_io_dataIn; // @[stackmanage_35.scala 66:47]
  wire  Stack_30_io_clear; // @[stackmanage_35.scala 66:47]
  wire [31:0] Stack_30_io_ray_id; // @[stackmanage_35.scala 66:47]
  wire [31:0] Stack_30_io_dataOut; // @[stackmanage_35.scala 66:47]
  wire  Stack_30_io_empty; // @[stackmanage_35.scala 66:47]
  wire [31:0] Stack_30_io_hit_in; // @[stackmanage_35.scala 66:47]
  wire [31:0] Stack_30_io_hit_out; // @[stackmanage_35.scala 66:47]
  wire [31:0] Stack_30_io_ray_out; // @[stackmanage_35.scala 66:47]
  wire  Stack_30_io_enable; // @[stackmanage_35.scala 66:47]
  wire  Stack_31_clock; // @[stackmanage_35.scala 67:47]
  wire  Stack_31_reset; // @[stackmanage_35.scala 67:47]
  wire  Stack_31_io_push; // @[stackmanage_35.scala 67:47]
  wire  Stack_31_io_pop; // @[stackmanage_35.scala 67:47]
  wire [31:0] Stack_31_io_dataIn; // @[stackmanage_35.scala 67:47]
  wire  Stack_31_io_clear; // @[stackmanage_35.scala 67:47]
  wire [31:0] Stack_31_io_ray_id; // @[stackmanage_35.scala 67:47]
  wire [31:0] Stack_31_io_dataOut; // @[stackmanage_35.scala 67:47]
  wire  Stack_31_io_empty; // @[stackmanage_35.scala 67:47]
  wire [31:0] Stack_31_io_hit_in; // @[stackmanage_35.scala 67:47]
  wire [31:0] Stack_31_io_hit_out; // @[stackmanage_35.scala 67:47]
  wire [31:0] Stack_31_io_ray_out; // @[stackmanage_35.scala 67:47]
  wire  Stack_31_io_enable; // @[stackmanage_35.scala 67:47]
  wire  Stack_32_clock; // @[stackmanage_35.scala 68:49]
  wire  Stack_32_reset; // @[stackmanage_35.scala 68:49]
  wire  Stack_32_io_push; // @[stackmanage_35.scala 68:49]
  wire  Stack_32_io_pop; // @[stackmanage_35.scala 68:49]
  wire [31:0] Stack_32_io_dataIn; // @[stackmanage_35.scala 68:49]
  wire  Stack_32_io_clear; // @[stackmanage_35.scala 68:49]
  wire [31:0] Stack_32_io_ray_id; // @[stackmanage_35.scala 68:49]
  wire [31:0] Stack_32_io_dataOut; // @[stackmanage_35.scala 68:49]
  wire  Stack_32_io_empty; // @[stackmanage_35.scala 68:49]
  wire [31:0] Stack_32_io_hit_in; // @[stackmanage_35.scala 68:49]
  wire [31:0] Stack_32_io_hit_out; // @[stackmanage_35.scala 68:49]
  wire [31:0] Stack_32_io_ray_out; // @[stackmanage_35.scala 68:49]
  wire  Stack_32_io_enable; // @[stackmanage_35.scala 68:49]
  wire  Stack_33_clock; // @[stackmanage_35.scala 69:48]
  wire  Stack_33_reset; // @[stackmanage_35.scala 69:48]
  wire  Stack_33_io_push; // @[stackmanage_35.scala 69:48]
  wire  Stack_33_io_pop; // @[stackmanage_35.scala 69:48]
  wire [31:0] Stack_33_io_dataIn; // @[stackmanage_35.scala 69:48]
  wire  Stack_33_io_clear; // @[stackmanage_35.scala 69:48]
  wire [31:0] Stack_33_io_ray_id; // @[stackmanage_35.scala 69:48]
  wire [31:0] Stack_33_io_dataOut; // @[stackmanage_35.scala 69:48]
  wire  Stack_33_io_empty; // @[stackmanage_35.scala 69:48]
  wire [31:0] Stack_33_io_hit_in; // @[stackmanage_35.scala 69:48]
  wire [31:0] Stack_33_io_hit_out; // @[stackmanage_35.scala 69:48]
  wire [31:0] Stack_33_io_ray_out; // @[stackmanage_35.scala 69:48]
  wire  Stack_33_io_enable; // @[stackmanage_35.scala 69:48]
  wire  Stack_34_clock; // @[stackmanage_35.scala 70:48]
  wire  Stack_34_reset; // @[stackmanage_35.scala 70:48]
  wire  Stack_34_io_push; // @[stackmanage_35.scala 70:48]
  wire  Stack_34_io_pop; // @[stackmanage_35.scala 70:48]
  wire [31:0] Stack_34_io_dataIn; // @[stackmanage_35.scala 70:48]
  wire  Stack_34_io_clear; // @[stackmanage_35.scala 70:48]
  wire [31:0] Stack_34_io_ray_id; // @[stackmanage_35.scala 70:48]
  wire [31:0] Stack_34_io_dataOut; // @[stackmanage_35.scala 70:48]
  wire  Stack_34_io_empty; // @[stackmanage_35.scala 70:48]
  wire [31:0] Stack_34_io_hit_in; // @[stackmanage_35.scala 70:48]
  wire [31:0] Stack_34_io_hit_out; // @[stackmanage_35.scala 70:48]
  wire [31:0] Stack_34_io_ray_out; // @[stackmanage_35.scala 70:48]
  wire  Stack_34_io_enable; // @[stackmanage_35.scala 70:48]
  reg [31:0] node_push_in_1; // @[stackmanage_35.scala 375:34]
  reg [31:0] node_push_in_2; // @[stackmanage_35.scala 376:34]
  wire  _T_1 = LUT_stack_io_push_en; // @[stackmanage_35.scala 383:57]
  wire [31:0] _GEN_0 = LUT_stack_io_push_34 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 1607:71 stackmanage_35.scala 1608:30 stackmanage_35.scala 1678:31]
  wire [31:0] _GEN_2 = LUT_stack_io_push_33 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 1571:71 stackmanage_35.scala 1572:30]
  wire [31:0] _GEN_4 = LUT_stack_io_push_33 & _T_1 ? $signed(32'sh0) : $signed(_GEN_0); // @[stackmanage_35.scala 1571:71 stackmanage_35.scala 1606:31]
  wire [31:0] _GEN_5 = LUT_stack_io_push_32 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 1535:71 stackmanage_35.scala 1536:30]
  wire [31:0] _GEN_7 = LUT_stack_io_push_32 & _T_1 ? $signed(32'sh0) : $signed(_GEN_2); // @[stackmanage_35.scala 1535:71 stackmanage_35.scala 1569:31]
  wire [31:0] _GEN_8 = LUT_stack_io_push_32 & _T_1 ? $signed(32'sh0) : $signed(_GEN_4); // @[stackmanage_35.scala 1535:71 stackmanage_35.scala 1570:31]
  wire [31:0] _GEN_9 = LUT_stack_io_push_31 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 1499:72 stackmanage_35.scala 1500:30]
  wire [31:0] _GEN_11 = LUT_stack_io_push_31 & _T_1 ? $signed(32'sh0) : $signed(_GEN_5); // @[stackmanage_35.scala 1499:72 stackmanage_35.scala 1532:31]
  wire [31:0] _GEN_12 = LUT_stack_io_push_31 & _T_1 ? $signed(32'sh0) : $signed(_GEN_7); // @[stackmanage_35.scala 1499:72 stackmanage_35.scala 1533:31]
  wire [31:0] _GEN_13 = LUT_stack_io_push_31 & _T_1 ? $signed(32'sh0) : $signed(_GEN_8); // @[stackmanage_35.scala 1499:72 stackmanage_35.scala 1534:31]
  wire [31:0] _GEN_14 = LUT_stack_io_push_30 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 1463:72 stackmanage_35.scala 1464:30]
  wire [31:0] _GEN_16 = LUT_stack_io_push_30 & _T_1 ? $signed(32'sh0) : $signed(_GEN_9); // @[stackmanage_35.scala 1463:72 stackmanage_35.scala 1495:31]
  wire [31:0] _GEN_17 = LUT_stack_io_push_30 & _T_1 ? $signed(32'sh0) : $signed(_GEN_11); // @[stackmanage_35.scala 1463:72 stackmanage_35.scala 1496:31]
  wire [31:0] _GEN_18 = LUT_stack_io_push_30 & _T_1 ? $signed(32'sh0) : $signed(_GEN_12); // @[stackmanage_35.scala 1463:72 stackmanage_35.scala 1497:31]
  wire [31:0] _GEN_19 = LUT_stack_io_push_30 & _T_1 ? $signed(32'sh0) : $signed(_GEN_13); // @[stackmanage_35.scala 1463:72 stackmanage_35.scala 1498:31]
  wire [31:0] _GEN_20 = LUT_stack_io_push_29 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 1427:72 stackmanage_35.scala 1428:30]
  wire [31:0] _GEN_22 = LUT_stack_io_push_29 & _T_1 ? $signed(32'sh0) : $signed(_GEN_14); // @[stackmanage_35.scala 1427:72 stackmanage_35.scala 1458:31]
  wire [31:0] _GEN_23 = LUT_stack_io_push_29 & _T_1 ? $signed(32'sh0) : $signed(_GEN_16); // @[stackmanage_35.scala 1427:72 stackmanage_35.scala 1459:31]
  wire [31:0] _GEN_24 = LUT_stack_io_push_29 & _T_1 ? $signed(32'sh0) : $signed(_GEN_17); // @[stackmanage_35.scala 1427:72 stackmanage_35.scala 1460:31]
  wire [31:0] _GEN_25 = LUT_stack_io_push_29 & _T_1 ? $signed(32'sh0) : $signed(_GEN_18); // @[stackmanage_35.scala 1427:72 stackmanage_35.scala 1461:31]
  wire [31:0] _GEN_26 = LUT_stack_io_push_29 & _T_1 ? $signed(32'sh0) : $signed(_GEN_19); // @[stackmanage_35.scala 1427:72 stackmanage_35.scala 1462:31]
  wire [31:0] _GEN_27 = LUT_stack_io_push_28 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 1391:72 stackmanage_35.scala 1392:30]
  wire [31:0] _GEN_29 = LUT_stack_io_push_28 & _T_1 ? $signed(32'sh0) : $signed(_GEN_20); // @[stackmanage_35.scala 1391:72 stackmanage_35.scala 1421:31]
  wire [31:0] _GEN_30 = LUT_stack_io_push_28 & _T_1 ? $signed(32'sh0) : $signed(_GEN_22); // @[stackmanage_35.scala 1391:72 stackmanage_35.scala 1422:31]
  wire [31:0] _GEN_31 = LUT_stack_io_push_28 & _T_1 ? $signed(32'sh0) : $signed(_GEN_23); // @[stackmanage_35.scala 1391:72 stackmanage_35.scala 1423:31]
  wire [31:0] _GEN_32 = LUT_stack_io_push_28 & _T_1 ? $signed(32'sh0) : $signed(_GEN_24); // @[stackmanage_35.scala 1391:72 stackmanage_35.scala 1424:31]
  wire [31:0] _GEN_33 = LUT_stack_io_push_28 & _T_1 ? $signed(32'sh0) : $signed(_GEN_25); // @[stackmanage_35.scala 1391:72 stackmanage_35.scala 1425:31]
  wire [31:0] _GEN_34 = LUT_stack_io_push_28 & _T_1 ? $signed(32'sh0) : $signed(_GEN_26); // @[stackmanage_35.scala 1391:72 stackmanage_35.scala 1426:31]
  wire [31:0] _GEN_35 = LUT_stack_io_push_27 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 1355:72 stackmanage_35.scala 1356:30]
  wire [31:0] _GEN_37 = LUT_stack_io_push_27 & _T_1 ? $signed(32'sh0) : $signed(_GEN_27); // @[stackmanage_35.scala 1355:72 stackmanage_35.scala 1384:31]
  wire [31:0] _GEN_38 = LUT_stack_io_push_27 & _T_1 ? $signed(32'sh0) : $signed(_GEN_29); // @[stackmanage_35.scala 1355:72 stackmanage_35.scala 1385:31]
  wire [31:0] _GEN_39 = LUT_stack_io_push_27 & _T_1 ? $signed(32'sh0) : $signed(_GEN_30); // @[stackmanage_35.scala 1355:72 stackmanage_35.scala 1386:31]
  wire [31:0] _GEN_40 = LUT_stack_io_push_27 & _T_1 ? $signed(32'sh0) : $signed(_GEN_31); // @[stackmanage_35.scala 1355:72 stackmanage_35.scala 1387:31]
  wire [31:0] _GEN_41 = LUT_stack_io_push_27 & _T_1 ? $signed(32'sh0) : $signed(_GEN_32); // @[stackmanage_35.scala 1355:72 stackmanage_35.scala 1388:31]
  wire [31:0] _GEN_42 = LUT_stack_io_push_27 & _T_1 ? $signed(32'sh0) : $signed(_GEN_33); // @[stackmanage_35.scala 1355:72 stackmanage_35.scala 1389:31]
  wire [31:0] _GEN_43 = LUT_stack_io_push_27 & _T_1 ? $signed(32'sh0) : $signed(_GEN_34); // @[stackmanage_35.scala 1355:72 stackmanage_35.scala 1390:31]
  wire [31:0] _GEN_44 = LUT_stack_io_push_26 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 1319:71 stackmanage_35.scala 1320:30]
  wire [31:0] _GEN_46 = LUT_stack_io_push_26 & _T_1 ? $signed(32'sh0) : $signed(_GEN_35); // @[stackmanage_35.scala 1319:71 stackmanage_35.scala 1347:31]
  wire [31:0] _GEN_47 = LUT_stack_io_push_26 & _T_1 ? $signed(32'sh0) : $signed(_GEN_37); // @[stackmanage_35.scala 1319:71 stackmanage_35.scala 1348:31]
  wire [31:0] _GEN_48 = LUT_stack_io_push_26 & _T_1 ? $signed(32'sh0) : $signed(_GEN_38); // @[stackmanage_35.scala 1319:71 stackmanage_35.scala 1349:31]
  wire [31:0] _GEN_49 = LUT_stack_io_push_26 & _T_1 ? $signed(32'sh0) : $signed(_GEN_39); // @[stackmanage_35.scala 1319:71 stackmanage_35.scala 1350:31]
  wire [31:0] _GEN_50 = LUT_stack_io_push_26 & _T_1 ? $signed(32'sh0) : $signed(_GEN_40); // @[stackmanage_35.scala 1319:71 stackmanage_35.scala 1351:31]
  wire [31:0] _GEN_51 = LUT_stack_io_push_26 & _T_1 ? $signed(32'sh0) : $signed(_GEN_41); // @[stackmanage_35.scala 1319:71 stackmanage_35.scala 1352:31]
  wire [31:0] _GEN_52 = LUT_stack_io_push_26 & _T_1 ? $signed(32'sh0) : $signed(_GEN_42); // @[stackmanage_35.scala 1319:71 stackmanage_35.scala 1353:31]
  wire [31:0] _GEN_53 = LUT_stack_io_push_26 & _T_1 ? $signed(32'sh0) : $signed(_GEN_43); // @[stackmanage_35.scala 1319:71 stackmanage_35.scala 1354:31]
  wire [31:0] _GEN_54 = LUT_stack_io_push_25 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 1283:71 stackmanage_35.scala 1284:30]
  wire [31:0] _GEN_56 = LUT_stack_io_push_25 & _T_1 ? $signed(32'sh0) : $signed(_GEN_44); // @[stackmanage_35.scala 1283:71 stackmanage_35.scala 1310:31]
  wire [31:0] _GEN_57 = LUT_stack_io_push_25 & _T_1 ? $signed(32'sh0) : $signed(_GEN_46); // @[stackmanage_35.scala 1283:71 stackmanage_35.scala 1311:31]
  wire [31:0] _GEN_58 = LUT_stack_io_push_25 & _T_1 ? $signed(32'sh0) : $signed(_GEN_47); // @[stackmanage_35.scala 1283:71 stackmanage_35.scala 1312:31]
  wire [31:0] _GEN_59 = LUT_stack_io_push_25 & _T_1 ? $signed(32'sh0) : $signed(_GEN_48); // @[stackmanage_35.scala 1283:71 stackmanage_35.scala 1313:31]
  wire [31:0] _GEN_60 = LUT_stack_io_push_25 & _T_1 ? $signed(32'sh0) : $signed(_GEN_49); // @[stackmanage_35.scala 1283:71 stackmanage_35.scala 1314:31]
  wire [31:0] _GEN_61 = LUT_stack_io_push_25 & _T_1 ? $signed(32'sh0) : $signed(_GEN_50); // @[stackmanage_35.scala 1283:71 stackmanage_35.scala 1315:31]
  wire [31:0] _GEN_62 = LUT_stack_io_push_25 & _T_1 ? $signed(32'sh0) : $signed(_GEN_51); // @[stackmanage_35.scala 1283:71 stackmanage_35.scala 1316:31]
  wire [31:0] _GEN_63 = LUT_stack_io_push_25 & _T_1 ? $signed(32'sh0) : $signed(_GEN_52); // @[stackmanage_35.scala 1283:71 stackmanage_35.scala 1317:31]
  wire [31:0] _GEN_64 = LUT_stack_io_push_25 & _T_1 ? $signed(32'sh0) : $signed(_GEN_53); // @[stackmanage_35.scala 1283:71 stackmanage_35.scala 1318:31]
  wire [31:0] _GEN_65 = LUT_stack_io_push_24 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 1247:71 stackmanage_35.scala 1248:30]
  wire [31:0] _GEN_67 = LUT_stack_io_push_24 & _T_1 ? $signed(32'sh0) : $signed(_GEN_54); // @[stackmanage_35.scala 1247:71 stackmanage_35.scala 1273:31]
  wire [31:0] _GEN_68 = LUT_stack_io_push_24 & _T_1 ? $signed(32'sh0) : $signed(_GEN_56); // @[stackmanage_35.scala 1247:71 stackmanage_35.scala 1274:31]
  wire [31:0] _GEN_69 = LUT_stack_io_push_24 & _T_1 ? $signed(32'sh0) : $signed(_GEN_57); // @[stackmanage_35.scala 1247:71 stackmanage_35.scala 1275:31]
  wire [31:0] _GEN_70 = LUT_stack_io_push_24 & _T_1 ? $signed(32'sh0) : $signed(_GEN_58); // @[stackmanage_35.scala 1247:71 stackmanage_35.scala 1276:31]
  wire [31:0] _GEN_71 = LUT_stack_io_push_24 & _T_1 ? $signed(32'sh0) : $signed(_GEN_59); // @[stackmanage_35.scala 1247:71 stackmanage_35.scala 1277:31]
  wire [31:0] _GEN_72 = LUT_stack_io_push_24 & _T_1 ? $signed(32'sh0) : $signed(_GEN_60); // @[stackmanage_35.scala 1247:71 stackmanage_35.scala 1278:31]
  wire [31:0] _GEN_73 = LUT_stack_io_push_24 & _T_1 ? $signed(32'sh0) : $signed(_GEN_61); // @[stackmanage_35.scala 1247:71 stackmanage_35.scala 1279:31]
  wire [31:0] _GEN_74 = LUT_stack_io_push_24 & _T_1 ? $signed(32'sh0) : $signed(_GEN_62); // @[stackmanage_35.scala 1247:71 stackmanage_35.scala 1280:31]
  wire [31:0] _GEN_75 = LUT_stack_io_push_24 & _T_1 ? $signed(32'sh0) : $signed(_GEN_63); // @[stackmanage_35.scala 1247:71 stackmanage_35.scala 1281:31]
  wire [31:0] _GEN_76 = LUT_stack_io_push_24 & _T_1 ? $signed(32'sh0) : $signed(_GEN_64); // @[stackmanage_35.scala 1247:71 stackmanage_35.scala 1282:31]
  wire [31:0] _GEN_77 = LUT_stack_io_push_23 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 1211:71 stackmanage_35.scala 1212:30]
  wire [31:0] _GEN_79 = LUT_stack_io_push_23 & _T_1 ? $signed(32'sh0) : $signed(_GEN_65); // @[stackmanage_35.scala 1211:71 stackmanage_35.scala 1236:31]
  wire [31:0] _GEN_80 = LUT_stack_io_push_23 & _T_1 ? $signed(32'sh0) : $signed(_GEN_67); // @[stackmanage_35.scala 1211:71 stackmanage_35.scala 1237:31]
  wire [31:0] _GEN_81 = LUT_stack_io_push_23 & _T_1 ? $signed(32'sh0) : $signed(_GEN_68); // @[stackmanage_35.scala 1211:71 stackmanage_35.scala 1238:31]
  wire [31:0] _GEN_82 = LUT_stack_io_push_23 & _T_1 ? $signed(32'sh0) : $signed(_GEN_69); // @[stackmanage_35.scala 1211:71 stackmanage_35.scala 1239:31]
  wire [31:0] _GEN_83 = LUT_stack_io_push_23 & _T_1 ? $signed(32'sh0) : $signed(_GEN_70); // @[stackmanage_35.scala 1211:71 stackmanage_35.scala 1240:31]
  wire [31:0] _GEN_84 = LUT_stack_io_push_23 & _T_1 ? $signed(32'sh0) : $signed(_GEN_71); // @[stackmanage_35.scala 1211:71 stackmanage_35.scala 1241:31]
  wire [31:0] _GEN_85 = LUT_stack_io_push_23 & _T_1 ? $signed(32'sh0) : $signed(_GEN_72); // @[stackmanage_35.scala 1211:71 stackmanage_35.scala 1242:31]
  wire [31:0] _GEN_86 = LUT_stack_io_push_23 & _T_1 ? $signed(32'sh0) : $signed(_GEN_73); // @[stackmanage_35.scala 1211:71 stackmanage_35.scala 1243:31]
  wire [31:0] _GEN_87 = LUT_stack_io_push_23 & _T_1 ? $signed(32'sh0) : $signed(_GEN_74); // @[stackmanage_35.scala 1211:71 stackmanage_35.scala 1244:31]
  wire [31:0] _GEN_88 = LUT_stack_io_push_23 & _T_1 ? $signed(32'sh0) : $signed(_GEN_75); // @[stackmanage_35.scala 1211:71 stackmanage_35.scala 1245:31]
  wire [31:0] _GEN_89 = LUT_stack_io_push_23 & _T_1 ? $signed(32'sh0) : $signed(_GEN_76); // @[stackmanage_35.scala 1211:71 stackmanage_35.scala 1246:31]
  wire [31:0] _GEN_90 = LUT_stack_io_push_22 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 1175:71 stackmanage_35.scala 1176:30]
  wire [31:0] _GEN_92 = LUT_stack_io_push_22 & _T_1 ? $signed(32'sh0) : $signed(_GEN_77); // @[stackmanage_35.scala 1175:71 stackmanage_35.scala 1199:31]
  wire [31:0] _GEN_93 = LUT_stack_io_push_22 & _T_1 ? $signed(32'sh0) : $signed(_GEN_79); // @[stackmanage_35.scala 1175:71 stackmanage_35.scala 1200:31]
  wire [31:0] _GEN_94 = LUT_stack_io_push_22 & _T_1 ? $signed(32'sh0) : $signed(_GEN_80); // @[stackmanage_35.scala 1175:71 stackmanage_35.scala 1201:31]
  wire [31:0] _GEN_95 = LUT_stack_io_push_22 & _T_1 ? $signed(32'sh0) : $signed(_GEN_81); // @[stackmanage_35.scala 1175:71 stackmanage_35.scala 1202:31]
  wire [31:0] _GEN_96 = LUT_stack_io_push_22 & _T_1 ? $signed(32'sh0) : $signed(_GEN_82); // @[stackmanage_35.scala 1175:71 stackmanage_35.scala 1203:31]
  wire [31:0] _GEN_97 = LUT_stack_io_push_22 & _T_1 ? $signed(32'sh0) : $signed(_GEN_83); // @[stackmanage_35.scala 1175:71 stackmanage_35.scala 1204:31]
  wire [31:0] _GEN_98 = LUT_stack_io_push_22 & _T_1 ? $signed(32'sh0) : $signed(_GEN_84); // @[stackmanage_35.scala 1175:71 stackmanage_35.scala 1205:31]
  wire [31:0] _GEN_99 = LUT_stack_io_push_22 & _T_1 ? $signed(32'sh0) : $signed(_GEN_85); // @[stackmanage_35.scala 1175:71 stackmanage_35.scala 1206:31]
  wire [31:0] _GEN_100 = LUT_stack_io_push_22 & _T_1 ? $signed(32'sh0) : $signed(_GEN_86); // @[stackmanage_35.scala 1175:71 stackmanage_35.scala 1207:31]
  wire [31:0] _GEN_101 = LUT_stack_io_push_22 & _T_1 ? $signed(32'sh0) : $signed(_GEN_87); // @[stackmanage_35.scala 1175:71 stackmanage_35.scala 1208:31]
  wire [31:0] _GEN_102 = LUT_stack_io_push_22 & _T_1 ? $signed(32'sh0) : $signed(_GEN_88); // @[stackmanage_35.scala 1175:71 stackmanage_35.scala 1209:31]
  wire [31:0] _GEN_103 = LUT_stack_io_push_22 & _T_1 ? $signed(32'sh0) : $signed(_GEN_89); // @[stackmanage_35.scala 1175:71 stackmanage_35.scala 1210:31]
  wire [31:0] _GEN_104 = LUT_stack_io_push_21 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 1139:71 stackmanage_35.scala 1140:30]
  wire [31:0] _GEN_106 = LUT_stack_io_push_21 & _T_1 ? $signed(32'sh0) : $signed(_GEN_90); // @[stackmanage_35.scala 1139:71 stackmanage_35.scala 1162:31]
  wire [31:0] _GEN_107 = LUT_stack_io_push_21 & _T_1 ? $signed(32'sh0) : $signed(_GEN_92); // @[stackmanage_35.scala 1139:71 stackmanage_35.scala 1163:31]
  wire [31:0] _GEN_108 = LUT_stack_io_push_21 & _T_1 ? $signed(32'sh0) : $signed(_GEN_93); // @[stackmanage_35.scala 1139:71 stackmanage_35.scala 1164:31]
  wire [31:0] _GEN_109 = LUT_stack_io_push_21 & _T_1 ? $signed(32'sh0) : $signed(_GEN_94); // @[stackmanage_35.scala 1139:71 stackmanage_35.scala 1165:31]
  wire [31:0] _GEN_110 = LUT_stack_io_push_21 & _T_1 ? $signed(32'sh0) : $signed(_GEN_95); // @[stackmanage_35.scala 1139:71 stackmanage_35.scala 1166:31]
  wire [31:0] _GEN_111 = LUT_stack_io_push_21 & _T_1 ? $signed(32'sh0) : $signed(_GEN_96); // @[stackmanage_35.scala 1139:71 stackmanage_35.scala 1167:31]
  wire [31:0] _GEN_112 = LUT_stack_io_push_21 & _T_1 ? $signed(32'sh0) : $signed(_GEN_97); // @[stackmanage_35.scala 1139:71 stackmanage_35.scala 1168:31]
  wire [31:0] _GEN_113 = LUT_stack_io_push_21 & _T_1 ? $signed(32'sh0) : $signed(_GEN_98); // @[stackmanage_35.scala 1139:71 stackmanage_35.scala 1169:31]
  wire [31:0] _GEN_114 = LUT_stack_io_push_21 & _T_1 ? $signed(32'sh0) : $signed(_GEN_99); // @[stackmanage_35.scala 1139:71 stackmanage_35.scala 1170:31]
  wire [31:0] _GEN_115 = LUT_stack_io_push_21 & _T_1 ? $signed(32'sh0) : $signed(_GEN_100); // @[stackmanage_35.scala 1139:71 stackmanage_35.scala 1171:31]
  wire [31:0] _GEN_116 = LUT_stack_io_push_21 & _T_1 ? $signed(32'sh0) : $signed(_GEN_101); // @[stackmanage_35.scala 1139:71 stackmanage_35.scala 1172:31]
  wire [31:0] _GEN_117 = LUT_stack_io_push_21 & _T_1 ? $signed(32'sh0) : $signed(_GEN_102); // @[stackmanage_35.scala 1139:71 stackmanage_35.scala 1173:31]
  wire [31:0] _GEN_118 = LUT_stack_io_push_21 & _T_1 ? $signed(32'sh0) : $signed(_GEN_103); // @[stackmanage_35.scala 1139:71 stackmanage_35.scala 1174:31]
  wire [31:0] _GEN_119 = LUT_stack_io_push_20 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 1103:71 stackmanage_35.scala 1104:30]
  wire [31:0] _GEN_121 = LUT_stack_io_push_20 & _T_1 ? $signed(32'sh0) : $signed(_GEN_104); // @[stackmanage_35.scala 1103:71 stackmanage_35.scala 1125:31]
  wire [31:0] _GEN_122 = LUT_stack_io_push_20 & _T_1 ? $signed(32'sh0) : $signed(_GEN_106); // @[stackmanage_35.scala 1103:71 stackmanage_35.scala 1126:31]
  wire [31:0] _GEN_123 = LUT_stack_io_push_20 & _T_1 ? $signed(32'sh0) : $signed(_GEN_107); // @[stackmanage_35.scala 1103:71 stackmanage_35.scala 1127:31]
  wire [31:0] _GEN_124 = LUT_stack_io_push_20 & _T_1 ? $signed(32'sh0) : $signed(_GEN_108); // @[stackmanage_35.scala 1103:71 stackmanage_35.scala 1128:31]
  wire [31:0] _GEN_125 = LUT_stack_io_push_20 & _T_1 ? $signed(32'sh0) : $signed(_GEN_109); // @[stackmanage_35.scala 1103:71 stackmanage_35.scala 1129:31]
  wire [31:0] _GEN_126 = LUT_stack_io_push_20 & _T_1 ? $signed(32'sh0) : $signed(_GEN_110); // @[stackmanage_35.scala 1103:71 stackmanage_35.scala 1130:31]
  wire [31:0] _GEN_127 = LUT_stack_io_push_20 & _T_1 ? $signed(32'sh0) : $signed(_GEN_111); // @[stackmanage_35.scala 1103:71 stackmanage_35.scala 1131:31]
  wire [31:0] _GEN_128 = LUT_stack_io_push_20 & _T_1 ? $signed(32'sh0) : $signed(_GEN_112); // @[stackmanage_35.scala 1103:71 stackmanage_35.scala 1132:31]
  wire [31:0] _GEN_129 = LUT_stack_io_push_20 & _T_1 ? $signed(32'sh0) : $signed(_GEN_113); // @[stackmanage_35.scala 1103:71 stackmanage_35.scala 1133:31]
  wire [31:0] _GEN_130 = LUT_stack_io_push_20 & _T_1 ? $signed(32'sh0) : $signed(_GEN_114); // @[stackmanage_35.scala 1103:71 stackmanage_35.scala 1134:31]
  wire [31:0] _GEN_131 = LUT_stack_io_push_20 & _T_1 ? $signed(32'sh0) : $signed(_GEN_115); // @[stackmanage_35.scala 1103:71 stackmanage_35.scala 1135:31]
  wire [31:0] _GEN_132 = LUT_stack_io_push_20 & _T_1 ? $signed(32'sh0) : $signed(_GEN_116); // @[stackmanage_35.scala 1103:71 stackmanage_35.scala 1136:31]
  wire [31:0] _GEN_133 = LUT_stack_io_push_20 & _T_1 ? $signed(32'sh0) : $signed(_GEN_117); // @[stackmanage_35.scala 1103:71 stackmanage_35.scala 1137:31]
  wire [31:0] _GEN_134 = LUT_stack_io_push_20 & _T_1 ? $signed(32'sh0) : $signed(_GEN_118); // @[stackmanage_35.scala 1103:71 stackmanage_35.scala 1138:31]
  wire [31:0] _GEN_135 = LUT_stack_io_push_19 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 1067:71 stackmanage_35.scala 1068:30]
  wire [31:0] _GEN_137 = LUT_stack_io_push_19 & _T_1 ? $signed(32'sh0) : $signed(_GEN_119); // @[stackmanage_35.scala 1067:71 stackmanage_35.scala 1088:31]
  wire [31:0] _GEN_138 = LUT_stack_io_push_19 & _T_1 ? $signed(32'sh0) : $signed(_GEN_121); // @[stackmanage_35.scala 1067:71 stackmanage_35.scala 1089:31]
  wire [31:0] _GEN_139 = LUT_stack_io_push_19 & _T_1 ? $signed(32'sh0) : $signed(_GEN_122); // @[stackmanage_35.scala 1067:71 stackmanage_35.scala 1090:31]
  wire [31:0] _GEN_140 = LUT_stack_io_push_19 & _T_1 ? $signed(32'sh0) : $signed(_GEN_123); // @[stackmanage_35.scala 1067:71 stackmanage_35.scala 1091:31]
  wire [31:0] _GEN_141 = LUT_stack_io_push_19 & _T_1 ? $signed(32'sh0) : $signed(_GEN_124); // @[stackmanage_35.scala 1067:71 stackmanage_35.scala 1092:31]
  wire [31:0] _GEN_142 = LUT_stack_io_push_19 & _T_1 ? $signed(32'sh0) : $signed(_GEN_125); // @[stackmanage_35.scala 1067:71 stackmanage_35.scala 1093:31]
  wire [31:0] _GEN_143 = LUT_stack_io_push_19 & _T_1 ? $signed(32'sh0) : $signed(_GEN_126); // @[stackmanage_35.scala 1067:71 stackmanage_35.scala 1094:31]
  wire [31:0] _GEN_144 = LUT_stack_io_push_19 & _T_1 ? $signed(32'sh0) : $signed(_GEN_127); // @[stackmanage_35.scala 1067:71 stackmanage_35.scala 1095:31]
  wire [31:0] _GEN_145 = LUT_stack_io_push_19 & _T_1 ? $signed(32'sh0) : $signed(_GEN_128); // @[stackmanage_35.scala 1067:71 stackmanage_35.scala 1096:31]
  wire [31:0] _GEN_146 = LUT_stack_io_push_19 & _T_1 ? $signed(32'sh0) : $signed(_GEN_129); // @[stackmanage_35.scala 1067:71 stackmanage_35.scala 1097:31]
  wire [31:0] _GEN_147 = LUT_stack_io_push_19 & _T_1 ? $signed(32'sh0) : $signed(_GEN_130); // @[stackmanage_35.scala 1067:71 stackmanage_35.scala 1098:31]
  wire [31:0] _GEN_148 = LUT_stack_io_push_19 & _T_1 ? $signed(32'sh0) : $signed(_GEN_131); // @[stackmanage_35.scala 1067:71 stackmanage_35.scala 1099:31]
  wire [31:0] _GEN_149 = LUT_stack_io_push_19 & _T_1 ? $signed(32'sh0) : $signed(_GEN_132); // @[stackmanage_35.scala 1067:71 stackmanage_35.scala 1100:31]
  wire [31:0] _GEN_150 = LUT_stack_io_push_19 & _T_1 ? $signed(32'sh0) : $signed(_GEN_133); // @[stackmanage_35.scala 1067:71 stackmanage_35.scala 1101:31]
  wire [31:0] _GEN_151 = LUT_stack_io_push_19 & _T_1 ? $signed(32'sh0) : $signed(_GEN_134); // @[stackmanage_35.scala 1067:71 stackmanage_35.scala 1102:31]
  wire [31:0] _GEN_152 = LUT_stack_io_push_18 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 1031:71 stackmanage_35.scala 1032:30]
  wire [31:0] _GEN_154 = LUT_stack_io_push_18 & _T_1 ? $signed(32'sh0) : $signed(_GEN_135); // @[stackmanage_35.scala 1031:71 stackmanage_35.scala 1051:31]
  wire [31:0] _GEN_155 = LUT_stack_io_push_18 & _T_1 ? $signed(32'sh0) : $signed(_GEN_137); // @[stackmanage_35.scala 1031:71 stackmanage_35.scala 1052:31]
  wire [31:0] _GEN_156 = LUT_stack_io_push_18 & _T_1 ? $signed(32'sh0) : $signed(_GEN_138); // @[stackmanage_35.scala 1031:71 stackmanage_35.scala 1053:31]
  wire [31:0] _GEN_157 = LUT_stack_io_push_18 & _T_1 ? $signed(32'sh0) : $signed(_GEN_139); // @[stackmanage_35.scala 1031:71 stackmanage_35.scala 1054:31]
  wire [31:0] _GEN_158 = LUT_stack_io_push_18 & _T_1 ? $signed(32'sh0) : $signed(_GEN_140); // @[stackmanage_35.scala 1031:71 stackmanage_35.scala 1055:31]
  wire [31:0] _GEN_159 = LUT_stack_io_push_18 & _T_1 ? $signed(32'sh0) : $signed(_GEN_141); // @[stackmanage_35.scala 1031:71 stackmanage_35.scala 1056:31]
  wire [31:0] _GEN_160 = LUT_stack_io_push_18 & _T_1 ? $signed(32'sh0) : $signed(_GEN_142); // @[stackmanage_35.scala 1031:71 stackmanage_35.scala 1057:31]
  wire [31:0] _GEN_161 = LUT_stack_io_push_18 & _T_1 ? $signed(32'sh0) : $signed(_GEN_143); // @[stackmanage_35.scala 1031:71 stackmanage_35.scala 1058:31]
  wire [31:0] _GEN_162 = LUT_stack_io_push_18 & _T_1 ? $signed(32'sh0) : $signed(_GEN_144); // @[stackmanage_35.scala 1031:71 stackmanage_35.scala 1059:31]
  wire [31:0] _GEN_163 = LUT_stack_io_push_18 & _T_1 ? $signed(32'sh0) : $signed(_GEN_145); // @[stackmanage_35.scala 1031:71 stackmanage_35.scala 1060:31]
  wire [31:0] _GEN_164 = LUT_stack_io_push_18 & _T_1 ? $signed(32'sh0) : $signed(_GEN_146); // @[stackmanage_35.scala 1031:71 stackmanage_35.scala 1061:31]
  wire [31:0] _GEN_165 = LUT_stack_io_push_18 & _T_1 ? $signed(32'sh0) : $signed(_GEN_147); // @[stackmanage_35.scala 1031:71 stackmanage_35.scala 1062:31]
  wire [31:0] _GEN_166 = LUT_stack_io_push_18 & _T_1 ? $signed(32'sh0) : $signed(_GEN_148); // @[stackmanage_35.scala 1031:71 stackmanage_35.scala 1063:31]
  wire [31:0] _GEN_167 = LUT_stack_io_push_18 & _T_1 ? $signed(32'sh0) : $signed(_GEN_149); // @[stackmanage_35.scala 1031:71 stackmanage_35.scala 1064:31]
  wire [31:0] _GEN_168 = LUT_stack_io_push_18 & _T_1 ? $signed(32'sh0) : $signed(_GEN_150); // @[stackmanage_35.scala 1031:71 stackmanage_35.scala 1065:31]
  wire [31:0] _GEN_169 = LUT_stack_io_push_18 & _T_1 ? $signed(32'sh0) : $signed(_GEN_151); // @[stackmanage_35.scala 1031:71 stackmanage_35.scala 1066:31]
  wire [31:0] _GEN_170 = LUT_stack_io_push_17 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 995:71 stackmanage_35.scala 996:30]
  wire [31:0] _GEN_172 = LUT_stack_io_push_17 & _T_1 ? $signed(32'sh0) : $signed(_GEN_152); // @[stackmanage_35.scala 995:71 stackmanage_35.scala 1014:31]
  wire [31:0] _GEN_173 = LUT_stack_io_push_17 & _T_1 ? $signed(32'sh0) : $signed(_GEN_154); // @[stackmanage_35.scala 995:71 stackmanage_35.scala 1015:31]
  wire [31:0] _GEN_174 = LUT_stack_io_push_17 & _T_1 ? $signed(32'sh0) : $signed(_GEN_155); // @[stackmanage_35.scala 995:71 stackmanage_35.scala 1016:31]
  wire [31:0] _GEN_175 = LUT_stack_io_push_17 & _T_1 ? $signed(32'sh0) : $signed(_GEN_156); // @[stackmanage_35.scala 995:71 stackmanage_35.scala 1017:31]
  wire [31:0] _GEN_176 = LUT_stack_io_push_17 & _T_1 ? $signed(32'sh0) : $signed(_GEN_157); // @[stackmanage_35.scala 995:71 stackmanage_35.scala 1018:31]
  wire [31:0] _GEN_177 = LUT_stack_io_push_17 & _T_1 ? $signed(32'sh0) : $signed(_GEN_158); // @[stackmanage_35.scala 995:71 stackmanage_35.scala 1019:31]
  wire [31:0] _GEN_178 = LUT_stack_io_push_17 & _T_1 ? $signed(32'sh0) : $signed(_GEN_159); // @[stackmanage_35.scala 995:71 stackmanage_35.scala 1020:31]
  wire [31:0] _GEN_179 = LUT_stack_io_push_17 & _T_1 ? $signed(32'sh0) : $signed(_GEN_160); // @[stackmanage_35.scala 995:71 stackmanage_35.scala 1021:31]
  wire [31:0] _GEN_180 = LUT_stack_io_push_17 & _T_1 ? $signed(32'sh0) : $signed(_GEN_161); // @[stackmanage_35.scala 995:71 stackmanage_35.scala 1022:31]
  wire [31:0] _GEN_181 = LUT_stack_io_push_17 & _T_1 ? $signed(32'sh0) : $signed(_GEN_162); // @[stackmanage_35.scala 995:71 stackmanage_35.scala 1023:31]
  wire [31:0] _GEN_182 = LUT_stack_io_push_17 & _T_1 ? $signed(32'sh0) : $signed(_GEN_163); // @[stackmanage_35.scala 995:71 stackmanage_35.scala 1024:31]
  wire [31:0] _GEN_183 = LUT_stack_io_push_17 & _T_1 ? $signed(32'sh0) : $signed(_GEN_164); // @[stackmanage_35.scala 995:71 stackmanage_35.scala 1025:31]
  wire [31:0] _GEN_184 = LUT_stack_io_push_17 & _T_1 ? $signed(32'sh0) : $signed(_GEN_165); // @[stackmanage_35.scala 995:71 stackmanage_35.scala 1026:31]
  wire [31:0] _GEN_185 = LUT_stack_io_push_17 & _T_1 ? $signed(32'sh0) : $signed(_GEN_166); // @[stackmanage_35.scala 995:71 stackmanage_35.scala 1027:31]
  wire [31:0] _GEN_186 = LUT_stack_io_push_17 & _T_1 ? $signed(32'sh0) : $signed(_GEN_167); // @[stackmanage_35.scala 995:71 stackmanage_35.scala 1028:31]
  wire [31:0] _GEN_187 = LUT_stack_io_push_17 & _T_1 ? $signed(32'sh0) : $signed(_GEN_168); // @[stackmanage_35.scala 995:71 stackmanage_35.scala 1029:31]
  wire [31:0] _GEN_188 = LUT_stack_io_push_17 & _T_1 ? $signed(32'sh0) : $signed(_GEN_169); // @[stackmanage_35.scala 995:71 stackmanage_35.scala 1030:31]
  wire [31:0] _GEN_189 = LUT_stack_io_push_16 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 959:71 stackmanage_35.scala 960:30]
  wire [31:0] _GEN_191 = LUT_stack_io_push_16 & _T_1 ? $signed(32'sh0) : $signed(_GEN_170); // @[stackmanage_35.scala 959:71 stackmanage_35.scala 977:31]
  wire [31:0] _GEN_192 = LUT_stack_io_push_16 & _T_1 ? $signed(32'sh0) : $signed(_GEN_172); // @[stackmanage_35.scala 959:71 stackmanage_35.scala 978:31]
  wire [31:0] _GEN_193 = LUT_stack_io_push_16 & _T_1 ? $signed(32'sh0) : $signed(_GEN_173); // @[stackmanage_35.scala 959:71 stackmanage_35.scala 979:31]
  wire [31:0] _GEN_194 = LUT_stack_io_push_16 & _T_1 ? $signed(32'sh0) : $signed(_GEN_174); // @[stackmanage_35.scala 959:71 stackmanage_35.scala 980:31]
  wire [31:0] _GEN_195 = LUT_stack_io_push_16 & _T_1 ? $signed(32'sh0) : $signed(_GEN_175); // @[stackmanage_35.scala 959:71 stackmanage_35.scala 981:31]
  wire [31:0] _GEN_196 = LUT_stack_io_push_16 & _T_1 ? $signed(32'sh0) : $signed(_GEN_176); // @[stackmanage_35.scala 959:71 stackmanage_35.scala 982:31]
  wire [31:0] _GEN_197 = LUT_stack_io_push_16 & _T_1 ? $signed(32'sh0) : $signed(_GEN_177); // @[stackmanage_35.scala 959:71 stackmanage_35.scala 983:31]
  wire [31:0] _GEN_198 = LUT_stack_io_push_16 & _T_1 ? $signed(32'sh0) : $signed(_GEN_178); // @[stackmanage_35.scala 959:71 stackmanage_35.scala 984:31]
  wire [31:0] _GEN_199 = LUT_stack_io_push_16 & _T_1 ? $signed(32'sh0) : $signed(_GEN_179); // @[stackmanage_35.scala 959:71 stackmanage_35.scala 985:31]
  wire [31:0] _GEN_200 = LUT_stack_io_push_16 & _T_1 ? $signed(32'sh0) : $signed(_GEN_180); // @[stackmanage_35.scala 959:71 stackmanage_35.scala 986:31]
  wire [31:0] _GEN_201 = LUT_stack_io_push_16 & _T_1 ? $signed(32'sh0) : $signed(_GEN_181); // @[stackmanage_35.scala 959:71 stackmanage_35.scala 987:31]
  wire [31:0] _GEN_202 = LUT_stack_io_push_16 & _T_1 ? $signed(32'sh0) : $signed(_GEN_182); // @[stackmanage_35.scala 959:71 stackmanage_35.scala 988:31]
  wire [31:0] _GEN_203 = LUT_stack_io_push_16 & _T_1 ? $signed(32'sh0) : $signed(_GEN_183); // @[stackmanage_35.scala 959:71 stackmanage_35.scala 989:31]
  wire [31:0] _GEN_204 = LUT_stack_io_push_16 & _T_1 ? $signed(32'sh0) : $signed(_GEN_184); // @[stackmanage_35.scala 959:71 stackmanage_35.scala 990:31]
  wire [31:0] _GEN_205 = LUT_stack_io_push_16 & _T_1 ? $signed(32'sh0) : $signed(_GEN_185); // @[stackmanage_35.scala 959:71 stackmanage_35.scala 991:31]
  wire [31:0] _GEN_206 = LUT_stack_io_push_16 & _T_1 ? $signed(32'sh0) : $signed(_GEN_186); // @[stackmanage_35.scala 959:71 stackmanage_35.scala 992:31]
  wire [31:0] _GEN_207 = LUT_stack_io_push_16 & _T_1 ? $signed(32'sh0) : $signed(_GEN_187); // @[stackmanage_35.scala 959:71 stackmanage_35.scala 993:31]
  wire [31:0] _GEN_208 = LUT_stack_io_push_16 & _T_1 ? $signed(32'sh0) : $signed(_GEN_188); // @[stackmanage_35.scala 959:71 stackmanage_35.scala 994:31]
  wire [31:0] _GEN_209 = LUT_stack_io_push_15 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 923:71 stackmanage_35.scala 924:30]
  wire [31:0] _GEN_211 = LUT_stack_io_push_15 & _T_1 ? $signed(32'sh0) : $signed(_GEN_189); // @[stackmanage_35.scala 923:71 stackmanage_35.scala 940:31]
  wire [31:0] _GEN_212 = LUT_stack_io_push_15 & _T_1 ? $signed(32'sh0) : $signed(_GEN_191); // @[stackmanage_35.scala 923:71 stackmanage_35.scala 941:31]
  wire [31:0] _GEN_213 = LUT_stack_io_push_15 & _T_1 ? $signed(32'sh0) : $signed(_GEN_192); // @[stackmanage_35.scala 923:71 stackmanage_35.scala 942:31]
  wire [31:0] _GEN_214 = LUT_stack_io_push_15 & _T_1 ? $signed(32'sh0) : $signed(_GEN_193); // @[stackmanage_35.scala 923:71 stackmanage_35.scala 943:31]
  wire [31:0] _GEN_215 = LUT_stack_io_push_15 & _T_1 ? $signed(32'sh0) : $signed(_GEN_194); // @[stackmanage_35.scala 923:71 stackmanage_35.scala 944:31]
  wire [31:0] _GEN_216 = LUT_stack_io_push_15 & _T_1 ? $signed(32'sh0) : $signed(_GEN_195); // @[stackmanage_35.scala 923:71 stackmanage_35.scala 945:31]
  wire [31:0] _GEN_217 = LUT_stack_io_push_15 & _T_1 ? $signed(32'sh0) : $signed(_GEN_196); // @[stackmanage_35.scala 923:71 stackmanage_35.scala 946:31]
  wire [31:0] _GEN_218 = LUT_stack_io_push_15 & _T_1 ? $signed(32'sh0) : $signed(_GEN_197); // @[stackmanage_35.scala 923:71 stackmanage_35.scala 947:31]
  wire [31:0] _GEN_219 = LUT_stack_io_push_15 & _T_1 ? $signed(32'sh0) : $signed(_GEN_198); // @[stackmanage_35.scala 923:71 stackmanage_35.scala 948:31]
  wire [31:0] _GEN_220 = LUT_stack_io_push_15 & _T_1 ? $signed(32'sh0) : $signed(_GEN_199); // @[stackmanage_35.scala 923:71 stackmanage_35.scala 949:31]
  wire [31:0] _GEN_221 = LUT_stack_io_push_15 & _T_1 ? $signed(32'sh0) : $signed(_GEN_200); // @[stackmanage_35.scala 923:71 stackmanage_35.scala 950:31]
  wire [31:0] _GEN_222 = LUT_stack_io_push_15 & _T_1 ? $signed(32'sh0) : $signed(_GEN_201); // @[stackmanage_35.scala 923:71 stackmanage_35.scala 951:31]
  wire [31:0] _GEN_223 = LUT_stack_io_push_15 & _T_1 ? $signed(32'sh0) : $signed(_GEN_202); // @[stackmanage_35.scala 923:71 stackmanage_35.scala 952:31]
  wire [31:0] _GEN_224 = LUT_stack_io_push_15 & _T_1 ? $signed(32'sh0) : $signed(_GEN_203); // @[stackmanage_35.scala 923:71 stackmanage_35.scala 953:31]
  wire [31:0] _GEN_225 = LUT_stack_io_push_15 & _T_1 ? $signed(32'sh0) : $signed(_GEN_204); // @[stackmanage_35.scala 923:71 stackmanage_35.scala 954:31]
  wire [31:0] _GEN_226 = LUT_stack_io_push_15 & _T_1 ? $signed(32'sh0) : $signed(_GEN_205); // @[stackmanage_35.scala 923:71 stackmanage_35.scala 955:31]
  wire [31:0] _GEN_227 = LUT_stack_io_push_15 & _T_1 ? $signed(32'sh0) : $signed(_GEN_206); // @[stackmanage_35.scala 923:71 stackmanage_35.scala 956:31]
  wire [31:0] _GEN_228 = LUT_stack_io_push_15 & _T_1 ? $signed(32'sh0) : $signed(_GEN_207); // @[stackmanage_35.scala 923:71 stackmanage_35.scala 957:31]
  wire [31:0] _GEN_229 = LUT_stack_io_push_15 & _T_1 ? $signed(32'sh0) : $signed(_GEN_208); // @[stackmanage_35.scala 923:71 stackmanage_35.scala 958:31]
  wire [31:0] _GEN_230 = LUT_stack_io_push_14 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 887:71 stackmanage_35.scala 888:30]
  wire [31:0] _GEN_232 = LUT_stack_io_push_14 & _T_1 ? $signed(32'sh0) : $signed(_GEN_209); // @[stackmanage_35.scala 887:71 stackmanage_35.scala 903:31]
  wire [31:0] _GEN_233 = LUT_stack_io_push_14 & _T_1 ? $signed(32'sh0) : $signed(_GEN_211); // @[stackmanage_35.scala 887:71 stackmanage_35.scala 904:31]
  wire [31:0] _GEN_234 = LUT_stack_io_push_14 & _T_1 ? $signed(32'sh0) : $signed(_GEN_212); // @[stackmanage_35.scala 887:71 stackmanage_35.scala 905:31]
  wire [31:0] _GEN_235 = LUT_stack_io_push_14 & _T_1 ? $signed(32'sh0) : $signed(_GEN_213); // @[stackmanage_35.scala 887:71 stackmanage_35.scala 906:31]
  wire [31:0] _GEN_236 = LUT_stack_io_push_14 & _T_1 ? $signed(32'sh0) : $signed(_GEN_214); // @[stackmanage_35.scala 887:71 stackmanage_35.scala 907:31]
  wire [31:0] _GEN_237 = LUT_stack_io_push_14 & _T_1 ? $signed(32'sh0) : $signed(_GEN_215); // @[stackmanage_35.scala 887:71 stackmanage_35.scala 908:31]
  wire [31:0] _GEN_238 = LUT_stack_io_push_14 & _T_1 ? $signed(32'sh0) : $signed(_GEN_216); // @[stackmanage_35.scala 887:71 stackmanage_35.scala 909:31]
  wire [31:0] _GEN_239 = LUT_stack_io_push_14 & _T_1 ? $signed(32'sh0) : $signed(_GEN_217); // @[stackmanage_35.scala 887:71 stackmanage_35.scala 910:31]
  wire [31:0] _GEN_240 = LUT_stack_io_push_14 & _T_1 ? $signed(32'sh0) : $signed(_GEN_218); // @[stackmanage_35.scala 887:71 stackmanage_35.scala 911:31]
  wire [31:0] _GEN_241 = LUT_stack_io_push_14 & _T_1 ? $signed(32'sh0) : $signed(_GEN_219); // @[stackmanage_35.scala 887:71 stackmanage_35.scala 912:31]
  wire [31:0] _GEN_242 = LUT_stack_io_push_14 & _T_1 ? $signed(32'sh0) : $signed(_GEN_220); // @[stackmanage_35.scala 887:71 stackmanage_35.scala 913:31]
  wire [31:0] _GEN_243 = LUT_stack_io_push_14 & _T_1 ? $signed(32'sh0) : $signed(_GEN_221); // @[stackmanage_35.scala 887:71 stackmanage_35.scala 914:31]
  wire [31:0] _GEN_244 = LUT_stack_io_push_14 & _T_1 ? $signed(32'sh0) : $signed(_GEN_222); // @[stackmanage_35.scala 887:71 stackmanage_35.scala 915:31]
  wire [31:0] _GEN_245 = LUT_stack_io_push_14 & _T_1 ? $signed(32'sh0) : $signed(_GEN_223); // @[stackmanage_35.scala 887:71 stackmanage_35.scala 916:31]
  wire [31:0] _GEN_246 = LUT_stack_io_push_14 & _T_1 ? $signed(32'sh0) : $signed(_GEN_224); // @[stackmanage_35.scala 887:71 stackmanage_35.scala 917:31]
  wire [31:0] _GEN_247 = LUT_stack_io_push_14 & _T_1 ? $signed(32'sh0) : $signed(_GEN_225); // @[stackmanage_35.scala 887:71 stackmanage_35.scala 918:31]
  wire [31:0] _GEN_248 = LUT_stack_io_push_14 & _T_1 ? $signed(32'sh0) : $signed(_GEN_226); // @[stackmanage_35.scala 887:71 stackmanage_35.scala 919:31]
  wire [31:0] _GEN_249 = LUT_stack_io_push_14 & _T_1 ? $signed(32'sh0) : $signed(_GEN_227); // @[stackmanage_35.scala 887:71 stackmanage_35.scala 920:31]
  wire [31:0] _GEN_250 = LUT_stack_io_push_14 & _T_1 ? $signed(32'sh0) : $signed(_GEN_228); // @[stackmanage_35.scala 887:71 stackmanage_35.scala 921:31]
  wire [31:0] _GEN_251 = LUT_stack_io_push_14 & _T_1 ? $signed(32'sh0) : $signed(_GEN_229); // @[stackmanage_35.scala 887:71 stackmanage_35.scala 922:31]
  wire [31:0] _GEN_252 = LUT_stack_io_push_13 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 851:71 stackmanage_35.scala 852:30]
  wire [31:0] _GEN_254 = LUT_stack_io_push_13 & _T_1 ? $signed(32'sh0) : $signed(_GEN_230); // @[stackmanage_35.scala 851:71 stackmanage_35.scala 866:31]
  wire [31:0] _GEN_255 = LUT_stack_io_push_13 & _T_1 ? $signed(32'sh0) : $signed(_GEN_232); // @[stackmanage_35.scala 851:71 stackmanage_35.scala 867:31]
  wire [31:0] _GEN_256 = LUT_stack_io_push_13 & _T_1 ? $signed(32'sh0) : $signed(_GEN_233); // @[stackmanage_35.scala 851:71 stackmanage_35.scala 868:31]
  wire [31:0] _GEN_257 = LUT_stack_io_push_13 & _T_1 ? $signed(32'sh0) : $signed(_GEN_234); // @[stackmanage_35.scala 851:71 stackmanage_35.scala 869:31]
  wire [31:0] _GEN_258 = LUT_stack_io_push_13 & _T_1 ? $signed(32'sh0) : $signed(_GEN_235); // @[stackmanage_35.scala 851:71 stackmanage_35.scala 870:31]
  wire [31:0] _GEN_259 = LUT_stack_io_push_13 & _T_1 ? $signed(32'sh0) : $signed(_GEN_236); // @[stackmanage_35.scala 851:71 stackmanage_35.scala 871:31]
  wire [31:0] _GEN_260 = LUT_stack_io_push_13 & _T_1 ? $signed(32'sh0) : $signed(_GEN_237); // @[stackmanage_35.scala 851:71 stackmanage_35.scala 872:31]
  wire [31:0] _GEN_261 = LUT_stack_io_push_13 & _T_1 ? $signed(32'sh0) : $signed(_GEN_238); // @[stackmanage_35.scala 851:71 stackmanage_35.scala 873:31]
  wire [31:0] _GEN_262 = LUT_stack_io_push_13 & _T_1 ? $signed(32'sh0) : $signed(_GEN_239); // @[stackmanage_35.scala 851:71 stackmanage_35.scala 874:31]
  wire [31:0] _GEN_263 = LUT_stack_io_push_13 & _T_1 ? $signed(32'sh0) : $signed(_GEN_240); // @[stackmanage_35.scala 851:71 stackmanage_35.scala 875:31]
  wire [31:0] _GEN_264 = LUT_stack_io_push_13 & _T_1 ? $signed(32'sh0) : $signed(_GEN_241); // @[stackmanage_35.scala 851:71 stackmanage_35.scala 876:31]
  wire [31:0] _GEN_265 = LUT_stack_io_push_13 & _T_1 ? $signed(32'sh0) : $signed(_GEN_242); // @[stackmanage_35.scala 851:71 stackmanage_35.scala 877:31]
  wire [31:0] _GEN_266 = LUT_stack_io_push_13 & _T_1 ? $signed(32'sh0) : $signed(_GEN_243); // @[stackmanage_35.scala 851:71 stackmanage_35.scala 878:31]
  wire [31:0] _GEN_267 = LUT_stack_io_push_13 & _T_1 ? $signed(32'sh0) : $signed(_GEN_244); // @[stackmanage_35.scala 851:71 stackmanage_35.scala 879:31]
  wire [31:0] _GEN_268 = LUT_stack_io_push_13 & _T_1 ? $signed(32'sh0) : $signed(_GEN_245); // @[stackmanage_35.scala 851:71 stackmanage_35.scala 880:31]
  wire [31:0] _GEN_269 = LUT_stack_io_push_13 & _T_1 ? $signed(32'sh0) : $signed(_GEN_246); // @[stackmanage_35.scala 851:71 stackmanage_35.scala 881:31]
  wire [31:0] _GEN_270 = LUT_stack_io_push_13 & _T_1 ? $signed(32'sh0) : $signed(_GEN_247); // @[stackmanage_35.scala 851:71 stackmanage_35.scala 882:31]
  wire [31:0] _GEN_271 = LUT_stack_io_push_13 & _T_1 ? $signed(32'sh0) : $signed(_GEN_248); // @[stackmanage_35.scala 851:71 stackmanage_35.scala 883:31]
  wire [31:0] _GEN_272 = LUT_stack_io_push_13 & _T_1 ? $signed(32'sh0) : $signed(_GEN_249); // @[stackmanage_35.scala 851:71 stackmanage_35.scala 884:31]
  wire [31:0] _GEN_273 = LUT_stack_io_push_13 & _T_1 ? $signed(32'sh0) : $signed(_GEN_250); // @[stackmanage_35.scala 851:71 stackmanage_35.scala 885:31]
  wire [31:0] _GEN_274 = LUT_stack_io_push_13 & _T_1 ? $signed(32'sh0) : $signed(_GEN_251); // @[stackmanage_35.scala 851:71 stackmanage_35.scala 886:31]
  wire [31:0] _GEN_275 = LUT_stack_io_push_12 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 815:71 stackmanage_35.scala 816:30]
  wire [31:0] _GEN_277 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_252); // @[stackmanage_35.scala 815:71 stackmanage_35.scala 829:31]
  wire [31:0] _GEN_278 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_254); // @[stackmanage_35.scala 815:71 stackmanage_35.scala 830:31]
  wire [31:0] _GEN_279 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_255); // @[stackmanage_35.scala 815:71 stackmanage_35.scala 831:31]
  wire [31:0] _GEN_280 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_256); // @[stackmanage_35.scala 815:71 stackmanage_35.scala 832:31]
  wire [31:0] _GEN_281 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_257); // @[stackmanage_35.scala 815:71 stackmanage_35.scala 833:31]
  wire [31:0] _GEN_282 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_258); // @[stackmanage_35.scala 815:71 stackmanage_35.scala 834:31]
  wire [31:0] _GEN_283 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_259); // @[stackmanage_35.scala 815:71 stackmanage_35.scala 835:31]
  wire [31:0] _GEN_284 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_260); // @[stackmanage_35.scala 815:71 stackmanage_35.scala 836:31]
  wire [31:0] _GEN_285 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_261); // @[stackmanage_35.scala 815:71 stackmanage_35.scala 837:31]
  wire [31:0] _GEN_286 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_262); // @[stackmanage_35.scala 815:71 stackmanage_35.scala 838:31]
  wire [31:0] _GEN_287 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_263); // @[stackmanage_35.scala 815:71 stackmanage_35.scala 839:31]
  wire [31:0] _GEN_288 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_264); // @[stackmanage_35.scala 815:71 stackmanage_35.scala 840:31]
  wire [31:0] _GEN_289 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_265); // @[stackmanage_35.scala 815:71 stackmanage_35.scala 841:31]
  wire [31:0] _GEN_290 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_266); // @[stackmanage_35.scala 815:71 stackmanage_35.scala 842:31]
  wire [31:0] _GEN_291 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_267); // @[stackmanage_35.scala 815:71 stackmanage_35.scala 843:31]
  wire [31:0] _GEN_292 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_268); // @[stackmanage_35.scala 815:71 stackmanage_35.scala 844:31]
  wire [31:0] _GEN_293 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_269); // @[stackmanage_35.scala 815:71 stackmanage_35.scala 845:31]
  wire [31:0] _GEN_294 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_270); // @[stackmanage_35.scala 815:71 stackmanage_35.scala 846:31]
  wire [31:0] _GEN_295 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_271); // @[stackmanage_35.scala 815:71 stackmanage_35.scala 847:31]
  wire [31:0] _GEN_296 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_272); // @[stackmanage_35.scala 815:71 stackmanage_35.scala 848:31]
  wire [31:0] _GEN_297 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_273); // @[stackmanage_35.scala 815:71 stackmanage_35.scala 849:31]
  wire [31:0] _GEN_298 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_274); // @[stackmanage_35.scala 815:71 stackmanage_35.scala 850:31]
  wire [31:0] _GEN_299 = LUT_stack_io_push_11 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 779:71 stackmanage_35.scala 780:30]
  wire [31:0] _GEN_301 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_275); // @[stackmanage_35.scala 779:71 stackmanage_35.scala 792:31]
  wire [31:0] _GEN_302 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_277); // @[stackmanage_35.scala 779:71 stackmanage_35.scala 793:31]
  wire [31:0] _GEN_303 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_278); // @[stackmanage_35.scala 779:71 stackmanage_35.scala 794:31]
  wire [31:0] _GEN_304 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_279); // @[stackmanage_35.scala 779:71 stackmanage_35.scala 795:31]
  wire [31:0] _GEN_305 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_280); // @[stackmanage_35.scala 779:71 stackmanage_35.scala 796:31]
  wire [31:0] _GEN_306 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_281); // @[stackmanage_35.scala 779:71 stackmanage_35.scala 797:31]
  wire [31:0] _GEN_307 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_282); // @[stackmanage_35.scala 779:71 stackmanage_35.scala 798:31]
  wire [31:0] _GEN_308 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_283); // @[stackmanage_35.scala 779:71 stackmanage_35.scala 799:31]
  wire [31:0] _GEN_309 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_284); // @[stackmanage_35.scala 779:71 stackmanage_35.scala 800:31]
  wire [31:0] _GEN_310 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_285); // @[stackmanage_35.scala 779:71 stackmanage_35.scala 801:31]
  wire [31:0] _GEN_311 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_286); // @[stackmanage_35.scala 779:71 stackmanage_35.scala 802:31]
  wire [31:0] _GEN_312 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_287); // @[stackmanage_35.scala 779:71 stackmanage_35.scala 803:31]
  wire [31:0] _GEN_313 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_288); // @[stackmanage_35.scala 779:71 stackmanage_35.scala 804:31]
  wire [31:0] _GEN_314 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_289); // @[stackmanage_35.scala 779:71 stackmanage_35.scala 805:31]
  wire [31:0] _GEN_315 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_290); // @[stackmanage_35.scala 779:71 stackmanage_35.scala 806:31]
  wire [31:0] _GEN_316 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_291); // @[stackmanage_35.scala 779:71 stackmanage_35.scala 807:31]
  wire [31:0] _GEN_317 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_292); // @[stackmanage_35.scala 779:71 stackmanage_35.scala 808:31]
  wire [31:0] _GEN_318 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_293); // @[stackmanage_35.scala 779:71 stackmanage_35.scala 809:31]
  wire [31:0] _GEN_319 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_294); // @[stackmanage_35.scala 779:71 stackmanage_35.scala 810:31]
  wire [31:0] _GEN_320 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_295); // @[stackmanage_35.scala 779:71 stackmanage_35.scala 811:31]
  wire [31:0] _GEN_321 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_296); // @[stackmanage_35.scala 779:71 stackmanage_35.scala 812:31]
  wire [31:0] _GEN_322 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_297); // @[stackmanage_35.scala 779:71 stackmanage_35.scala 813:31]
  wire [31:0] _GEN_323 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_298); // @[stackmanage_35.scala 779:71 stackmanage_35.scala 814:31]
  wire [31:0] _GEN_324 = LUT_stack_io_push_10 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 743:71 stackmanage_35.scala 744:30]
  wire [31:0] _GEN_326 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_299); // @[stackmanage_35.scala 743:71 stackmanage_35.scala 755:31]
  wire [31:0] _GEN_327 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_301); // @[stackmanage_35.scala 743:71 stackmanage_35.scala 756:31]
  wire [31:0] _GEN_328 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_302); // @[stackmanage_35.scala 743:71 stackmanage_35.scala 757:31]
  wire [31:0] _GEN_329 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_303); // @[stackmanage_35.scala 743:71 stackmanage_35.scala 758:31]
  wire [31:0] _GEN_330 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_304); // @[stackmanage_35.scala 743:71 stackmanage_35.scala 759:31]
  wire [31:0] _GEN_331 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_305); // @[stackmanage_35.scala 743:71 stackmanage_35.scala 760:31]
  wire [31:0] _GEN_332 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_306); // @[stackmanage_35.scala 743:71 stackmanage_35.scala 761:31]
  wire [31:0] _GEN_333 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_307); // @[stackmanage_35.scala 743:71 stackmanage_35.scala 762:31]
  wire [31:0] _GEN_334 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_308); // @[stackmanage_35.scala 743:71 stackmanage_35.scala 763:31]
  wire [31:0] _GEN_335 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_309); // @[stackmanage_35.scala 743:71 stackmanage_35.scala 764:31]
  wire [31:0] _GEN_336 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_310); // @[stackmanage_35.scala 743:71 stackmanage_35.scala 765:31]
  wire [31:0] _GEN_337 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_311); // @[stackmanage_35.scala 743:71 stackmanage_35.scala 766:31]
  wire [31:0] _GEN_338 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_312); // @[stackmanage_35.scala 743:71 stackmanage_35.scala 767:31]
  wire [31:0] _GEN_339 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_313); // @[stackmanage_35.scala 743:71 stackmanage_35.scala 768:31]
  wire [31:0] _GEN_340 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_314); // @[stackmanage_35.scala 743:71 stackmanage_35.scala 769:31]
  wire [31:0] _GEN_341 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_315); // @[stackmanage_35.scala 743:71 stackmanage_35.scala 770:31]
  wire [31:0] _GEN_342 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_316); // @[stackmanage_35.scala 743:71 stackmanage_35.scala 771:31]
  wire [31:0] _GEN_343 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_317); // @[stackmanage_35.scala 743:71 stackmanage_35.scala 772:31]
  wire [31:0] _GEN_344 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_318); // @[stackmanage_35.scala 743:71 stackmanage_35.scala 773:31]
  wire [31:0] _GEN_345 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_319); // @[stackmanage_35.scala 743:71 stackmanage_35.scala 774:31]
  wire [31:0] _GEN_346 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_320); // @[stackmanage_35.scala 743:71 stackmanage_35.scala 775:31]
  wire [31:0] _GEN_347 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_321); // @[stackmanage_35.scala 743:71 stackmanage_35.scala 776:31]
  wire [31:0] _GEN_348 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_322); // @[stackmanage_35.scala 743:71 stackmanage_35.scala 777:31]
  wire [31:0] _GEN_349 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_323); // @[stackmanage_35.scala 743:71 stackmanage_35.scala 778:31]
  wire [31:0] _GEN_350 = LUT_stack_io_push_9 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 707:70 stackmanage_35.scala 708:29]
  wire [31:0] _GEN_352 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_324); // @[stackmanage_35.scala 707:70 stackmanage_35.scala 718:31]
  wire [31:0] _GEN_353 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_326); // @[stackmanage_35.scala 707:70 stackmanage_35.scala 719:31]
  wire [31:0] _GEN_354 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_327); // @[stackmanage_35.scala 707:70 stackmanage_35.scala 720:31]
  wire [31:0] _GEN_355 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_328); // @[stackmanage_35.scala 707:70 stackmanage_35.scala 721:31]
  wire [31:0] _GEN_356 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_329); // @[stackmanage_35.scala 707:70 stackmanage_35.scala 722:31]
  wire [31:0] _GEN_357 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_330); // @[stackmanage_35.scala 707:70 stackmanage_35.scala 723:31]
  wire [31:0] _GEN_358 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_331); // @[stackmanage_35.scala 707:70 stackmanage_35.scala 724:31]
  wire [31:0] _GEN_359 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_332); // @[stackmanage_35.scala 707:70 stackmanage_35.scala 725:31]
  wire [31:0] _GEN_360 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_333); // @[stackmanage_35.scala 707:70 stackmanage_35.scala 726:31]
  wire [31:0] _GEN_361 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_334); // @[stackmanage_35.scala 707:70 stackmanage_35.scala 727:31]
  wire [31:0] _GEN_362 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_335); // @[stackmanage_35.scala 707:70 stackmanage_35.scala 728:31]
  wire [31:0] _GEN_363 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_336); // @[stackmanage_35.scala 707:70 stackmanage_35.scala 729:31]
  wire [31:0] _GEN_364 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_337); // @[stackmanage_35.scala 707:70 stackmanage_35.scala 730:31]
  wire [31:0] _GEN_365 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_338); // @[stackmanage_35.scala 707:70 stackmanage_35.scala 731:31]
  wire [31:0] _GEN_366 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_339); // @[stackmanage_35.scala 707:70 stackmanage_35.scala 732:31]
  wire [31:0] _GEN_367 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_340); // @[stackmanage_35.scala 707:70 stackmanage_35.scala 733:31]
  wire [31:0] _GEN_368 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_341); // @[stackmanage_35.scala 707:70 stackmanage_35.scala 734:31]
  wire [31:0] _GEN_369 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_342); // @[stackmanage_35.scala 707:70 stackmanage_35.scala 735:31]
  wire [31:0] _GEN_370 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_343); // @[stackmanage_35.scala 707:70 stackmanage_35.scala 736:31]
  wire [31:0] _GEN_371 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_344); // @[stackmanage_35.scala 707:70 stackmanage_35.scala 737:31]
  wire [31:0] _GEN_372 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_345); // @[stackmanage_35.scala 707:70 stackmanage_35.scala 738:31]
  wire [31:0] _GEN_373 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_346); // @[stackmanage_35.scala 707:70 stackmanage_35.scala 739:31]
  wire [31:0] _GEN_374 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_347); // @[stackmanage_35.scala 707:70 stackmanage_35.scala 740:31]
  wire [31:0] _GEN_375 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_348); // @[stackmanage_35.scala 707:70 stackmanage_35.scala 741:31]
  wire [31:0] _GEN_376 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_349); // @[stackmanage_35.scala 707:70 stackmanage_35.scala 742:31]
  wire [31:0] _GEN_377 = LUT_stack_io_push_8 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 671:70 stackmanage_35.scala 672:29]
  wire [31:0] _GEN_379 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_350); // @[stackmanage_35.scala 671:70 stackmanage_35.scala 681:30]
  wire [31:0] _GEN_380 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_352); // @[stackmanage_35.scala 671:70 stackmanage_35.scala 682:31]
  wire [31:0] _GEN_381 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_353); // @[stackmanage_35.scala 671:70 stackmanage_35.scala 683:31]
  wire [31:0] _GEN_382 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_354); // @[stackmanage_35.scala 671:70 stackmanage_35.scala 684:31]
  wire [31:0] _GEN_383 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_355); // @[stackmanage_35.scala 671:70 stackmanage_35.scala 685:31]
  wire [31:0] _GEN_384 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_356); // @[stackmanage_35.scala 671:70 stackmanage_35.scala 686:31]
  wire [31:0] _GEN_385 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_357); // @[stackmanage_35.scala 671:70 stackmanage_35.scala 687:31]
  wire [31:0] _GEN_386 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_358); // @[stackmanage_35.scala 671:70 stackmanage_35.scala 688:31]
  wire [31:0] _GEN_387 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_359); // @[stackmanage_35.scala 671:70 stackmanage_35.scala 689:31]
  wire [31:0] _GEN_388 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_360); // @[stackmanage_35.scala 671:70 stackmanage_35.scala 690:31]
  wire [31:0] _GEN_389 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_361); // @[stackmanage_35.scala 671:70 stackmanage_35.scala 691:31]
  wire [31:0] _GEN_390 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_362); // @[stackmanage_35.scala 671:70 stackmanage_35.scala 692:31]
  wire [31:0] _GEN_391 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_363); // @[stackmanage_35.scala 671:70 stackmanage_35.scala 693:31]
  wire [31:0] _GEN_392 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_364); // @[stackmanage_35.scala 671:70 stackmanage_35.scala 694:31]
  wire [31:0] _GEN_393 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_365); // @[stackmanage_35.scala 671:70 stackmanage_35.scala 695:31]
  wire [31:0] _GEN_394 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_366); // @[stackmanage_35.scala 671:70 stackmanage_35.scala 696:31]
  wire [31:0] _GEN_395 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_367); // @[stackmanage_35.scala 671:70 stackmanage_35.scala 697:31]
  wire [31:0] _GEN_396 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_368); // @[stackmanage_35.scala 671:70 stackmanage_35.scala 698:31]
  wire [31:0] _GEN_397 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_369); // @[stackmanage_35.scala 671:70 stackmanage_35.scala 699:31]
  wire [31:0] _GEN_398 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_370); // @[stackmanage_35.scala 671:70 stackmanage_35.scala 700:31]
  wire [31:0] _GEN_399 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_371); // @[stackmanage_35.scala 671:70 stackmanage_35.scala 701:31]
  wire [31:0] _GEN_400 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_372); // @[stackmanage_35.scala 671:70 stackmanage_35.scala 702:31]
  wire [31:0] _GEN_401 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_373); // @[stackmanage_35.scala 671:70 stackmanage_35.scala 703:31]
  wire [31:0] _GEN_402 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_374); // @[stackmanage_35.scala 671:70 stackmanage_35.scala 704:31]
  wire [31:0] _GEN_403 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_375); // @[stackmanage_35.scala 671:70 stackmanage_35.scala 705:31]
  wire [31:0] _GEN_404 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_376); // @[stackmanage_35.scala 671:70 stackmanage_35.scala 706:31]
  wire [31:0] _GEN_405 = LUT_stack_io_push_7 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 635:70 stackmanage_35.scala 636:29]
  wire [31:0] _GEN_407 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_377); // @[stackmanage_35.scala 635:70 stackmanage_35.scala 644:30]
  wire [31:0] _GEN_408 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_379); // @[stackmanage_35.scala 635:70 stackmanage_35.scala 645:30]
  wire [31:0] _GEN_409 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_380); // @[stackmanage_35.scala 635:70 stackmanage_35.scala 646:31]
  wire [31:0] _GEN_410 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_381); // @[stackmanage_35.scala 635:70 stackmanage_35.scala 647:31]
  wire [31:0] _GEN_411 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_382); // @[stackmanage_35.scala 635:70 stackmanage_35.scala 648:31]
  wire [31:0] _GEN_412 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_383); // @[stackmanage_35.scala 635:70 stackmanage_35.scala 649:31]
  wire [31:0] _GEN_413 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_384); // @[stackmanage_35.scala 635:70 stackmanage_35.scala 650:31]
  wire [31:0] _GEN_414 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_385); // @[stackmanage_35.scala 635:70 stackmanage_35.scala 651:31]
  wire [31:0] _GEN_415 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_386); // @[stackmanage_35.scala 635:70 stackmanage_35.scala 652:31]
  wire [31:0] _GEN_416 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_387); // @[stackmanage_35.scala 635:70 stackmanage_35.scala 653:31]
  wire [31:0] _GEN_417 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_388); // @[stackmanage_35.scala 635:70 stackmanage_35.scala 654:31]
  wire [31:0] _GEN_418 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_389); // @[stackmanage_35.scala 635:70 stackmanage_35.scala 655:31]
  wire [31:0] _GEN_419 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_390); // @[stackmanage_35.scala 635:70 stackmanage_35.scala 656:31]
  wire [31:0] _GEN_420 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_391); // @[stackmanage_35.scala 635:70 stackmanage_35.scala 657:31]
  wire [31:0] _GEN_421 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_392); // @[stackmanage_35.scala 635:70 stackmanage_35.scala 658:31]
  wire [31:0] _GEN_422 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_393); // @[stackmanage_35.scala 635:70 stackmanage_35.scala 659:31]
  wire [31:0] _GEN_423 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_394); // @[stackmanage_35.scala 635:70 stackmanage_35.scala 660:31]
  wire [31:0] _GEN_424 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_395); // @[stackmanage_35.scala 635:70 stackmanage_35.scala 661:31]
  wire [31:0] _GEN_425 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_396); // @[stackmanage_35.scala 635:70 stackmanage_35.scala 662:31]
  wire [31:0] _GEN_426 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_397); // @[stackmanage_35.scala 635:70 stackmanage_35.scala 663:31]
  wire [31:0] _GEN_427 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_398); // @[stackmanage_35.scala 635:70 stackmanage_35.scala 664:31]
  wire [31:0] _GEN_428 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_399); // @[stackmanage_35.scala 635:70 stackmanage_35.scala 665:31]
  wire [31:0] _GEN_429 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_400); // @[stackmanage_35.scala 635:70 stackmanage_35.scala 666:31]
  wire [31:0] _GEN_430 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_401); // @[stackmanage_35.scala 635:70 stackmanage_35.scala 667:31]
  wire [31:0] _GEN_431 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_402); // @[stackmanage_35.scala 635:70 stackmanage_35.scala 668:31]
  wire [31:0] _GEN_432 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_403); // @[stackmanage_35.scala 635:70 stackmanage_35.scala 669:31]
  wire [31:0] _GEN_433 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_404); // @[stackmanage_35.scala 635:70 stackmanage_35.scala 670:31]
  wire [31:0] _GEN_434 = LUT_stack_io_push_6 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 599:70 stackmanage_35.scala 600:29]
  wire [31:0] _GEN_436 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_405); // @[stackmanage_35.scala 599:70 stackmanage_35.scala 607:30]
  wire [31:0] _GEN_437 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_407); // @[stackmanage_35.scala 599:70 stackmanage_35.scala 608:30]
  wire [31:0] _GEN_438 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_408); // @[stackmanage_35.scala 599:70 stackmanage_35.scala 609:30]
  wire [31:0] _GEN_439 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_409); // @[stackmanage_35.scala 599:70 stackmanage_35.scala 610:31]
  wire [31:0] _GEN_440 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_410); // @[stackmanage_35.scala 599:70 stackmanage_35.scala 611:31]
  wire [31:0] _GEN_441 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_411); // @[stackmanage_35.scala 599:70 stackmanage_35.scala 612:31]
  wire [31:0] _GEN_442 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_412); // @[stackmanage_35.scala 599:70 stackmanage_35.scala 613:31]
  wire [31:0] _GEN_443 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_413); // @[stackmanage_35.scala 599:70 stackmanage_35.scala 614:31]
  wire [31:0] _GEN_444 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_414); // @[stackmanage_35.scala 599:70 stackmanage_35.scala 615:31]
  wire [31:0] _GEN_445 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_415); // @[stackmanage_35.scala 599:70 stackmanage_35.scala 616:31]
  wire [31:0] _GEN_446 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_416); // @[stackmanage_35.scala 599:70 stackmanage_35.scala 617:31]
  wire [31:0] _GEN_447 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_417); // @[stackmanage_35.scala 599:70 stackmanage_35.scala 618:31]
  wire [31:0] _GEN_448 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_418); // @[stackmanage_35.scala 599:70 stackmanage_35.scala 619:31]
  wire [31:0] _GEN_449 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_419); // @[stackmanage_35.scala 599:70 stackmanage_35.scala 620:31]
  wire [31:0] _GEN_450 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_420); // @[stackmanage_35.scala 599:70 stackmanage_35.scala 621:31]
  wire [31:0] _GEN_451 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_421); // @[stackmanage_35.scala 599:70 stackmanage_35.scala 622:31]
  wire [31:0] _GEN_452 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_422); // @[stackmanage_35.scala 599:70 stackmanage_35.scala 623:31]
  wire [31:0] _GEN_453 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_423); // @[stackmanage_35.scala 599:70 stackmanage_35.scala 624:31]
  wire [31:0] _GEN_454 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_424); // @[stackmanage_35.scala 599:70 stackmanage_35.scala 625:31]
  wire [31:0] _GEN_455 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_425); // @[stackmanage_35.scala 599:70 stackmanage_35.scala 626:31]
  wire [31:0] _GEN_456 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_426); // @[stackmanage_35.scala 599:70 stackmanage_35.scala 627:31]
  wire [31:0] _GEN_457 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_427); // @[stackmanage_35.scala 599:70 stackmanage_35.scala 628:31]
  wire [31:0] _GEN_458 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_428); // @[stackmanage_35.scala 599:70 stackmanage_35.scala 629:31]
  wire [31:0] _GEN_459 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_429); // @[stackmanage_35.scala 599:70 stackmanage_35.scala 630:31]
  wire [31:0] _GEN_460 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_430); // @[stackmanage_35.scala 599:70 stackmanage_35.scala 631:31]
  wire [31:0] _GEN_461 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_431); // @[stackmanage_35.scala 599:70 stackmanage_35.scala 632:31]
  wire [31:0] _GEN_462 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_432); // @[stackmanage_35.scala 599:70 stackmanage_35.scala 633:31]
  wire [31:0] _GEN_463 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_433); // @[stackmanage_35.scala 599:70 stackmanage_35.scala 634:31]
  wire [31:0] _GEN_464 = LUT_stack_io_push_5 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 563:70 stackmanage_35.scala 564:29]
  wire [31:0] _GEN_466 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_434); // @[stackmanage_35.scala 563:70 stackmanage_35.scala 570:30]
  wire [31:0] _GEN_467 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_436); // @[stackmanage_35.scala 563:70 stackmanage_35.scala 571:30]
  wire [31:0] _GEN_468 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_437); // @[stackmanage_35.scala 563:70 stackmanage_35.scala 572:30]
  wire [31:0] _GEN_469 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_438); // @[stackmanage_35.scala 563:70 stackmanage_35.scala 573:30]
  wire [31:0] _GEN_470 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_439); // @[stackmanage_35.scala 563:70 stackmanage_35.scala 574:31]
  wire [31:0] _GEN_471 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_440); // @[stackmanage_35.scala 563:70 stackmanage_35.scala 575:31]
  wire [31:0] _GEN_472 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_441); // @[stackmanage_35.scala 563:70 stackmanage_35.scala 576:31]
  wire [31:0] _GEN_473 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_442); // @[stackmanage_35.scala 563:70 stackmanage_35.scala 577:31]
  wire [31:0] _GEN_474 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_443); // @[stackmanage_35.scala 563:70 stackmanage_35.scala 578:31]
  wire [31:0] _GEN_475 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_444); // @[stackmanage_35.scala 563:70 stackmanage_35.scala 579:31]
  wire [31:0] _GEN_476 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_445); // @[stackmanage_35.scala 563:70 stackmanage_35.scala 580:31]
  wire [31:0] _GEN_477 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_446); // @[stackmanage_35.scala 563:70 stackmanage_35.scala 581:31]
  wire [31:0] _GEN_478 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_447); // @[stackmanage_35.scala 563:70 stackmanage_35.scala 582:31]
  wire [31:0] _GEN_479 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_448); // @[stackmanage_35.scala 563:70 stackmanage_35.scala 583:31]
  wire [31:0] _GEN_480 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_449); // @[stackmanage_35.scala 563:70 stackmanage_35.scala 584:31]
  wire [31:0] _GEN_481 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_450); // @[stackmanage_35.scala 563:70 stackmanage_35.scala 585:31]
  wire [31:0] _GEN_482 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_451); // @[stackmanage_35.scala 563:70 stackmanage_35.scala 586:31]
  wire [31:0] _GEN_483 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_452); // @[stackmanage_35.scala 563:70 stackmanage_35.scala 587:31]
  wire [31:0] _GEN_484 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_453); // @[stackmanage_35.scala 563:70 stackmanage_35.scala 588:31]
  wire [31:0] _GEN_485 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_454); // @[stackmanage_35.scala 563:70 stackmanage_35.scala 589:31]
  wire [31:0] _GEN_486 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_455); // @[stackmanage_35.scala 563:70 stackmanage_35.scala 590:31]
  wire [31:0] _GEN_487 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_456); // @[stackmanage_35.scala 563:70 stackmanage_35.scala 591:31]
  wire [31:0] _GEN_488 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_457); // @[stackmanage_35.scala 563:70 stackmanage_35.scala 592:31]
  wire [31:0] _GEN_489 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_458); // @[stackmanage_35.scala 563:70 stackmanage_35.scala 593:31]
  wire [31:0] _GEN_490 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_459); // @[stackmanage_35.scala 563:70 stackmanage_35.scala 594:31]
  wire [31:0] _GEN_491 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_460); // @[stackmanage_35.scala 563:70 stackmanage_35.scala 595:31]
  wire [31:0] _GEN_492 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_461); // @[stackmanage_35.scala 563:70 stackmanage_35.scala 596:31]
  wire [31:0] _GEN_493 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_462); // @[stackmanage_35.scala 563:70 stackmanage_35.scala 597:31]
  wire [31:0] _GEN_494 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_463); // @[stackmanage_35.scala 563:70 stackmanage_35.scala 598:31]
  wire [31:0] _GEN_495 = LUT_stack_io_push_4 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 527:70 stackmanage_35.scala 528:29]
  wire [31:0] _GEN_497 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_464); // @[stackmanage_35.scala 527:70 stackmanage_35.scala 533:30]
  wire [31:0] _GEN_498 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_466); // @[stackmanage_35.scala 527:70 stackmanage_35.scala 534:30]
  wire [31:0] _GEN_499 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_467); // @[stackmanage_35.scala 527:70 stackmanage_35.scala 535:30]
  wire [31:0] _GEN_500 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_468); // @[stackmanage_35.scala 527:70 stackmanage_35.scala 536:30]
  wire [31:0] _GEN_501 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_469); // @[stackmanage_35.scala 527:70 stackmanage_35.scala 537:30]
  wire [31:0] _GEN_502 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_470); // @[stackmanage_35.scala 527:70 stackmanage_35.scala 538:31]
  wire [31:0] _GEN_503 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_471); // @[stackmanage_35.scala 527:70 stackmanage_35.scala 539:31]
  wire [31:0] _GEN_504 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_472); // @[stackmanage_35.scala 527:70 stackmanage_35.scala 540:31]
  wire [31:0] _GEN_505 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_473); // @[stackmanage_35.scala 527:70 stackmanage_35.scala 541:31]
  wire [31:0] _GEN_506 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_474); // @[stackmanage_35.scala 527:70 stackmanage_35.scala 542:31]
  wire [31:0] _GEN_507 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_475); // @[stackmanage_35.scala 527:70 stackmanage_35.scala 543:31]
  wire [31:0] _GEN_508 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_476); // @[stackmanage_35.scala 527:70 stackmanage_35.scala 544:31]
  wire [31:0] _GEN_509 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_477); // @[stackmanage_35.scala 527:70 stackmanage_35.scala 545:31]
  wire [31:0] _GEN_510 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_478); // @[stackmanage_35.scala 527:70 stackmanage_35.scala 546:31]
  wire [31:0] _GEN_511 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_479); // @[stackmanage_35.scala 527:70 stackmanage_35.scala 547:31]
  wire [31:0] _GEN_512 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_480); // @[stackmanage_35.scala 527:70 stackmanage_35.scala 548:31]
  wire [31:0] _GEN_513 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_481); // @[stackmanage_35.scala 527:70 stackmanage_35.scala 549:31]
  wire [31:0] _GEN_514 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_482); // @[stackmanage_35.scala 527:70 stackmanage_35.scala 550:31]
  wire [31:0] _GEN_515 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_483); // @[stackmanage_35.scala 527:70 stackmanage_35.scala 551:31]
  wire [31:0] _GEN_516 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_484); // @[stackmanage_35.scala 527:70 stackmanage_35.scala 552:31]
  wire [31:0] _GEN_517 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_485); // @[stackmanage_35.scala 527:70 stackmanage_35.scala 553:31]
  wire [31:0] _GEN_518 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_486); // @[stackmanage_35.scala 527:70 stackmanage_35.scala 554:31]
  wire [31:0] _GEN_519 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_487); // @[stackmanage_35.scala 527:70 stackmanage_35.scala 555:31]
  wire [31:0] _GEN_520 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_488); // @[stackmanage_35.scala 527:70 stackmanage_35.scala 556:31]
  wire [31:0] _GEN_521 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_489); // @[stackmanage_35.scala 527:70 stackmanage_35.scala 557:31]
  wire [31:0] _GEN_522 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_490); // @[stackmanage_35.scala 527:70 stackmanage_35.scala 558:31]
  wire [31:0] _GEN_523 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_491); // @[stackmanage_35.scala 527:70 stackmanage_35.scala 559:31]
  wire [31:0] _GEN_524 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_492); // @[stackmanage_35.scala 527:70 stackmanage_35.scala 560:31]
  wire [31:0] _GEN_525 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_493); // @[stackmanage_35.scala 527:70 stackmanage_35.scala 561:31]
  wire [31:0] _GEN_526 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_494); // @[stackmanage_35.scala 527:70 stackmanage_35.scala 562:31]
  wire [31:0] _GEN_527 = LUT_stack_io_push_3 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 491:70 stackmanage_35.scala 492:29]
  wire [31:0] _GEN_529 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_495); // @[stackmanage_35.scala 491:70 stackmanage_35.scala 496:30]
  wire [31:0] _GEN_530 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_497); // @[stackmanage_35.scala 491:70 stackmanage_35.scala 497:30]
  wire [31:0] _GEN_531 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_498); // @[stackmanage_35.scala 491:70 stackmanage_35.scala 498:30]
  wire [31:0] _GEN_532 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_499); // @[stackmanage_35.scala 491:70 stackmanage_35.scala 499:30]
  wire [31:0] _GEN_533 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_500); // @[stackmanage_35.scala 491:70 stackmanage_35.scala 500:30]
  wire [31:0] _GEN_534 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_501); // @[stackmanage_35.scala 491:70 stackmanage_35.scala 501:30]
  wire [31:0] _GEN_535 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_502); // @[stackmanage_35.scala 491:70 stackmanage_35.scala 502:31]
  wire [31:0] _GEN_536 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_503); // @[stackmanage_35.scala 491:70 stackmanage_35.scala 503:31]
  wire [31:0] _GEN_537 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_504); // @[stackmanage_35.scala 491:70 stackmanage_35.scala 504:31]
  wire [31:0] _GEN_538 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_505); // @[stackmanage_35.scala 491:70 stackmanage_35.scala 505:31]
  wire [31:0] _GEN_539 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_506); // @[stackmanage_35.scala 491:70 stackmanage_35.scala 506:31]
  wire [31:0] _GEN_540 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_507); // @[stackmanage_35.scala 491:70 stackmanage_35.scala 507:31]
  wire [31:0] _GEN_541 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_508); // @[stackmanage_35.scala 491:70 stackmanage_35.scala 508:31]
  wire [31:0] _GEN_542 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_509); // @[stackmanage_35.scala 491:70 stackmanage_35.scala 509:31]
  wire [31:0] _GEN_543 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_510); // @[stackmanage_35.scala 491:70 stackmanage_35.scala 510:31]
  wire [31:0] _GEN_544 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_511); // @[stackmanage_35.scala 491:70 stackmanage_35.scala 511:31]
  wire [31:0] _GEN_545 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_512); // @[stackmanage_35.scala 491:70 stackmanage_35.scala 512:31]
  wire [31:0] _GEN_546 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_513); // @[stackmanage_35.scala 491:70 stackmanage_35.scala 513:31]
  wire [31:0] _GEN_547 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_514); // @[stackmanage_35.scala 491:70 stackmanage_35.scala 514:31]
  wire [31:0] _GEN_548 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_515); // @[stackmanage_35.scala 491:70 stackmanage_35.scala 515:31]
  wire [31:0] _GEN_549 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_516); // @[stackmanage_35.scala 491:70 stackmanage_35.scala 516:31]
  wire [31:0] _GEN_550 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_517); // @[stackmanage_35.scala 491:70 stackmanage_35.scala 517:31]
  wire [31:0] _GEN_551 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_518); // @[stackmanage_35.scala 491:70 stackmanage_35.scala 518:31]
  wire [31:0] _GEN_552 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_519); // @[stackmanage_35.scala 491:70 stackmanage_35.scala 519:31]
  wire [31:0] _GEN_553 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_520); // @[stackmanage_35.scala 491:70 stackmanage_35.scala 520:31]
  wire [31:0] _GEN_554 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_521); // @[stackmanage_35.scala 491:70 stackmanage_35.scala 521:31]
  wire [31:0] _GEN_555 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_522); // @[stackmanage_35.scala 491:70 stackmanage_35.scala 522:31]
  wire [31:0] _GEN_556 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_523); // @[stackmanage_35.scala 491:70 stackmanage_35.scala 523:31]
  wire [31:0] _GEN_557 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_524); // @[stackmanage_35.scala 491:70 stackmanage_35.scala 524:31]
  wire [31:0] _GEN_558 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_525); // @[stackmanage_35.scala 491:70 stackmanage_35.scala 525:31]
  wire [31:0] _GEN_559 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_526); // @[stackmanage_35.scala 491:70 stackmanage_35.scala 526:31]
  wire [31:0] _GEN_560 = LUT_stack_io_push_2 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 455:70 stackmanage_35.scala 456:29]
  wire [31:0] _GEN_562 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_527); // @[stackmanage_35.scala 455:70 stackmanage_35.scala 459:30]
  wire [31:0] _GEN_563 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_529); // @[stackmanage_35.scala 455:70 stackmanage_35.scala 460:30]
  wire [31:0] _GEN_564 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_530); // @[stackmanage_35.scala 455:70 stackmanage_35.scala 461:30]
  wire [31:0] _GEN_565 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_531); // @[stackmanage_35.scala 455:70 stackmanage_35.scala 462:30]
  wire [31:0] _GEN_566 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_532); // @[stackmanage_35.scala 455:70 stackmanage_35.scala 463:30]
  wire [31:0] _GEN_567 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_533); // @[stackmanage_35.scala 455:70 stackmanage_35.scala 464:30]
  wire [31:0] _GEN_568 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_534); // @[stackmanage_35.scala 455:70 stackmanage_35.scala 465:30]
  wire [31:0] _GEN_569 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_535); // @[stackmanage_35.scala 455:70 stackmanage_35.scala 466:31]
  wire [31:0] _GEN_570 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_536); // @[stackmanage_35.scala 455:70 stackmanage_35.scala 467:31]
  wire [31:0] _GEN_571 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_537); // @[stackmanage_35.scala 455:70 stackmanage_35.scala 468:31]
  wire [31:0] _GEN_572 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_538); // @[stackmanage_35.scala 455:70 stackmanage_35.scala 469:31]
  wire [31:0] _GEN_573 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_539); // @[stackmanage_35.scala 455:70 stackmanage_35.scala 470:31]
  wire [31:0] _GEN_574 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_540); // @[stackmanage_35.scala 455:70 stackmanage_35.scala 471:31]
  wire [31:0] _GEN_575 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_541); // @[stackmanage_35.scala 455:70 stackmanage_35.scala 472:31]
  wire [31:0] _GEN_576 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_542); // @[stackmanage_35.scala 455:70 stackmanage_35.scala 473:31]
  wire [31:0] _GEN_577 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_543); // @[stackmanage_35.scala 455:70 stackmanage_35.scala 474:31]
  wire [31:0] _GEN_578 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_544); // @[stackmanage_35.scala 455:70 stackmanage_35.scala 475:31]
  wire [31:0] _GEN_579 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_545); // @[stackmanage_35.scala 455:70 stackmanage_35.scala 476:31]
  wire [31:0] _GEN_580 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_546); // @[stackmanage_35.scala 455:70 stackmanage_35.scala 477:31]
  wire [31:0] _GEN_581 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_547); // @[stackmanage_35.scala 455:70 stackmanage_35.scala 478:31]
  wire [31:0] _GEN_582 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_548); // @[stackmanage_35.scala 455:70 stackmanage_35.scala 479:31]
  wire [31:0] _GEN_583 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_549); // @[stackmanage_35.scala 455:70 stackmanage_35.scala 480:31]
  wire [31:0] _GEN_584 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_550); // @[stackmanage_35.scala 455:70 stackmanage_35.scala 481:31]
  wire [31:0] _GEN_585 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_551); // @[stackmanage_35.scala 455:70 stackmanage_35.scala 482:31]
  wire [31:0] _GEN_586 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_552); // @[stackmanage_35.scala 455:70 stackmanage_35.scala 483:31]
  wire [31:0] _GEN_587 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_553); // @[stackmanage_35.scala 455:70 stackmanage_35.scala 484:31]
  wire [31:0] _GEN_588 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_554); // @[stackmanage_35.scala 455:70 stackmanage_35.scala 485:31]
  wire [31:0] _GEN_589 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_555); // @[stackmanage_35.scala 455:70 stackmanage_35.scala 486:31]
  wire [31:0] _GEN_590 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_556); // @[stackmanage_35.scala 455:70 stackmanage_35.scala 487:31]
  wire [31:0] _GEN_591 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_557); // @[stackmanage_35.scala 455:70 stackmanage_35.scala 488:31]
  wire [31:0] _GEN_592 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_558); // @[stackmanage_35.scala 455:70 stackmanage_35.scala 489:31]
  wire [31:0] _GEN_593 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_559); // @[stackmanage_35.scala 455:70 stackmanage_35.scala 490:31]
  wire [31:0] _GEN_594 = LUT_stack_io_push_1 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 419:70 stackmanage_35.scala 420:29]
  wire [31:0] _GEN_596 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_560); // @[stackmanage_35.scala 419:70 stackmanage_35.scala 422:30]
  wire [31:0] _GEN_597 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_562); // @[stackmanage_35.scala 419:70 stackmanage_35.scala 423:30]
  wire [31:0] _GEN_598 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_563); // @[stackmanage_35.scala 419:70 stackmanage_35.scala 424:30]
  wire [31:0] _GEN_599 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_564); // @[stackmanage_35.scala 419:70 stackmanage_35.scala 425:30]
  wire [31:0] _GEN_600 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_565); // @[stackmanage_35.scala 419:70 stackmanage_35.scala 426:30]
  wire [31:0] _GEN_601 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_566); // @[stackmanage_35.scala 419:70 stackmanage_35.scala 427:30]
  wire [31:0] _GEN_602 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_567); // @[stackmanage_35.scala 419:70 stackmanage_35.scala 428:30]
  wire [31:0] _GEN_603 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_568); // @[stackmanage_35.scala 419:70 stackmanage_35.scala 429:30]
  wire [31:0] _GEN_604 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_569); // @[stackmanage_35.scala 419:70 stackmanage_35.scala 430:31]
  wire [31:0] _GEN_605 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_570); // @[stackmanage_35.scala 419:70 stackmanage_35.scala 431:31]
  wire [31:0] _GEN_606 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_571); // @[stackmanage_35.scala 419:70 stackmanage_35.scala 432:31]
  wire [31:0] _GEN_607 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_572); // @[stackmanage_35.scala 419:70 stackmanage_35.scala 433:31]
  wire [31:0] _GEN_608 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_573); // @[stackmanage_35.scala 419:70 stackmanage_35.scala 434:31]
  wire [31:0] _GEN_609 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_574); // @[stackmanage_35.scala 419:70 stackmanage_35.scala 435:31]
  wire [31:0] _GEN_610 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_575); // @[stackmanage_35.scala 419:70 stackmanage_35.scala 436:31]
  wire [31:0] _GEN_611 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_576); // @[stackmanage_35.scala 419:70 stackmanage_35.scala 437:31]
  wire [31:0] _GEN_612 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_577); // @[stackmanage_35.scala 419:70 stackmanage_35.scala 438:31]
  wire [31:0] _GEN_613 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_578); // @[stackmanage_35.scala 419:70 stackmanage_35.scala 439:31]
  wire [31:0] _GEN_614 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_579); // @[stackmanage_35.scala 419:70 stackmanage_35.scala 440:31]
  wire [31:0] _GEN_615 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_580); // @[stackmanage_35.scala 419:70 stackmanage_35.scala 441:31]
  wire [31:0] _GEN_616 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_581); // @[stackmanage_35.scala 419:70 stackmanage_35.scala 442:31]
  wire [31:0] _GEN_617 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_582); // @[stackmanage_35.scala 419:70 stackmanage_35.scala 443:31]
  wire [31:0] _GEN_618 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_583); // @[stackmanage_35.scala 419:70 stackmanage_35.scala 444:31]
  wire [31:0] _GEN_619 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_584); // @[stackmanage_35.scala 419:70 stackmanage_35.scala 445:31]
  wire [31:0] _GEN_620 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_585); // @[stackmanage_35.scala 419:70 stackmanage_35.scala 446:31]
  wire [31:0] _GEN_621 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_586); // @[stackmanage_35.scala 419:70 stackmanage_35.scala 447:31]
  wire [31:0] _GEN_622 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_587); // @[stackmanage_35.scala 419:70 stackmanage_35.scala 448:31]
  wire [31:0] _GEN_623 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_588); // @[stackmanage_35.scala 419:70 stackmanage_35.scala 449:31]
  wire [31:0] _GEN_624 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_589); // @[stackmanage_35.scala 419:70 stackmanage_35.scala 450:31]
  wire [31:0] _GEN_625 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_590); // @[stackmanage_35.scala 419:70 stackmanage_35.scala 451:31]
  wire [31:0] _GEN_626 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_591); // @[stackmanage_35.scala 419:70 stackmanage_35.scala 452:31]
  wire [31:0] _GEN_627 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_592); // @[stackmanage_35.scala 419:70 stackmanage_35.scala 453:31]
  wire [31:0] _GEN_628 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_593); // @[stackmanage_35.scala 419:70 stackmanage_35.scala 454:31]
  reg [31:0] hitT_out_temp; // @[stackmanage_35.scala 1682:34]
  reg [31:0] ray_out_temp; // @[stackmanage_35.scala 1683:35]
  reg [31:0] node_out_temp; // @[stackmanage_35.scala 1684:32]
  reg  pop_valid_1; // @[stackmanage_35.scala 1685:38]
  wire  _T_105 = LUT_stack_io_pop_en; // @[stackmanage_35.scala 1686:29]
  wire [31:0] _GEN_664 = _T_105 & LUT_stack_io_pop_34 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 4100:69 stackmanage_35.scala 4101:29 stackmanage_35.scala 4240:29]
  wire [31:0] _GEN_665 = _T_105 & LUT_stack_io_pop_34 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 4100:69 stackmanage_35.scala 4102:28 stackmanage_35.scala 4241:28]
  wire [31:0] _GEN_667 = _T_105 & LUT_stack_io_pop_33 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 4029:69 stackmanage_35.scala 4030:29]
  wire [31:0] _GEN_668 = _T_105 & LUT_stack_io_pop_33 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 4029:69 stackmanage_35.scala 4031:28]
  wire [31:0] _GEN_670 = _T_105 & LUT_stack_io_pop_33 ? 32'h0 : _GEN_664; // @[stackmanage_35.scala 4029:69 stackmanage_35.scala 4098:29]
  wire [31:0] _GEN_671 = _T_105 & LUT_stack_io_pop_33 ? 32'h0 : _GEN_665; // @[stackmanage_35.scala 4029:69 stackmanage_35.scala 4099:28]
  wire [31:0] _GEN_672 = _T_105 & LUT_stack_io_pop_32 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 3958:69 stackmanage_35.scala 3959:29]
  wire [31:0] _GEN_673 = _T_105 & LUT_stack_io_pop_32 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 3958:69 stackmanage_35.scala 3960:28]
  wire [31:0] _GEN_675 = _T_105 & LUT_stack_io_pop_32 ? 32'h0 : _GEN_667; // @[stackmanage_35.scala 3958:69 stackmanage_35.scala 4025:29]
  wire [31:0] _GEN_676 = _T_105 & LUT_stack_io_pop_32 ? 32'h0 : _GEN_668; // @[stackmanage_35.scala 3958:69 stackmanage_35.scala 4026:28]
  wire [31:0] _GEN_677 = _T_105 & LUT_stack_io_pop_32 ? 32'h0 : _GEN_670; // @[stackmanage_35.scala 3958:69 stackmanage_35.scala 4027:29]
  wire [31:0] _GEN_678 = _T_105 & LUT_stack_io_pop_32 ? 32'h0 : _GEN_671; // @[stackmanage_35.scala 3958:69 stackmanage_35.scala 4028:28]
  wire [31:0] _GEN_679 = _T_105 & LUT_stack_io_pop_31 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 3887:69 stackmanage_35.scala 3888:29]
  wire [31:0] _GEN_680 = _T_105 & LUT_stack_io_pop_31 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 3887:69 stackmanage_35.scala 3889:28]
  wire [31:0] _GEN_682 = _T_105 & LUT_stack_io_pop_31 ? 32'h0 : _GEN_672; // @[stackmanage_35.scala 3887:69 stackmanage_35.scala 3952:29]
  wire [31:0] _GEN_683 = _T_105 & LUT_stack_io_pop_31 ? 32'h0 : _GEN_673; // @[stackmanage_35.scala 3887:69 stackmanage_35.scala 3953:28]
  wire [31:0] _GEN_684 = _T_105 & LUT_stack_io_pop_31 ? 32'h0 : _GEN_675; // @[stackmanage_35.scala 3887:69 stackmanage_35.scala 3954:29]
  wire [31:0] _GEN_685 = _T_105 & LUT_stack_io_pop_31 ? 32'h0 : _GEN_676; // @[stackmanage_35.scala 3887:69 stackmanage_35.scala 3955:28]
  wire [31:0] _GEN_686 = _T_105 & LUT_stack_io_pop_31 ? 32'h0 : _GEN_677; // @[stackmanage_35.scala 3887:69 stackmanage_35.scala 3956:29]
  wire [31:0] _GEN_687 = _T_105 & LUT_stack_io_pop_31 ? 32'h0 : _GEN_678; // @[stackmanage_35.scala 3887:69 stackmanage_35.scala 3957:28]
  wire [31:0] _GEN_688 = _T_105 & LUT_stack_io_pop_30 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 3816:69 stackmanage_35.scala 3817:29]
  wire [31:0] _GEN_689 = _T_105 & LUT_stack_io_pop_30 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 3816:69 stackmanage_35.scala 3818:28]
  wire [31:0] _GEN_691 = _T_105 & LUT_stack_io_pop_30 ? 32'h0 : _GEN_679; // @[stackmanage_35.scala 3816:69 stackmanage_35.scala 3879:29]
  wire [31:0] _GEN_692 = _T_105 & LUT_stack_io_pop_30 ? 32'h0 : _GEN_680; // @[stackmanage_35.scala 3816:69 stackmanage_35.scala 3880:28]
  wire [31:0] _GEN_693 = _T_105 & LUT_stack_io_pop_30 ? 32'h0 : _GEN_682; // @[stackmanage_35.scala 3816:69 stackmanage_35.scala 3881:29]
  wire [31:0] _GEN_694 = _T_105 & LUT_stack_io_pop_30 ? 32'h0 : _GEN_683; // @[stackmanage_35.scala 3816:69 stackmanage_35.scala 3882:28]
  wire [31:0] _GEN_695 = _T_105 & LUT_stack_io_pop_30 ? 32'h0 : _GEN_684; // @[stackmanage_35.scala 3816:69 stackmanage_35.scala 3883:29]
  wire [31:0] _GEN_696 = _T_105 & LUT_stack_io_pop_30 ? 32'h0 : _GEN_685; // @[stackmanage_35.scala 3816:69 stackmanage_35.scala 3884:28]
  wire [31:0] _GEN_697 = _T_105 & LUT_stack_io_pop_30 ? 32'h0 : _GEN_686; // @[stackmanage_35.scala 3816:69 stackmanage_35.scala 3885:29]
  wire [31:0] _GEN_698 = _T_105 & LUT_stack_io_pop_30 ? 32'h0 : _GEN_687; // @[stackmanage_35.scala 3816:69 stackmanage_35.scala 3886:28]
  wire [31:0] _GEN_699 = _T_105 & LUT_stack_io_pop_29 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 3745:69 stackmanage_35.scala 3746:29]
  wire [31:0] _GEN_700 = _T_105 & LUT_stack_io_pop_29 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 3745:69 stackmanage_35.scala 3747:28]
  wire [31:0] _GEN_702 = _T_105 & LUT_stack_io_pop_29 ? 32'h0 : _GEN_688; // @[stackmanage_35.scala 3745:69 stackmanage_35.scala 3806:29]
  wire [31:0] _GEN_703 = _T_105 & LUT_stack_io_pop_29 ? 32'h0 : _GEN_689; // @[stackmanage_35.scala 3745:69 stackmanage_35.scala 3807:29]
  wire [31:0] _GEN_704 = _T_105 & LUT_stack_io_pop_29 ? 32'h0 : _GEN_691; // @[stackmanage_35.scala 3745:69 stackmanage_35.scala 3808:29]
  wire [31:0] _GEN_705 = _T_105 & LUT_stack_io_pop_29 ? 32'h0 : _GEN_692; // @[stackmanage_35.scala 3745:69 stackmanage_35.scala 3809:28]
  wire [31:0] _GEN_706 = _T_105 & LUT_stack_io_pop_29 ? 32'h0 : _GEN_693; // @[stackmanage_35.scala 3745:69 stackmanage_35.scala 3810:29]
  wire [31:0] _GEN_707 = _T_105 & LUT_stack_io_pop_29 ? 32'h0 : _GEN_694; // @[stackmanage_35.scala 3745:69 stackmanage_35.scala 3811:28]
  wire [31:0] _GEN_708 = _T_105 & LUT_stack_io_pop_29 ? 32'h0 : _GEN_695; // @[stackmanage_35.scala 3745:69 stackmanage_35.scala 3812:29]
  wire [31:0] _GEN_709 = _T_105 & LUT_stack_io_pop_29 ? 32'h0 : _GEN_696; // @[stackmanage_35.scala 3745:69 stackmanage_35.scala 3813:28]
  wire [31:0] _GEN_710 = _T_105 & LUT_stack_io_pop_29 ? 32'h0 : _GEN_697; // @[stackmanage_35.scala 3745:69 stackmanage_35.scala 3814:29]
  wire [31:0] _GEN_711 = _T_105 & LUT_stack_io_pop_29 ? 32'h0 : _GEN_698; // @[stackmanage_35.scala 3745:69 stackmanage_35.scala 3815:28]
  wire [31:0] _GEN_712 = _T_105 & LUT_stack_io_pop_28 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 3674:70 stackmanage_35.scala 3675:29]
  wire [31:0] _GEN_713 = _T_105 & LUT_stack_io_pop_28 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 3674:70 stackmanage_35.scala 3676:28]
  wire [31:0] _GEN_715 = _T_105 & LUT_stack_io_pop_28 ? 32'h0 : _GEN_699; // @[stackmanage_35.scala 3674:70 stackmanage_35.scala 3733:29]
  wire [31:0] _GEN_716 = _T_105 & LUT_stack_io_pop_28 ? 32'h0 : _GEN_700; // @[stackmanage_35.scala 3674:70 stackmanage_35.scala 3734:28]
  wire [31:0] _GEN_717 = _T_105 & LUT_stack_io_pop_28 ? 32'h0 : _GEN_702; // @[stackmanage_35.scala 3674:70 stackmanage_35.scala 3735:29]
  wire [31:0] _GEN_718 = _T_105 & LUT_stack_io_pop_28 ? 32'h0 : _GEN_703; // @[stackmanage_35.scala 3674:70 stackmanage_35.scala 3736:29]
  wire [31:0] _GEN_719 = _T_105 & LUT_stack_io_pop_28 ? 32'h0 : _GEN_704; // @[stackmanage_35.scala 3674:70 stackmanage_35.scala 3737:29]
  wire [31:0] _GEN_720 = _T_105 & LUT_stack_io_pop_28 ? 32'h0 : _GEN_705; // @[stackmanage_35.scala 3674:70 stackmanage_35.scala 3738:28]
  wire [31:0] _GEN_721 = _T_105 & LUT_stack_io_pop_28 ? 32'h0 : _GEN_706; // @[stackmanage_35.scala 3674:70 stackmanage_35.scala 3739:29]
  wire [31:0] _GEN_722 = _T_105 & LUT_stack_io_pop_28 ? 32'h0 : _GEN_707; // @[stackmanage_35.scala 3674:70 stackmanage_35.scala 3740:28]
  wire [31:0] _GEN_723 = _T_105 & LUT_stack_io_pop_28 ? 32'h0 : _GEN_708; // @[stackmanage_35.scala 3674:70 stackmanage_35.scala 3741:29]
  wire [31:0] _GEN_724 = _T_105 & LUT_stack_io_pop_28 ? 32'h0 : _GEN_709; // @[stackmanage_35.scala 3674:70 stackmanage_35.scala 3742:28]
  wire [31:0] _GEN_725 = _T_105 & LUT_stack_io_pop_28 ? 32'h0 : _GEN_710; // @[stackmanage_35.scala 3674:70 stackmanage_35.scala 3743:29]
  wire [31:0] _GEN_726 = _T_105 & LUT_stack_io_pop_28 ? 32'h0 : _GEN_711; // @[stackmanage_35.scala 3674:70 stackmanage_35.scala 3744:28]
  wire [31:0] _GEN_727 = _T_105 & LUT_stack_io_pop_27 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 3603:69 stackmanage_35.scala 3604:29]
  wire [31:0] _GEN_728 = _T_105 & LUT_stack_io_pop_27 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 3603:69 stackmanage_35.scala 3605:28]
  wire [31:0] _GEN_730 = _T_105 & LUT_stack_io_pop_27 ? 32'h0 : _GEN_712; // @[stackmanage_35.scala 3603:69 stackmanage_35.scala 3660:29]
  wire [31:0] _GEN_731 = _T_105 & LUT_stack_io_pop_27 ? 32'h0 : _GEN_713; // @[stackmanage_35.scala 3603:69 stackmanage_35.scala 3661:28]
  wire [31:0] _GEN_732 = _T_105 & LUT_stack_io_pop_27 ? 32'h0 : _GEN_715; // @[stackmanage_35.scala 3603:69 stackmanage_35.scala 3662:29]
  wire [31:0] _GEN_733 = _T_105 & LUT_stack_io_pop_27 ? 32'h0 : _GEN_716; // @[stackmanage_35.scala 3603:69 stackmanage_35.scala 3663:28]
  wire [31:0] _GEN_734 = _T_105 & LUT_stack_io_pop_27 ? 32'h0 : _GEN_717; // @[stackmanage_35.scala 3603:69 stackmanage_35.scala 3664:29]
  wire [31:0] _GEN_735 = _T_105 & LUT_stack_io_pop_27 ? 32'h0 : _GEN_718; // @[stackmanage_35.scala 3603:69 stackmanage_35.scala 3665:29]
  wire [31:0] _GEN_736 = _T_105 & LUT_stack_io_pop_27 ? 32'h0 : _GEN_719; // @[stackmanage_35.scala 3603:69 stackmanage_35.scala 3666:29]
  wire [31:0] _GEN_737 = _T_105 & LUT_stack_io_pop_27 ? 32'h0 : _GEN_720; // @[stackmanage_35.scala 3603:69 stackmanage_35.scala 3667:28]
  wire [31:0] _GEN_738 = _T_105 & LUT_stack_io_pop_27 ? 32'h0 : _GEN_721; // @[stackmanage_35.scala 3603:69 stackmanage_35.scala 3668:29]
  wire [31:0] _GEN_739 = _T_105 & LUT_stack_io_pop_27 ? 32'h0 : _GEN_722; // @[stackmanage_35.scala 3603:69 stackmanage_35.scala 3669:28]
  wire [31:0] _GEN_740 = _T_105 & LUT_stack_io_pop_27 ? 32'h0 : _GEN_723; // @[stackmanage_35.scala 3603:69 stackmanage_35.scala 3670:29]
  wire [31:0] _GEN_741 = _T_105 & LUT_stack_io_pop_27 ? 32'h0 : _GEN_724; // @[stackmanage_35.scala 3603:69 stackmanage_35.scala 3671:28]
  wire [31:0] _GEN_742 = _T_105 & LUT_stack_io_pop_27 ? 32'h0 : _GEN_725; // @[stackmanage_35.scala 3603:69 stackmanage_35.scala 3672:29]
  wire [31:0] _GEN_743 = _T_105 & LUT_stack_io_pop_27 ? 32'h0 : _GEN_726; // @[stackmanage_35.scala 3603:69 stackmanage_35.scala 3673:28]
  wire [31:0] _GEN_744 = _T_105 & LUT_stack_io_pop_26 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 3532:70 stackmanage_35.scala 3533:29]
  wire [31:0] _GEN_745 = _T_105 & LUT_stack_io_pop_26 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 3532:70 stackmanage_35.scala 3534:28]
  wire [31:0] _GEN_747 = _T_105 & LUT_stack_io_pop_26 ? 32'h0 : _GEN_727; // @[stackmanage_35.scala 3532:70 stackmanage_35.scala 3587:29]
  wire [31:0] _GEN_748 = _T_105 & LUT_stack_io_pop_26 ? 32'h0 : _GEN_728; // @[stackmanage_35.scala 3532:70 stackmanage_35.scala 3588:28]
  wire [31:0] _GEN_749 = _T_105 & LUT_stack_io_pop_26 ? 32'h0 : _GEN_730; // @[stackmanage_35.scala 3532:70 stackmanage_35.scala 3589:29]
  wire [31:0] _GEN_750 = _T_105 & LUT_stack_io_pop_26 ? 32'h0 : _GEN_731; // @[stackmanage_35.scala 3532:70 stackmanage_35.scala 3590:28]
  wire [31:0] _GEN_751 = _T_105 & LUT_stack_io_pop_26 ? 32'h0 : _GEN_732; // @[stackmanage_35.scala 3532:70 stackmanage_35.scala 3591:29]
  wire [31:0] _GEN_752 = _T_105 & LUT_stack_io_pop_26 ? 32'h0 : _GEN_733; // @[stackmanage_35.scala 3532:70 stackmanage_35.scala 3592:28]
  wire [31:0] _GEN_753 = _T_105 & LUT_stack_io_pop_26 ? 32'h0 : _GEN_734; // @[stackmanage_35.scala 3532:70 stackmanage_35.scala 3593:29]
  wire [31:0] _GEN_754 = _T_105 & LUT_stack_io_pop_26 ? 32'h0 : _GEN_735; // @[stackmanage_35.scala 3532:70 stackmanage_35.scala 3594:29]
  wire [31:0] _GEN_755 = _T_105 & LUT_stack_io_pop_26 ? 32'h0 : _GEN_736; // @[stackmanage_35.scala 3532:70 stackmanage_35.scala 3595:29]
  wire [31:0] _GEN_756 = _T_105 & LUT_stack_io_pop_26 ? 32'h0 : _GEN_737; // @[stackmanage_35.scala 3532:70 stackmanage_35.scala 3596:28]
  wire [31:0] _GEN_757 = _T_105 & LUT_stack_io_pop_26 ? 32'h0 : _GEN_738; // @[stackmanage_35.scala 3532:70 stackmanage_35.scala 3597:29]
  wire [31:0] _GEN_758 = _T_105 & LUT_stack_io_pop_26 ? 32'h0 : _GEN_739; // @[stackmanage_35.scala 3532:70 stackmanage_35.scala 3598:28]
  wire [31:0] _GEN_759 = _T_105 & LUT_stack_io_pop_26 ? 32'h0 : _GEN_740; // @[stackmanage_35.scala 3532:70 stackmanage_35.scala 3599:29]
  wire [31:0] _GEN_760 = _T_105 & LUT_stack_io_pop_26 ? 32'h0 : _GEN_741; // @[stackmanage_35.scala 3532:70 stackmanage_35.scala 3600:28]
  wire [31:0] _GEN_761 = _T_105 & LUT_stack_io_pop_26 ? 32'h0 : _GEN_742; // @[stackmanage_35.scala 3532:70 stackmanage_35.scala 3601:29]
  wire [31:0] _GEN_762 = _T_105 & LUT_stack_io_pop_26 ? 32'h0 : _GEN_743; // @[stackmanage_35.scala 3532:70 stackmanage_35.scala 3602:28]
  wire [31:0] _GEN_763 = _T_105 & LUT_stack_io_pop_25 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 3461:69 stackmanage_35.scala 3462:29]
  wire [31:0] _GEN_764 = _T_105 & LUT_stack_io_pop_25 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 3461:69 stackmanage_35.scala 3463:28]
  wire [31:0] _GEN_766 = _T_105 & LUT_stack_io_pop_25 ? 32'h0 : _GEN_744; // @[stackmanage_35.scala 3461:69 stackmanage_35.scala 3514:29]
  wire [31:0] _GEN_767 = _T_105 & LUT_stack_io_pop_25 ? 32'h0 : _GEN_745; // @[stackmanage_35.scala 3461:69 stackmanage_35.scala 3515:28]
  wire [31:0] _GEN_768 = _T_105 & LUT_stack_io_pop_25 ? 32'h0 : _GEN_747; // @[stackmanage_35.scala 3461:69 stackmanage_35.scala 3516:29]
  wire [31:0] _GEN_769 = _T_105 & LUT_stack_io_pop_25 ? 32'h0 : _GEN_748; // @[stackmanage_35.scala 3461:69 stackmanage_35.scala 3517:28]
  wire [31:0] _GEN_770 = _T_105 & LUT_stack_io_pop_25 ? 32'h0 : _GEN_749; // @[stackmanage_35.scala 3461:69 stackmanage_35.scala 3518:29]
  wire [31:0] _GEN_771 = _T_105 & LUT_stack_io_pop_25 ? 32'h0 : _GEN_750; // @[stackmanage_35.scala 3461:69 stackmanage_35.scala 3519:28]
  wire [31:0] _GEN_772 = _T_105 & LUT_stack_io_pop_25 ? 32'h0 : _GEN_751; // @[stackmanage_35.scala 3461:69 stackmanage_35.scala 3520:29]
  wire [31:0] _GEN_773 = _T_105 & LUT_stack_io_pop_25 ? 32'h0 : _GEN_752; // @[stackmanage_35.scala 3461:69 stackmanage_35.scala 3521:28]
  wire [31:0] _GEN_774 = _T_105 & LUT_stack_io_pop_25 ? 32'h0 : _GEN_753; // @[stackmanage_35.scala 3461:69 stackmanage_35.scala 3522:29]
  wire [31:0] _GEN_775 = _T_105 & LUT_stack_io_pop_25 ? 32'h0 : _GEN_754; // @[stackmanage_35.scala 3461:69 stackmanage_35.scala 3523:29]
  wire [31:0] _GEN_776 = _T_105 & LUT_stack_io_pop_25 ? 32'h0 : _GEN_755; // @[stackmanage_35.scala 3461:69 stackmanage_35.scala 3524:29]
  wire [31:0] _GEN_777 = _T_105 & LUT_stack_io_pop_25 ? 32'h0 : _GEN_756; // @[stackmanage_35.scala 3461:69 stackmanage_35.scala 3525:28]
  wire [31:0] _GEN_778 = _T_105 & LUT_stack_io_pop_25 ? 32'h0 : _GEN_757; // @[stackmanage_35.scala 3461:69 stackmanage_35.scala 3526:29]
  wire [31:0] _GEN_779 = _T_105 & LUT_stack_io_pop_25 ? 32'h0 : _GEN_758; // @[stackmanage_35.scala 3461:69 stackmanage_35.scala 3527:28]
  wire [31:0] _GEN_780 = _T_105 & LUT_stack_io_pop_25 ? 32'h0 : _GEN_759; // @[stackmanage_35.scala 3461:69 stackmanage_35.scala 3528:29]
  wire [31:0] _GEN_781 = _T_105 & LUT_stack_io_pop_25 ? 32'h0 : _GEN_760; // @[stackmanage_35.scala 3461:69 stackmanage_35.scala 3529:28]
  wire [31:0] _GEN_782 = _T_105 & LUT_stack_io_pop_25 ? 32'h0 : _GEN_761; // @[stackmanage_35.scala 3461:69 stackmanage_35.scala 3530:29]
  wire [31:0] _GEN_783 = _T_105 & LUT_stack_io_pop_25 ? 32'h0 : _GEN_762; // @[stackmanage_35.scala 3461:69 stackmanage_35.scala 3531:28]
  wire [31:0] _GEN_784 = _T_105 & LUT_stack_io_pop_24 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 3390:69 stackmanage_35.scala 3391:29]
  wire [31:0] _GEN_785 = _T_105 & LUT_stack_io_pop_24 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 3390:69 stackmanage_35.scala 3392:28]
  wire [31:0] _GEN_787 = _T_105 & LUT_stack_io_pop_24 ? 32'h0 : _GEN_763; // @[stackmanage_35.scala 3390:69 stackmanage_35.scala 3441:29]
  wire [31:0] _GEN_788 = _T_105 & LUT_stack_io_pop_24 ? 32'h0 : _GEN_764; // @[stackmanage_35.scala 3390:69 stackmanage_35.scala 3442:28]
  wire [31:0] _GEN_789 = _T_105 & LUT_stack_io_pop_24 ? 32'h0 : _GEN_766; // @[stackmanage_35.scala 3390:69 stackmanage_35.scala 3443:29]
  wire [31:0] _GEN_790 = _T_105 & LUT_stack_io_pop_24 ? 32'h0 : _GEN_767; // @[stackmanage_35.scala 3390:69 stackmanage_35.scala 3444:28]
  wire [31:0] _GEN_791 = _T_105 & LUT_stack_io_pop_24 ? 32'h0 : _GEN_768; // @[stackmanage_35.scala 3390:69 stackmanage_35.scala 3445:29]
  wire [31:0] _GEN_792 = _T_105 & LUT_stack_io_pop_24 ? 32'h0 : _GEN_769; // @[stackmanage_35.scala 3390:69 stackmanage_35.scala 3446:28]
  wire [31:0] _GEN_793 = _T_105 & LUT_stack_io_pop_24 ? 32'h0 : _GEN_770; // @[stackmanage_35.scala 3390:69 stackmanage_35.scala 3447:29]
  wire [31:0] _GEN_794 = _T_105 & LUT_stack_io_pop_24 ? 32'h0 : _GEN_771; // @[stackmanage_35.scala 3390:69 stackmanage_35.scala 3448:28]
  wire [31:0] _GEN_795 = _T_105 & LUT_stack_io_pop_24 ? 32'h0 : _GEN_772; // @[stackmanage_35.scala 3390:69 stackmanage_35.scala 3449:29]
  wire [31:0] _GEN_796 = _T_105 & LUT_stack_io_pop_24 ? 32'h0 : _GEN_773; // @[stackmanage_35.scala 3390:69 stackmanage_35.scala 3450:28]
  wire [31:0] _GEN_797 = _T_105 & LUT_stack_io_pop_24 ? 32'h0 : _GEN_774; // @[stackmanage_35.scala 3390:69 stackmanage_35.scala 3451:29]
  wire [31:0] _GEN_798 = _T_105 & LUT_stack_io_pop_24 ? 32'h0 : _GEN_775; // @[stackmanage_35.scala 3390:69 stackmanage_35.scala 3452:29]
  wire [31:0] _GEN_799 = _T_105 & LUT_stack_io_pop_24 ? 32'h0 : _GEN_776; // @[stackmanage_35.scala 3390:69 stackmanage_35.scala 3453:29]
  wire [31:0] _GEN_800 = _T_105 & LUT_stack_io_pop_24 ? 32'h0 : _GEN_777; // @[stackmanage_35.scala 3390:69 stackmanage_35.scala 3454:28]
  wire [31:0] _GEN_801 = _T_105 & LUT_stack_io_pop_24 ? 32'h0 : _GEN_778; // @[stackmanage_35.scala 3390:69 stackmanage_35.scala 3455:29]
  wire [31:0] _GEN_802 = _T_105 & LUT_stack_io_pop_24 ? 32'h0 : _GEN_779; // @[stackmanage_35.scala 3390:69 stackmanage_35.scala 3456:28]
  wire [31:0] _GEN_803 = _T_105 & LUT_stack_io_pop_24 ? 32'h0 : _GEN_780; // @[stackmanage_35.scala 3390:69 stackmanage_35.scala 3457:29]
  wire [31:0] _GEN_804 = _T_105 & LUT_stack_io_pop_24 ? 32'h0 : _GEN_781; // @[stackmanage_35.scala 3390:69 stackmanage_35.scala 3458:28]
  wire [31:0] _GEN_805 = _T_105 & LUT_stack_io_pop_24 ? 32'h0 : _GEN_782; // @[stackmanage_35.scala 3390:69 stackmanage_35.scala 3459:29]
  wire [31:0] _GEN_806 = _T_105 & LUT_stack_io_pop_24 ? 32'h0 : _GEN_783; // @[stackmanage_35.scala 3390:69 stackmanage_35.scala 3460:28]
  wire [31:0] _GEN_807 = _T_105 & LUT_stack_io_pop_23 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 3319:69 stackmanage_35.scala 3320:29]
  wire [31:0] _GEN_808 = _T_105 & LUT_stack_io_pop_23 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 3319:69 stackmanage_35.scala 3321:28]
  wire [31:0] _GEN_810 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_784; // @[stackmanage_35.scala 3319:69 stackmanage_35.scala 3368:29]
  wire [31:0] _GEN_811 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_785; // @[stackmanage_35.scala 3319:69 stackmanage_35.scala 3369:28]
  wire [31:0] _GEN_812 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_787; // @[stackmanage_35.scala 3319:69 stackmanage_35.scala 3370:29]
  wire [31:0] _GEN_813 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_788; // @[stackmanage_35.scala 3319:69 stackmanage_35.scala 3371:28]
  wire [31:0] _GEN_814 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_789; // @[stackmanage_35.scala 3319:69 stackmanage_35.scala 3372:29]
  wire [31:0] _GEN_815 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_790; // @[stackmanage_35.scala 3319:69 stackmanage_35.scala 3373:28]
  wire [31:0] _GEN_816 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_791; // @[stackmanage_35.scala 3319:69 stackmanage_35.scala 3374:29]
  wire [31:0] _GEN_817 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_792; // @[stackmanage_35.scala 3319:69 stackmanage_35.scala 3375:28]
  wire [31:0] _GEN_818 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_793; // @[stackmanage_35.scala 3319:69 stackmanage_35.scala 3376:29]
  wire [31:0] _GEN_819 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_794; // @[stackmanage_35.scala 3319:69 stackmanage_35.scala 3377:28]
  wire [31:0] _GEN_820 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_795; // @[stackmanage_35.scala 3319:69 stackmanage_35.scala 3378:29]
  wire [31:0] _GEN_821 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_796; // @[stackmanage_35.scala 3319:69 stackmanage_35.scala 3379:28]
  wire [31:0] _GEN_822 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_797; // @[stackmanage_35.scala 3319:69 stackmanage_35.scala 3380:29]
  wire [31:0] _GEN_823 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_798; // @[stackmanage_35.scala 3319:69 stackmanage_35.scala 3381:29]
  wire [31:0] _GEN_824 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_799; // @[stackmanage_35.scala 3319:69 stackmanage_35.scala 3382:29]
  wire [31:0] _GEN_825 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_800; // @[stackmanage_35.scala 3319:69 stackmanage_35.scala 3383:28]
  wire [31:0] _GEN_826 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_801; // @[stackmanage_35.scala 3319:69 stackmanage_35.scala 3384:29]
  wire [31:0] _GEN_827 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_802; // @[stackmanage_35.scala 3319:69 stackmanage_35.scala 3385:28]
  wire [31:0] _GEN_828 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_803; // @[stackmanage_35.scala 3319:69 stackmanage_35.scala 3386:29]
  wire [31:0] _GEN_829 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_804; // @[stackmanage_35.scala 3319:69 stackmanage_35.scala 3387:28]
  wire [31:0] _GEN_830 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_805; // @[stackmanage_35.scala 3319:69 stackmanage_35.scala 3388:29]
  wire [31:0] _GEN_831 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_806; // @[stackmanage_35.scala 3319:69 stackmanage_35.scala 3389:28]
  wire [31:0] _GEN_832 = _T_105 & LUT_stack_io_pop_22 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 3248:69 stackmanage_35.scala 3249:29]
  wire [31:0] _GEN_833 = _T_105 & LUT_stack_io_pop_22 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 3248:69 stackmanage_35.scala 3250:28]
  wire [31:0] _GEN_835 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_807; // @[stackmanage_35.scala 3248:69 stackmanage_35.scala 3295:29]
  wire [31:0] _GEN_836 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_808; // @[stackmanage_35.scala 3248:69 stackmanage_35.scala 3296:28]
  wire [31:0] _GEN_837 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_810; // @[stackmanage_35.scala 3248:69 stackmanage_35.scala 3297:29]
  wire [31:0] _GEN_838 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_811; // @[stackmanage_35.scala 3248:69 stackmanage_35.scala 3298:28]
  wire [31:0] _GEN_839 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_812; // @[stackmanage_35.scala 3248:69 stackmanage_35.scala 3299:29]
  wire [31:0] _GEN_840 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_813; // @[stackmanage_35.scala 3248:69 stackmanage_35.scala 3300:28]
  wire [31:0] _GEN_841 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_814; // @[stackmanage_35.scala 3248:69 stackmanage_35.scala 3301:29]
  wire [31:0] _GEN_842 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_815; // @[stackmanage_35.scala 3248:69 stackmanage_35.scala 3302:28]
  wire [31:0] _GEN_843 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_816; // @[stackmanage_35.scala 3248:69 stackmanage_35.scala 3303:29]
  wire [31:0] _GEN_844 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_817; // @[stackmanage_35.scala 3248:69 stackmanage_35.scala 3304:28]
  wire [31:0] _GEN_845 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_818; // @[stackmanage_35.scala 3248:69 stackmanage_35.scala 3305:29]
  wire [31:0] _GEN_846 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_819; // @[stackmanage_35.scala 3248:69 stackmanage_35.scala 3306:28]
  wire [31:0] _GEN_847 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_820; // @[stackmanage_35.scala 3248:69 stackmanage_35.scala 3307:29]
  wire [31:0] _GEN_848 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_821; // @[stackmanage_35.scala 3248:69 stackmanage_35.scala 3308:28]
  wire [31:0] _GEN_849 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_822; // @[stackmanage_35.scala 3248:69 stackmanage_35.scala 3309:29]
  wire [31:0] _GEN_850 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_823; // @[stackmanage_35.scala 3248:69 stackmanage_35.scala 3310:29]
  wire [31:0] _GEN_851 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_824; // @[stackmanage_35.scala 3248:69 stackmanage_35.scala 3311:29]
  wire [31:0] _GEN_852 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_825; // @[stackmanage_35.scala 3248:69 stackmanage_35.scala 3312:28]
  wire [31:0] _GEN_853 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_826; // @[stackmanage_35.scala 3248:69 stackmanage_35.scala 3313:29]
  wire [31:0] _GEN_854 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_827; // @[stackmanage_35.scala 3248:69 stackmanage_35.scala 3314:28]
  wire [31:0] _GEN_855 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_828; // @[stackmanage_35.scala 3248:69 stackmanage_35.scala 3315:29]
  wire [31:0] _GEN_856 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_829; // @[stackmanage_35.scala 3248:69 stackmanage_35.scala 3316:28]
  wire [31:0] _GEN_857 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_830; // @[stackmanage_35.scala 3248:69 stackmanage_35.scala 3317:29]
  wire [31:0] _GEN_858 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_831; // @[stackmanage_35.scala 3248:69 stackmanage_35.scala 3318:28]
  wire [31:0] _GEN_859 = _T_105 & LUT_stack_io_pop_21 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 3177:69 stackmanage_35.scala 3178:29]
  wire [31:0] _GEN_860 = _T_105 & LUT_stack_io_pop_21 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 3177:69 stackmanage_35.scala 3179:28]
  wire [31:0] _GEN_862 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_832; // @[stackmanage_35.scala 3177:69 stackmanage_35.scala 3222:29]
  wire [31:0] _GEN_863 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_833; // @[stackmanage_35.scala 3177:69 stackmanage_35.scala 3223:28]
  wire [31:0] _GEN_864 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_835; // @[stackmanage_35.scala 3177:69 stackmanage_35.scala 3224:29]
  wire [31:0] _GEN_865 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_836; // @[stackmanage_35.scala 3177:69 stackmanage_35.scala 3225:28]
  wire [31:0] _GEN_866 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_837; // @[stackmanage_35.scala 3177:69 stackmanage_35.scala 3226:29]
  wire [31:0] _GEN_867 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_838; // @[stackmanage_35.scala 3177:69 stackmanage_35.scala 3227:28]
  wire [31:0] _GEN_868 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_839; // @[stackmanage_35.scala 3177:69 stackmanage_35.scala 3228:29]
  wire [31:0] _GEN_869 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_840; // @[stackmanage_35.scala 3177:69 stackmanage_35.scala 3229:28]
  wire [31:0] _GEN_870 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_841; // @[stackmanage_35.scala 3177:69 stackmanage_35.scala 3230:29]
  wire [31:0] _GEN_871 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_842; // @[stackmanage_35.scala 3177:69 stackmanage_35.scala 3231:28]
  wire [31:0] _GEN_872 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_843; // @[stackmanage_35.scala 3177:69 stackmanage_35.scala 3232:29]
  wire [31:0] _GEN_873 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_844; // @[stackmanage_35.scala 3177:69 stackmanage_35.scala 3233:28]
  wire [31:0] _GEN_874 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_845; // @[stackmanage_35.scala 3177:69 stackmanage_35.scala 3234:29]
  wire [31:0] _GEN_875 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_846; // @[stackmanage_35.scala 3177:69 stackmanage_35.scala 3235:28]
  wire [31:0] _GEN_876 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_847; // @[stackmanage_35.scala 3177:69 stackmanage_35.scala 3236:29]
  wire [31:0] _GEN_877 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_848; // @[stackmanage_35.scala 3177:69 stackmanage_35.scala 3237:28]
  wire [31:0] _GEN_878 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_849; // @[stackmanage_35.scala 3177:69 stackmanage_35.scala 3238:29]
  wire [31:0] _GEN_879 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_850; // @[stackmanage_35.scala 3177:69 stackmanage_35.scala 3239:29]
  wire [31:0] _GEN_880 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_851; // @[stackmanage_35.scala 3177:69 stackmanage_35.scala 3240:29]
  wire [31:0] _GEN_881 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_852; // @[stackmanage_35.scala 3177:69 stackmanage_35.scala 3241:28]
  wire [31:0] _GEN_882 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_853; // @[stackmanage_35.scala 3177:69 stackmanage_35.scala 3242:29]
  wire [31:0] _GEN_883 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_854; // @[stackmanage_35.scala 3177:69 stackmanage_35.scala 3243:28]
  wire [31:0] _GEN_884 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_855; // @[stackmanage_35.scala 3177:69 stackmanage_35.scala 3244:29]
  wire [31:0] _GEN_885 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_856; // @[stackmanage_35.scala 3177:69 stackmanage_35.scala 3245:28]
  wire [31:0] _GEN_886 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_857; // @[stackmanage_35.scala 3177:69 stackmanage_35.scala 3246:29]
  wire [31:0] _GEN_887 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_858; // @[stackmanage_35.scala 3177:69 stackmanage_35.scala 3247:28]
  wire [31:0] _GEN_888 = _T_105 & LUT_stack_io_pop_20 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 3106:69 stackmanage_35.scala 3107:29]
  wire [31:0] _GEN_889 = _T_105 & LUT_stack_io_pop_20 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 3106:69 stackmanage_35.scala 3108:28]
  wire [31:0] _GEN_891 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_859; // @[stackmanage_35.scala 3106:69 stackmanage_35.scala 3149:29]
  wire [31:0] _GEN_892 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_860; // @[stackmanage_35.scala 3106:69 stackmanage_35.scala 3150:28]
  wire [31:0] _GEN_893 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_862; // @[stackmanage_35.scala 3106:69 stackmanage_35.scala 3151:29]
  wire [31:0] _GEN_894 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_863; // @[stackmanage_35.scala 3106:69 stackmanage_35.scala 3152:28]
  wire [31:0] _GEN_895 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_864; // @[stackmanage_35.scala 3106:69 stackmanage_35.scala 3153:29]
  wire [31:0] _GEN_896 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_865; // @[stackmanage_35.scala 3106:69 stackmanage_35.scala 3154:28]
  wire [31:0] _GEN_897 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_866; // @[stackmanage_35.scala 3106:69 stackmanage_35.scala 3155:29]
  wire [31:0] _GEN_898 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_867; // @[stackmanage_35.scala 3106:69 stackmanage_35.scala 3156:28]
  wire [31:0] _GEN_899 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_868; // @[stackmanage_35.scala 3106:69 stackmanage_35.scala 3157:29]
  wire [31:0] _GEN_900 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_869; // @[stackmanage_35.scala 3106:69 stackmanage_35.scala 3158:28]
  wire [31:0] _GEN_901 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_870; // @[stackmanage_35.scala 3106:69 stackmanage_35.scala 3159:29]
  wire [31:0] _GEN_902 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_871; // @[stackmanage_35.scala 3106:69 stackmanage_35.scala 3160:28]
  wire [31:0] _GEN_903 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_872; // @[stackmanage_35.scala 3106:69 stackmanage_35.scala 3161:29]
  wire [31:0] _GEN_904 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_873; // @[stackmanage_35.scala 3106:69 stackmanage_35.scala 3162:28]
  wire [31:0] _GEN_905 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_874; // @[stackmanage_35.scala 3106:69 stackmanage_35.scala 3163:29]
  wire [31:0] _GEN_906 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_875; // @[stackmanage_35.scala 3106:69 stackmanage_35.scala 3164:28]
  wire [31:0] _GEN_907 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_876; // @[stackmanage_35.scala 3106:69 stackmanage_35.scala 3165:29]
  wire [31:0] _GEN_908 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_877; // @[stackmanage_35.scala 3106:69 stackmanage_35.scala 3166:28]
  wire [31:0] _GEN_909 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_878; // @[stackmanage_35.scala 3106:69 stackmanage_35.scala 3167:29]
  wire [31:0] _GEN_910 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_879; // @[stackmanage_35.scala 3106:69 stackmanage_35.scala 3168:29]
  wire [31:0] _GEN_911 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_880; // @[stackmanage_35.scala 3106:69 stackmanage_35.scala 3169:29]
  wire [31:0] _GEN_912 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_881; // @[stackmanage_35.scala 3106:69 stackmanage_35.scala 3170:28]
  wire [31:0] _GEN_913 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_882; // @[stackmanage_35.scala 3106:69 stackmanage_35.scala 3171:29]
  wire [31:0] _GEN_914 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_883; // @[stackmanage_35.scala 3106:69 stackmanage_35.scala 3172:28]
  wire [31:0] _GEN_915 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_884; // @[stackmanage_35.scala 3106:69 stackmanage_35.scala 3173:29]
  wire [31:0] _GEN_916 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_885; // @[stackmanage_35.scala 3106:69 stackmanage_35.scala 3174:28]
  wire [31:0] _GEN_917 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_886; // @[stackmanage_35.scala 3106:69 stackmanage_35.scala 3175:29]
  wire [31:0] _GEN_918 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_887; // @[stackmanage_35.scala 3106:69 stackmanage_35.scala 3176:28]
  wire [31:0] _GEN_919 = _T_105 & LUT_stack_io_pop_19 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 3035:69 stackmanage_35.scala 3036:29]
  wire [31:0] _GEN_920 = _T_105 & LUT_stack_io_pop_19 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 3035:69 stackmanage_35.scala 3037:28]
  wire [31:0] _GEN_922 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_888; // @[stackmanage_35.scala 3035:69 stackmanage_35.scala 3076:29]
  wire [31:0] _GEN_923 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_889; // @[stackmanage_35.scala 3035:69 stackmanage_35.scala 3077:29]
  wire [31:0] _GEN_924 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_891; // @[stackmanage_35.scala 3035:69 stackmanage_35.scala 3078:29]
  wire [31:0] _GEN_925 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_892; // @[stackmanage_35.scala 3035:69 stackmanage_35.scala 3079:28]
  wire [31:0] _GEN_926 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_893; // @[stackmanage_35.scala 3035:69 stackmanage_35.scala 3080:29]
  wire [31:0] _GEN_927 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_894; // @[stackmanage_35.scala 3035:69 stackmanage_35.scala 3081:28]
  wire [31:0] _GEN_928 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_895; // @[stackmanage_35.scala 3035:69 stackmanage_35.scala 3082:29]
  wire [31:0] _GEN_929 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_896; // @[stackmanage_35.scala 3035:69 stackmanage_35.scala 3083:28]
  wire [31:0] _GEN_930 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_897; // @[stackmanage_35.scala 3035:69 stackmanage_35.scala 3084:29]
  wire [31:0] _GEN_931 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_898; // @[stackmanage_35.scala 3035:69 stackmanage_35.scala 3085:28]
  wire [31:0] _GEN_932 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_899; // @[stackmanage_35.scala 3035:69 stackmanage_35.scala 3086:29]
  wire [31:0] _GEN_933 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_900; // @[stackmanage_35.scala 3035:69 stackmanage_35.scala 3087:28]
  wire [31:0] _GEN_934 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_901; // @[stackmanage_35.scala 3035:69 stackmanage_35.scala 3088:29]
  wire [31:0] _GEN_935 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_902; // @[stackmanage_35.scala 3035:69 stackmanage_35.scala 3089:28]
  wire [31:0] _GEN_936 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_903; // @[stackmanage_35.scala 3035:69 stackmanage_35.scala 3090:29]
  wire [31:0] _GEN_937 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_904; // @[stackmanage_35.scala 3035:69 stackmanage_35.scala 3091:28]
  wire [31:0] _GEN_938 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_905; // @[stackmanage_35.scala 3035:69 stackmanage_35.scala 3092:29]
  wire [31:0] _GEN_939 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_906; // @[stackmanage_35.scala 3035:69 stackmanage_35.scala 3093:28]
  wire [31:0] _GEN_940 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_907; // @[stackmanage_35.scala 3035:69 stackmanage_35.scala 3094:29]
  wire [31:0] _GEN_941 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_908; // @[stackmanage_35.scala 3035:69 stackmanage_35.scala 3095:28]
  wire [31:0] _GEN_942 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_909; // @[stackmanage_35.scala 3035:69 stackmanage_35.scala 3096:29]
  wire [31:0] _GEN_943 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_910; // @[stackmanage_35.scala 3035:69 stackmanage_35.scala 3097:29]
  wire [31:0] _GEN_944 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_911; // @[stackmanage_35.scala 3035:69 stackmanage_35.scala 3098:29]
  wire [31:0] _GEN_945 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_912; // @[stackmanage_35.scala 3035:69 stackmanage_35.scala 3099:28]
  wire [31:0] _GEN_946 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_913; // @[stackmanage_35.scala 3035:69 stackmanage_35.scala 3100:29]
  wire [31:0] _GEN_947 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_914; // @[stackmanage_35.scala 3035:69 stackmanage_35.scala 3101:28]
  wire [31:0] _GEN_948 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_915; // @[stackmanage_35.scala 3035:69 stackmanage_35.scala 3102:29]
  wire [31:0] _GEN_949 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_916; // @[stackmanage_35.scala 3035:69 stackmanage_35.scala 3103:28]
  wire [31:0] _GEN_950 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_917; // @[stackmanage_35.scala 3035:69 stackmanage_35.scala 3104:29]
  wire [31:0] _GEN_951 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_918; // @[stackmanage_35.scala 3035:69 stackmanage_35.scala 3105:28]
  wire [31:0] _GEN_952 = _T_105 & LUT_stack_io_pop_18 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 2964:69 stackmanage_35.scala 2965:29]
  wire [31:0] _GEN_953 = _T_105 & LUT_stack_io_pop_18 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 2964:69 stackmanage_35.scala 2966:28]
  wire [31:0] _GEN_955 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_919; // @[stackmanage_35.scala 2964:69 stackmanage_35.scala 3003:29]
  wire [31:0] _GEN_956 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_920; // @[stackmanage_35.scala 2964:69 stackmanage_35.scala 3004:28]
  wire [31:0] _GEN_957 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_922; // @[stackmanage_35.scala 2964:69 stackmanage_35.scala 3005:29]
  wire [31:0] _GEN_958 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_923; // @[stackmanage_35.scala 2964:69 stackmanage_35.scala 3006:29]
  wire [31:0] _GEN_959 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_924; // @[stackmanage_35.scala 2964:69 stackmanage_35.scala 3007:29]
  wire [31:0] _GEN_960 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_925; // @[stackmanage_35.scala 2964:69 stackmanage_35.scala 3008:28]
  wire [31:0] _GEN_961 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_926; // @[stackmanage_35.scala 2964:69 stackmanage_35.scala 3009:29]
  wire [31:0] _GEN_962 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_927; // @[stackmanage_35.scala 2964:69 stackmanage_35.scala 3010:28]
  wire [31:0] _GEN_963 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_928; // @[stackmanage_35.scala 2964:69 stackmanage_35.scala 3011:29]
  wire [31:0] _GEN_964 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_929; // @[stackmanage_35.scala 2964:69 stackmanage_35.scala 3012:28]
  wire [31:0] _GEN_965 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_930; // @[stackmanage_35.scala 2964:69 stackmanage_35.scala 3013:29]
  wire [31:0] _GEN_966 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_931; // @[stackmanage_35.scala 2964:69 stackmanage_35.scala 3014:28]
  wire [31:0] _GEN_967 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_932; // @[stackmanage_35.scala 2964:69 stackmanage_35.scala 3015:29]
  wire [31:0] _GEN_968 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_933; // @[stackmanage_35.scala 2964:69 stackmanage_35.scala 3016:28]
  wire [31:0] _GEN_969 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_934; // @[stackmanage_35.scala 2964:69 stackmanage_35.scala 3017:29]
  wire [31:0] _GEN_970 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_935; // @[stackmanage_35.scala 2964:69 stackmanage_35.scala 3018:28]
  wire [31:0] _GEN_971 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_936; // @[stackmanage_35.scala 2964:69 stackmanage_35.scala 3019:29]
  wire [31:0] _GEN_972 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_937; // @[stackmanage_35.scala 2964:69 stackmanage_35.scala 3020:28]
  wire [31:0] _GEN_973 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_938; // @[stackmanage_35.scala 2964:69 stackmanage_35.scala 3021:29]
  wire [31:0] _GEN_974 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_939; // @[stackmanage_35.scala 2964:69 stackmanage_35.scala 3022:28]
  wire [31:0] _GEN_975 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_940; // @[stackmanage_35.scala 2964:69 stackmanage_35.scala 3023:29]
  wire [31:0] _GEN_976 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_941; // @[stackmanage_35.scala 2964:69 stackmanage_35.scala 3024:28]
  wire [31:0] _GEN_977 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_942; // @[stackmanage_35.scala 2964:69 stackmanage_35.scala 3025:29]
  wire [31:0] _GEN_978 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_943; // @[stackmanage_35.scala 2964:69 stackmanage_35.scala 3026:29]
  wire [31:0] _GEN_979 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_944; // @[stackmanage_35.scala 2964:69 stackmanage_35.scala 3027:29]
  wire [31:0] _GEN_980 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_945; // @[stackmanage_35.scala 2964:69 stackmanage_35.scala 3028:28]
  wire [31:0] _GEN_981 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_946; // @[stackmanage_35.scala 2964:69 stackmanage_35.scala 3029:29]
  wire [31:0] _GEN_982 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_947; // @[stackmanage_35.scala 2964:69 stackmanage_35.scala 3030:28]
  wire [31:0] _GEN_983 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_948; // @[stackmanage_35.scala 2964:69 stackmanage_35.scala 3031:29]
  wire [31:0] _GEN_984 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_949; // @[stackmanage_35.scala 2964:69 stackmanage_35.scala 3032:28]
  wire [31:0] _GEN_985 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_950; // @[stackmanage_35.scala 2964:69 stackmanage_35.scala 3033:29]
  wire [31:0] _GEN_986 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_951; // @[stackmanage_35.scala 2964:69 stackmanage_35.scala 3034:28]
  wire [31:0] _GEN_987 = _T_105 & LUT_stack_io_pop_17 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 2893:69 stackmanage_35.scala 2894:29]
  wire [31:0] _GEN_988 = _T_105 & LUT_stack_io_pop_17 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 2893:69 stackmanage_35.scala 2895:28]
  wire [31:0] _GEN_990 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_952; // @[stackmanage_35.scala 2893:69 stackmanage_35.scala 2930:29]
  wire [31:0] _GEN_991 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_953; // @[stackmanage_35.scala 2893:69 stackmanage_35.scala 2931:28]
  wire [31:0] _GEN_992 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_955; // @[stackmanage_35.scala 2893:69 stackmanage_35.scala 2932:29]
  wire [31:0] _GEN_993 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_956; // @[stackmanage_35.scala 2893:69 stackmanage_35.scala 2933:28]
  wire [31:0] _GEN_994 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_957; // @[stackmanage_35.scala 2893:69 stackmanage_35.scala 2934:29]
  wire [31:0] _GEN_995 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_958; // @[stackmanage_35.scala 2893:69 stackmanage_35.scala 2935:29]
  wire [31:0] _GEN_996 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_959; // @[stackmanage_35.scala 2893:69 stackmanage_35.scala 2936:29]
  wire [31:0] _GEN_997 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_960; // @[stackmanage_35.scala 2893:69 stackmanage_35.scala 2937:28]
  wire [31:0] _GEN_998 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_961; // @[stackmanage_35.scala 2893:69 stackmanage_35.scala 2938:29]
  wire [31:0] _GEN_999 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_962; // @[stackmanage_35.scala 2893:69 stackmanage_35.scala 2939:28]
  wire [31:0] _GEN_1000 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_963; // @[stackmanage_35.scala 2893:69 stackmanage_35.scala 2940:29]
  wire [31:0] _GEN_1001 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_964; // @[stackmanage_35.scala 2893:69 stackmanage_35.scala 2941:28]
  wire [31:0] _GEN_1002 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_965; // @[stackmanage_35.scala 2893:69 stackmanage_35.scala 2942:29]
  wire [31:0] _GEN_1003 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_966; // @[stackmanage_35.scala 2893:69 stackmanage_35.scala 2943:28]
  wire [31:0] _GEN_1004 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_967; // @[stackmanage_35.scala 2893:69 stackmanage_35.scala 2944:29]
  wire [31:0] _GEN_1005 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_968; // @[stackmanage_35.scala 2893:69 stackmanage_35.scala 2945:28]
  wire [31:0] _GEN_1006 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_969; // @[stackmanage_35.scala 2893:69 stackmanage_35.scala 2946:29]
  wire [31:0] _GEN_1007 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_970; // @[stackmanage_35.scala 2893:69 stackmanage_35.scala 2947:28]
  wire [31:0] _GEN_1008 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_971; // @[stackmanage_35.scala 2893:69 stackmanage_35.scala 2948:29]
  wire [31:0] _GEN_1009 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_972; // @[stackmanage_35.scala 2893:69 stackmanage_35.scala 2949:28]
  wire [31:0] _GEN_1010 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_973; // @[stackmanage_35.scala 2893:69 stackmanage_35.scala 2950:29]
  wire [31:0] _GEN_1011 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_974; // @[stackmanage_35.scala 2893:69 stackmanage_35.scala 2951:28]
  wire [31:0] _GEN_1012 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_975; // @[stackmanage_35.scala 2893:69 stackmanage_35.scala 2952:29]
  wire [31:0] _GEN_1013 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_976; // @[stackmanage_35.scala 2893:69 stackmanage_35.scala 2953:28]
  wire [31:0] _GEN_1014 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_977; // @[stackmanage_35.scala 2893:69 stackmanage_35.scala 2954:29]
  wire [31:0] _GEN_1015 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_978; // @[stackmanage_35.scala 2893:69 stackmanage_35.scala 2955:29]
  wire [31:0] _GEN_1016 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_979; // @[stackmanage_35.scala 2893:69 stackmanage_35.scala 2956:29]
  wire [31:0] _GEN_1017 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_980; // @[stackmanage_35.scala 2893:69 stackmanage_35.scala 2957:28]
  wire [31:0] _GEN_1018 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_981; // @[stackmanage_35.scala 2893:69 stackmanage_35.scala 2958:29]
  wire [31:0] _GEN_1019 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_982; // @[stackmanage_35.scala 2893:69 stackmanage_35.scala 2959:28]
  wire [31:0] _GEN_1020 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_983; // @[stackmanage_35.scala 2893:69 stackmanage_35.scala 2960:29]
  wire [31:0] _GEN_1021 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_984; // @[stackmanage_35.scala 2893:69 stackmanage_35.scala 2961:28]
  wire [31:0] _GEN_1022 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_985; // @[stackmanage_35.scala 2893:69 stackmanage_35.scala 2962:29]
  wire [31:0] _GEN_1023 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_986; // @[stackmanage_35.scala 2893:69 stackmanage_35.scala 2963:28]
  wire [31:0] _GEN_1024 = _T_105 & LUT_stack_io_pop_16 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 2822:69 stackmanage_35.scala 2823:29]
  wire [31:0] _GEN_1025 = _T_105 & LUT_stack_io_pop_16 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 2822:69 stackmanage_35.scala 2824:28]
  wire [31:0] _GEN_1027 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_987; // @[stackmanage_35.scala 2822:69 stackmanage_35.scala 2857:29]
  wire [31:0] _GEN_1028 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_988; // @[stackmanage_35.scala 2822:69 stackmanage_35.scala 2858:28]
  wire [31:0] _GEN_1029 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_990; // @[stackmanage_35.scala 2822:69 stackmanage_35.scala 2859:29]
  wire [31:0] _GEN_1030 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_991; // @[stackmanage_35.scala 2822:69 stackmanage_35.scala 2860:28]
  wire [31:0] _GEN_1031 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_992; // @[stackmanage_35.scala 2822:69 stackmanage_35.scala 2861:29]
  wire [31:0] _GEN_1032 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_993; // @[stackmanage_35.scala 2822:69 stackmanage_35.scala 2862:28]
  wire [31:0] _GEN_1033 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_994; // @[stackmanage_35.scala 2822:69 stackmanage_35.scala 2863:29]
  wire [31:0] _GEN_1034 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_995; // @[stackmanage_35.scala 2822:69 stackmanage_35.scala 2864:29]
  wire [31:0] _GEN_1035 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_996; // @[stackmanage_35.scala 2822:69 stackmanage_35.scala 2865:29]
  wire [31:0] _GEN_1036 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_997; // @[stackmanage_35.scala 2822:69 stackmanage_35.scala 2866:28]
  wire [31:0] _GEN_1037 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_998; // @[stackmanage_35.scala 2822:69 stackmanage_35.scala 2867:29]
  wire [31:0] _GEN_1038 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_999; // @[stackmanage_35.scala 2822:69 stackmanage_35.scala 2868:28]
  wire [31:0] _GEN_1039 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1000; // @[stackmanage_35.scala 2822:69 stackmanage_35.scala 2869:29]
  wire [31:0] _GEN_1040 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1001; // @[stackmanage_35.scala 2822:69 stackmanage_35.scala 2870:28]
  wire [31:0] _GEN_1041 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1002; // @[stackmanage_35.scala 2822:69 stackmanage_35.scala 2871:29]
  wire [31:0] _GEN_1042 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1003; // @[stackmanage_35.scala 2822:69 stackmanage_35.scala 2872:28]
  wire [31:0] _GEN_1043 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1004; // @[stackmanage_35.scala 2822:69 stackmanage_35.scala 2873:29]
  wire [31:0] _GEN_1044 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1005; // @[stackmanage_35.scala 2822:69 stackmanage_35.scala 2874:28]
  wire [31:0] _GEN_1045 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1006; // @[stackmanage_35.scala 2822:69 stackmanage_35.scala 2875:29]
  wire [31:0] _GEN_1046 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1007; // @[stackmanage_35.scala 2822:69 stackmanage_35.scala 2876:28]
  wire [31:0] _GEN_1047 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1008; // @[stackmanage_35.scala 2822:69 stackmanage_35.scala 2877:29]
  wire [31:0] _GEN_1048 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1009; // @[stackmanage_35.scala 2822:69 stackmanage_35.scala 2878:28]
  wire [31:0] _GEN_1049 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1010; // @[stackmanage_35.scala 2822:69 stackmanage_35.scala 2879:29]
  wire [31:0] _GEN_1050 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1011; // @[stackmanage_35.scala 2822:69 stackmanage_35.scala 2880:28]
  wire [31:0] _GEN_1051 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1012; // @[stackmanage_35.scala 2822:69 stackmanage_35.scala 2881:29]
  wire [31:0] _GEN_1052 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1013; // @[stackmanage_35.scala 2822:69 stackmanage_35.scala 2882:28]
  wire [31:0] _GEN_1053 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1014; // @[stackmanage_35.scala 2822:69 stackmanage_35.scala 2883:29]
  wire [31:0] _GEN_1054 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1015; // @[stackmanage_35.scala 2822:69 stackmanage_35.scala 2884:29]
  wire [31:0] _GEN_1055 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1016; // @[stackmanage_35.scala 2822:69 stackmanage_35.scala 2885:29]
  wire [31:0] _GEN_1056 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1017; // @[stackmanage_35.scala 2822:69 stackmanage_35.scala 2886:28]
  wire [31:0] _GEN_1057 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1018; // @[stackmanage_35.scala 2822:69 stackmanage_35.scala 2887:29]
  wire [31:0] _GEN_1058 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1019; // @[stackmanage_35.scala 2822:69 stackmanage_35.scala 2888:28]
  wire [31:0] _GEN_1059 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1020; // @[stackmanage_35.scala 2822:69 stackmanage_35.scala 2889:29]
  wire [31:0] _GEN_1060 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1021; // @[stackmanage_35.scala 2822:69 stackmanage_35.scala 2890:28]
  wire [31:0] _GEN_1061 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1022; // @[stackmanage_35.scala 2822:69 stackmanage_35.scala 2891:29]
  wire [31:0] _GEN_1062 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1023; // @[stackmanage_35.scala 2822:69 stackmanage_35.scala 2892:28]
  wire [31:0] _GEN_1063 = _T_105 & LUT_stack_io_pop_15 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 2751:69 stackmanage_35.scala 2752:29]
  wire [31:0] _GEN_1064 = _T_105 & LUT_stack_io_pop_15 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 2751:69 stackmanage_35.scala 2753:28]
  wire [31:0] _GEN_1066 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1024; // @[stackmanage_35.scala 2751:69 stackmanage_35.scala 2784:29]
  wire [31:0] _GEN_1067 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1025; // @[stackmanage_35.scala 2751:69 stackmanage_35.scala 2785:28]
  wire [31:0] _GEN_1068 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1027; // @[stackmanage_35.scala 2751:69 stackmanage_35.scala 2786:29]
  wire [31:0] _GEN_1069 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1028; // @[stackmanage_35.scala 2751:69 stackmanage_35.scala 2787:28]
  wire [31:0] _GEN_1070 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1029; // @[stackmanage_35.scala 2751:69 stackmanage_35.scala 2788:29]
  wire [31:0] _GEN_1071 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1030; // @[stackmanage_35.scala 2751:69 stackmanage_35.scala 2789:28]
  wire [31:0] _GEN_1072 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1031; // @[stackmanage_35.scala 2751:69 stackmanage_35.scala 2790:29]
  wire [31:0] _GEN_1073 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1032; // @[stackmanage_35.scala 2751:69 stackmanage_35.scala 2791:28]
  wire [31:0] _GEN_1074 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1033; // @[stackmanage_35.scala 2751:69 stackmanage_35.scala 2792:29]
  wire [31:0] _GEN_1075 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1034; // @[stackmanage_35.scala 2751:69 stackmanage_35.scala 2793:29]
  wire [31:0] _GEN_1076 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1035; // @[stackmanage_35.scala 2751:69 stackmanage_35.scala 2794:29]
  wire [31:0] _GEN_1077 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1036; // @[stackmanage_35.scala 2751:69 stackmanage_35.scala 2795:28]
  wire [31:0] _GEN_1078 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1037; // @[stackmanage_35.scala 2751:69 stackmanage_35.scala 2796:29]
  wire [31:0] _GEN_1079 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1038; // @[stackmanage_35.scala 2751:69 stackmanage_35.scala 2797:28]
  wire [31:0] _GEN_1080 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1039; // @[stackmanage_35.scala 2751:69 stackmanage_35.scala 2798:29]
  wire [31:0] _GEN_1081 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1040; // @[stackmanage_35.scala 2751:69 stackmanage_35.scala 2799:28]
  wire [31:0] _GEN_1082 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1041; // @[stackmanage_35.scala 2751:69 stackmanage_35.scala 2800:29]
  wire [31:0] _GEN_1083 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1042; // @[stackmanage_35.scala 2751:69 stackmanage_35.scala 2801:28]
  wire [31:0] _GEN_1084 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1043; // @[stackmanage_35.scala 2751:69 stackmanage_35.scala 2802:29]
  wire [31:0] _GEN_1085 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1044; // @[stackmanage_35.scala 2751:69 stackmanage_35.scala 2803:28]
  wire [31:0] _GEN_1086 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1045; // @[stackmanage_35.scala 2751:69 stackmanage_35.scala 2804:29]
  wire [31:0] _GEN_1087 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1046; // @[stackmanage_35.scala 2751:69 stackmanage_35.scala 2805:28]
  wire [31:0] _GEN_1088 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1047; // @[stackmanage_35.scala 2751:69 stackmanage_35.scala 2806:29]
  wire [31:0] _GEN_1089 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1048; // @[stackmanage_35.scala 2751:69 stackmanage_35.scala 2807:28]
  wire [31:0] _GEN_1090 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1049; // @[stackmanage_35.scala 2751:69 stackmanage_35.scala 2808:29]
  wire [31:0] _GEN_1091 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1050; // @[stackmanage_35.scala 2751:69 stackmanage_35.scala 2809:28]
  wire [31:0] _GEN_1092 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1051; // @[stackmanage_35.scala 2751:69 stackmanage_35.scala 2810:29]
  wire [31:0] _GEN_1093 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1052; // @[stackmanage_35.scala 2751:69 stackmanage_35.scala 2811:28]
  wire [31:0] _GEN_1094 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1053; // @[stackmanage_35.scala 2751:69 stackmanage_35.scala 2812:29]
  wire [31:0] _GEN_1095 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1054; // @[stackmanage_35.scala 2751:69 stackmanage_35.scala 2813:29]
  wire [31:0] _GEN_1096 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1055; // @[stackmanage_35.scala 2751:69 stackmanage_35.scala 2814:29]
  wire [31:0] _GEN_1097 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1056; // @[stackmanage_35.scala 2751:69 stackmanage_35.scala 2815:28]
  wire [31:0] _GEN_1098 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1057; // @[stackmanage_35.scala 2751:69 stackmanage_35.scala 2816:29]
  wire [31:0] _GEN_1099 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1058; // @[stackmanage_35.scala 2751:69 stackmanage_35.scala 2817:28]
  wire [31:0] _GEN_1100 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1059; // @[stackmanage_35.scala 2751:69 stackmanage_35.scala 2818:29]
  wire [31:0] _GEN_1101 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1060; // @[stackmanage_35.scala 2751:69 stackmanage_35.scala 2819:28]
  wire [31:0] _GEN_1102 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1061; // @[stackmanage_35.scala 2751:69 stackmanage_35.scala 2820:29]
  wire [31:0] _GEN_1103 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1062; // @[stackmanage_35.scala 2751:69 stackmanage_35.scala 2821:28]
  wire [31:0] _GEN_1104 = _T_105 & LUT_stack_io_pop_14 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 2680:69 stackmanage_35.scala 2681:29]
  wire [31:0] _GEN_1105 = _T_105 & LUT_stack_io_pop_14 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 2680:69 stackmanage_35.scala 2682:28]
  wire [31:0] _GEN_1107 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1063; // @[stackmanage_35.scala 2680:69 stackmanage_35.scala 2711:29]
  wire [31:0] _GEN_1108 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1064; // @[stackmanage_35.scala 2680:69 stackmanage_35.scala 2712:28]
  wire [31:0] _GEN_1109 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1066; // @[stackmanage_35.scala 2680:69 stackmanage_35.scala 2713:29]
  wire [31:0] _GEN_1110 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1067; // @[stackmanage_35.scala 2680:69 stackmanage_35.scala 2714:28]
  wire [31:0] _GEN_1111 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1068; // @[stackmanage_35.scala 2680:69 stackmanage_35.scala 2715:29]
  wire [31:0] _GEN_1112 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1069; // @[stackmanage_35.scala 2680:69 stackmanage_35.scala 2716:28]
  wire [31:0] _GEN_1113 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1070; // @[stackmanage_35.scala 2680:69 stackmanage_35.scala 2717:29]
  wire [31:0] _GEN_1114 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1071; // @[stackmanage_35.scala 2680:69 stackmanage_35.scala 2718:28]
  wire [31:0] _GEN_1115 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1072; // @[stackmanage_35.scala 2680:69 stackmanage_35.scala 2719:29]
  wire [31:0] _GEN_1116 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1073; // @[stackmanage_35.scala 2680:69 stackmanage_35.scala 2720:28]
  wire [31:0] _GEN_1117 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1074; // @[stackmanage_35.scala 2680:69 stackmanage_35.scala 2721:29]
  wire [31:0] _GEN_1118 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1075; // @[stackmanage_35.scala 2680:69 stackmanage_35.scala 2722:29]
  wire [31:0] _GEN_1119 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1076; // @[stackmanage_35.scala 2680:69 stackmanage_35.scala 2723:29]
  wire [31:0] _GEN_1120 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1077; // @[stackmanage_35.scala 2680:69 stackmanage_35.scala 2724:28]
  wire [31:0] _GEN_1121 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1078; // @[stackmanage_35.scala 2680:69 stackmanage_35.scala 2725:29]
  wire [31:0] _GEN_1122 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1079; // @[stackmanage_35.scala 2680:69 stackmanage_35.scala 2726:28]
  wire [31:0] _GEN_1123 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1080; // @[stackmanage_35.scala 2680:69 stackmanage_35.scala 2727:29]
  wire [31:0] _GEN_1124 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1081; // @[stackmanage_35.scala 2680:69 stackmanage_35.scala 2728:28]
  wire [31:0] _GEN_1125 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1082; // @[stackmanage_35.scala 2680:69 stackmanage_35.scala 2729:29]
  wire [31:0] _GEN_1126 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1083; // @[stackmanage_35.scala 2680:69 stackmanage_35.scala 2730:28]
  wire [31:0] _GEN_1127 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1084; // @[stackmanage_35.scala 2680:69 stackmanage_35.scala 2731:29]
  wire [31:0] _GEN_1128 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1085; // @[stackmanage_35.scala 2680:69 stackmanage_35.scala 2732:28]
  wire [31:0] _GEN_1129 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1086; // @[stackmanage_35.scala 2680:69 stackmanage_35.scala 2733:29]
  wire [31:0] _GEN_1130 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1087; // @[stackmanage_35.scala 2680:69 stackmanage_35.scala 2734:28]
  wire [31:0] _GEN_1131 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1088; // @[stackmanage_35.scala 2680:69 stackmanage_35.scala 2735:29]
  wire [31:0] _GEN_1132 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1089; // @[stackmanage_35.scala 2680:69 stackmanage_35.scala 2736:28]
  wire [31:0] _GEN_1133 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1090; // @[stackmanage_35.scala 2680:69 stackmanage_35.scala 2737:29]
  wire [31:0] _GEN_1134 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1091; // @[stackmanage_35.scala 2680:69 stackmanage_35.scala 2738:28]
  wire [31:0] _GEN_1135 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1092; // @[stackmanage_35.scala 2680:69 stackmanage_35.scala 2739:29]
  wire [31:0] _GEN_1136 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1093; // @[stackmanage_35.scala 2680:69 stackmanage_35.scala 2740:28]
  wire [31:0] _GEN_1137 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1094; // @[stackmanage_35.scala 2680:69 stackmanage_35.scala 2741:29]
  wire [31:0] _GEN_1138 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1095; // @[stackmanage_35.scala 2680:69 stackmanage_35.scala 2742:29]
  wire [31:0] _GEN_1139 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1096; // @[stackmanage_35.scala 2680:69 stackmanage_35.scala 2743:29]
  wire [31:0] _GEN_1140 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1097; // @[stackmanage_35.scala 2680:69 stackmanage_35.scala 2744:28]
  wire [31:0] _GEN_1141 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1098; // @[stackmanage_35.scala 2680:69 stackmanage_35.scala 2745:29]
  wire [31:0] _GEN_1142 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1099; // @[stackmanage_35.scala 2680:69 stackmanage_35.scala 2746:28]
  wire [31:0] _GEN_1143 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1100; // @[stackmanage_35.scala 2680:69 stackmanage_35.scala 2747:29]
  wire [31:0] _GEN_1144 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1101; // @[stackmanage_35.scala 2680:69 stackmanage_35.scala 2748:28]
  wire [31:0] _GEN_1145 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1102; // @[stackmanage_35.scala 2680:69 stackmanage_35.scala 2749:29]
  wire [31:0] _GEN_1146 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1103; // @[stackmanage_35.scala 2680:69 stackmanage_35.scala 2750:28]
  wire [31:0] _GEN_1147 = _T_105 & LUT_stack_io_pop_13 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2610:29]
  wire [31:0] _GEN_1148 = _T_105 & LUT_stack_io_pop_13 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2611:28]
  wire [31:0] _GEN_1150 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1104; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2638:29]
  wire [31:0] _GEN_1151 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1105; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2639:28]
  wire [31:0] _GEN_1152 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1107; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2640:29]
  wire [31:0] _GEN_1153 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1108; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2641:28]
  wire [31:0] _GEN_1154 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1109; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2642:29]
  wire [31:0] _GEN_1155 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1110; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2643:28]
  wire [31:0] _GEN_1156 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1111; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2644:29]
  wire [31:0] _GEN_1157 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1112; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2645:28]
  wire [31:0] _GEN_1158 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1113; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2646:29]
  wire [31:0] _GEN_1159 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1114; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2647:28]
  wire [31:0] _GEN_1160 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1115; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2648:29]
  wire [31:0] _GEN_1161 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1116; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2649:28]
  wire [31:0] _GEN_1162 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1117; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2650:29]
  wire [31:0] _GEN_1163 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1118; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2651:29]
  wire [31:0] _GEN_1164 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1119; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2652:29]
  wire [31:0] _GEN_1165 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1120; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2653:28]
  wire [31:0] _GEN_1166 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1121; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2654:29]
  wire [31:0] _GEN_1167 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1122; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2655:28]
  wire [31:0] _GEN_1168 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1123; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2656:29]
  wire [31:0] _GEN_1169 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1124; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2657:28]
  wire [31:0] _GEN_1170 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1125; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2658:29]
  wire [31:0] _GEN_1171 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1126; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2659:28]
  wire [31:0] _GEN_1172 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1127; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2660:29]
  wire [31:0] _GEN_1173 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1128; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2661:28]
  wire [31:0] _GEN_1174 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1129; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2662:29]
  wire [31:0] _GEN_1175 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1130; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2663:28]
  wire [31:0] _GEN_1176 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1131; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2664:29]
  wire [31:0] _GEN_1177 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1132; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2665:28]
  wire [31:0] _GEN_1178 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1133; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2666:29]
  wire [31:0] _GEN_1179 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1134; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2667:28]
  wire [31:0] _GEN_1180 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1135; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2668:29]
  wire [31:0] _GEN_1181 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1136; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2669:28]
  wire [31:0] _GEN_1182 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1137; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2670:29]
  wire [31:0] _GEN_1183 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1138; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2671:29]
  wire [31:0] _GEN_1184 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1139; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2672:29]
  wire [31:0] _GEN_1185 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1140; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2673:28]
  wire [31:0] _GEN_1186 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1141; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2674:29]
  wire [31:0] _GEN_1187 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1142; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2675:28]
  wire [31:0] _GEN_1188 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1143; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2676:29]
  wire [31:0] _GEN_1189 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1144; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2677:28]
  wire [31:0] _GEN_1190 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1145; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2678:29]
  wire [31:0] _GEN_1191 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1146; // @[stackmanage_35.scala 2609:69 stackmanage_35.scala 2679:28]
  wire [31:0] _GEN_1192 = _T_105 & LUT_stack_io_pop_12 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2539:29]
  wire [31:0] _GEN_1193 = _T_105 & LUT_stack_io_pop_12 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2540:28]
  wire [31:0] _GEN_1195 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1147; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2565:29]
  wire [31:0] _GEN_1196 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1148; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2566:28]
  wire [31:0] _GEN_1197 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1150; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2567:29]
  wire [31:0] _GEN_1198 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1151; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2568:28]
  wire [31:0] _GEN_1199 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1152; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2569:29]
  wire [31:0] _GEN_1200 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1153; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2570:28]
  wire [31:0] _GEN_1201 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1154; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2571:29]
  wire [31:0] _GEN_1202 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1155; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2572:28]
  wire [31:0] _GEN_1203 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1156; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2573:29]
  wire [31:0] _GEN_1204 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1157; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2574:28]
  wire [31:0] _GEN_1205 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1158; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2575:29]
  wire [31:0] _GEN_1206 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1159; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2576:28]
  wire [31:0] _GEN_1207 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1160; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2577:29]
  wire [31:0] _GEN_1208 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1161; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2578:28]
  wire [31:0] _GEN_1209 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1162; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2579:29]
  wire [31:0] _GEN_1210 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1163; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2580:29]
  wire [31:0] _GEN_1211 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1164; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2581:29]
  wire [31:0] _GEN_1212 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1165; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2582:28]
  wire [31:0] _GEN_1213 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1166; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2583:29]
  wire [31:0] _GEN_1214 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1167; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2584:28]
  wire [31:0] _GEN_1215 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1168; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2585:29]
  wire [31:0] _GEN_1216 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1169; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2586:28]
  wire [31:0] _GEN_1217 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1170; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2587:29]
  wire [31:0] _GEN_1218 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1171; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2588:28]
  wire [31:0] _GEN_1219 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1172; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2589:29]
  wire [31:0] _GEN_1220 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1173; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2590:28]
  wire [31:0] _GEN_1221 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1174; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2591:29]
  wire [31:0] _GEN_1222 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1175; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2592:28]
  wire [31:0] _GEN_1223 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1176; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2593:29]
  wire [31:0] _GEN_1224 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1177; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2594:28]
  wire [31:0] _GEN_1225 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1178; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2595:29]
  wire [31:0] _GEN_1226 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1179; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2596:28]
  wire [31:0] _GEN_1227 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1180; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2597:29]
  wire [31:0] _GEN_1228 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1181; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2598:28]
  wire [31:0] _GEN_1229 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1182; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2599:29]
  wire [31:0] _GEN_1230 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1183; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2600:29]
  wire [31:0] _GEN_1231 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1184; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2601:29]
  wire [31:0] _GEN_1232 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1185; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2602:28]
  wire [31:0] _GEN_1233 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1186; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2603:29]
  wire [31:0] _GEN_1234 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1187; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2604:28]
  wire [31:0] _GEN_1235 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1188; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2605:29]
  wire [31:0] _GEN_1236 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1189; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2606:28]
  wire [31:0] _GEN_1237 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1190; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2607:29]
  wire [31:0] _GEN_1238 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1191; // @[stackmanage_35.scala 2538:69 stackmanage_35.scala 2608:28]
  wire [31:0] _GEN_1239 = _T_105 & LUT_stack_io_pop_11 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2468:29]
  wire [31:0] _GEN_1240 = _T_105 & LUT_stack_io_pop_11 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2469:28]
  wire [31:0] _GEN_1242 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1192; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2492:29]
  wire [31:0] _GEN_1243 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1193; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2493:28]
  wire [31:0] _GEN_1244 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1195; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2494:29]
  wire [31:0] _GEN_1245 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1196; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2495:28]
  wire [31:0] _GEN_1246 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1197; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2496:29]
  wire [31:0] _GEN_1247 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1198; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2497:28]
  wire [31:0] _GEN_1248 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1199; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2498:29]
  wire [31:0] _GEN_1249 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1200; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2499:28]
  wire [31:0] _GEN_1250 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1201; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2500:29]
  wire [31:0] _GEN_1251 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1202; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2501:28]
  wire [31:0] _GEN_1252 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1203; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2502:29]
  wire [31:0] _GEN_1253 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1204; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2503:28]
  wire [31:0] _GEN_1254 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1205; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2504:29]
  wire [31:0] _GEN_1255 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1206; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2505:28]
  wire [31:0] _GEN_1256 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1207; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2506:29]
  wire [31:0] _GEN_1257 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1208; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2507:28]
  wire [31:0] _GEN_1258 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1209; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2508:29]
  wire [31:0] _GEN_1259 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1210; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2509:29]
  wire [31:0] _GEN_1260 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1211; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2510:29]
  wire [31:0] _GEN_1261 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1212; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2511:28]
  wire [31:0] _GEN_1262 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1213; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2512:29]
  wire [31:0] _GEN_1263 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1214; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2513:28]
  wire [31:0] _GEN_1264 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1215; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2514:29]
  wire [31:0] _GEN_1265 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1216; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2515:28]
  wire [31:0] _GEN_1266 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1217; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2516:29]
  wire [31:0] _GEN_1267 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1218; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2517:28]
  wire [31:0] _GEN_1268 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1219; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2518:29]
  wire [31:0] _GEN_1269 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1220; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2519:28]
  wire [31:0] _GEN_1270 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1221; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2520:29]
  wire [31:0] _GEN_1271 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1222; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2521:28]
  wire [31:0] _GEN_1272 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1223; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2522:29]
  wire [31:0] _GEN_1273 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1224; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2523:28]
  wire [31:0] _GEN_1274 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1225; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2524:29]
  wire [31:0] _GEN_1275 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1226; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2525:28]
  wire [31:0] _GEN_1276 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1227; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2526:29]
  wire [31:0] _GEN_1277 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1228; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2527:28]
  wire [31:0] _GEN_1278 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1229; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2528:29]
  wire [31:0] _GEN_1279 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1230; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2529:29]
  wire [31:0] _GEN_1280 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1231; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2530:29]
  wire [31:0] _GEN_1281 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1232; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2531:28]
  wire [31:0] _GEN_1282 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1233; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2532:29]
  wire [31:0] _GEN_1283 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1234; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2533:28]
  wire [31:0] _GEN_1284 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1235; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2534:29]
  wire [31:0] _GEN_1285 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1236; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2535:28]
  wire [31:0] _GEN_1286 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1237; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2536:29]
  wire [31:0] _GEN_1287 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1238; // @[stackmanage_35.scala 2467:69 stackmanage_35.scala 2537:28]
  wire [31:0] _GEN_1288 = _T_105 & LUT_stack_io_pop_10 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2397:29]
  wire [31:0] _GEN_1289 = _T_105 & LUT_stack_io_pop_10 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2398:28]
  wire [31:0] _GEN_1291 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1239; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2419:29]
  wire [31:0] _GEN_1292 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1240; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2420:28]
  wire [31:0] _GEN_1293 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1242; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2421:29]
  wire [31:0] _GEN_1294 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1243; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2422:28]
  wire [31:0] _GEN_1295 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1244; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2423:29]
  wire [31:0] _GEN_1296 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1245; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2424:28]
  wire [31:0] _GEN_1297 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1246; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2425:29]
  wire [31:0] _GEN_1298 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1247; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2426:28]
  wire [31:0] _GEN_1299 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1248; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2427:29]
  wire [31:0] _GEN_1300 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1249; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2428:28]
  wire [31:0] _GEN_1301 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1250; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2429:29]
  wire [31:0] _GEN_1302 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1251; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2430:28]
  wire [31:0] _GEN_1303 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1252; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2431:29]
  wire [31:0] _GEN_1304 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1253; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2432:28]
  wire [31:0] _GEN_1305 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1254; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2433:29]
  wire [31:0] _GEN_1306 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1255; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2434:28]
  wire [31:0] _GEN_1307 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1256; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2435:29]
  wire [31:0] _GEN_1308 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1257; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2436:28]
  wire [31:0] _GEN_1309 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1258; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2437:29]
  wire [31:0] _GEN_1310 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1259; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2438:29]
  wire [31:0] _GEN_1311 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1260; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2439:29]
  wire [31:0] _GEN_1312 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1261; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2440:28]
  wire [31:0] _GEN_1313 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1262; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2441:29]
  wire [31:0] _GEN_1314 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1263; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2442:28]
  wire [31:0] _GEN_1315 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1264; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2443:29]
  wire [31:0] _GEN_1316 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1265; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2444:28]
  wire [31:0] _GEN_1317 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1266; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2445:29]
  wire [31:0] _GEN_1318 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1267; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2446:28]
  wire [31:0] _GEN_1319 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1268; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2447:29]
  wire [31:0] _GEN_1320 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1269; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2448:28]
  wire [31:0] _GEN_1321 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1270; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2449:29]
  wire [31:0] _GEN_1322 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1271; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2450:28]
  wire [31:0] _GEN_1323 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1272; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2451:29]
  wire [31:0] _GEN_1324 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1273; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2452:28]
  wire [31:0] _GEN_1325 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1274; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2453:29]
  wire [31:0] _GEN_1326 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1275; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2454:28]
  wire [31:0] _GEN_1327 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1276; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2455:29]
  wire [31:0] _GEN_1328 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1277; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2456:28]
  wire [31:0] _GEN_1329 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1278; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2457:29]
  wire [31:0] _GEN_1330 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1279; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2458:29]
  wire [31:0] _GEN_1331 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1280; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2459:29]
  wire [31:0] _GEN_1332 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1281; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2460:28]
  wire [31:0] _GEN_1333 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1282; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2461:29]
  wire [31:0] _GEN_1334 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1283; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2462:28]
  wire [31:0] _GEN_1335 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1284; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2463:29]
  wire [31:0] _GEN_1336 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1285; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2464:28]
  wire [31:0] _GEN_1337 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1286; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2465:29]
  wire [31:0] _GEN_1338 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1287; // @[stackmanage_35.scala 2396:69 stackmanage_35.scala 2466:28]
  wire [31:0] _GEN_1339 = _T_105 & LUT_stack_io_pop_9 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2326:28]
  wire [31:0] _GEN_1340 = _T_105 & LUT_stack_io_pop_9 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2327:27]
  wire [31:0] _GEN_1342 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1288; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2346:29]
  wire [31:0] _GEN_1343 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1289; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2347:29]
  wire [31:0] _GEN_1344 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1291; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2348:29]
  wire [31:0] _GEN_1345 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1292; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2349:28]
  wire [31:0] _GEN_1346 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1293; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2350:29]
  wire [31:0] _GEN_1347 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1294; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2351:28]
  wire [31:0] _GEN_1348 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1295; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2352:29]
  wire [31:0] _GEN_1349 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1296; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2353:28]
  wire [31:0] _GEN_1350 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1297; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2354:29]
  wire [31:0] _GEN_1351 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1298; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2355:28]
  wire [31:0] _GEN_1352 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1299; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2356:29]
  wire [31:0] _GEN_1353 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1300; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2357:28]
  wire [31:0] _GEN_1354 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1301; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2358:29]
  wire [31:0] _GEN_1355 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1302; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2359:28]
  wire [31:0] _GEN_1356 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1303; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2360:29]
  wire [31:0] _GEN_1357 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1304; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2361:28]
  wire [31:0] _GEN_1358 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1305; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2362:29]
  wire [31:0] _GEN_1359 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1306; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2363:28]
  wire [31:0] _GEN_1360 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1307; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2364:29]
  wire [31:0] _GEN_1361 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1308; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2365:28]
  wire [31:0] _GEN_1362 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1309; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2366:29]
  wire [31:0] _GEN_1363 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1310; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2367:29]
  wire [31:0] _GEN_1364 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1311; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2368:29]
  wire [31:0] _GEN_1365 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1312; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2369:28]
  wire [31:0] _GEN_1366 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1313; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2370:29]
  wire [31:0] _GEN_1367 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1314; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2371:28]
  wire [31:0] _GEN_1368 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1315; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2372:29]
  wire [31:0] _GEN_1369 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1316; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2373:28]
  wire [31:0] _GEN_1370 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1317; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2374:29]
  wire [31:0] _GEN_1371 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1318; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2375:28]
  wire [31:0] _GEN_1372 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1319; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2376:29]
  wire [31:0] _GEN_1373 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1320; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2377:28]
  wire [31:0] _GEN_1374 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1321; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2378:29]
  wire [31:0] _GEN_1375 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1322; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2379:28]
  wire [31:0] _GEN_1376 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1323; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2380:29]
  wire [31:0] _GEN_1377 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1324; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2381:28]
  wire [31:0] _GEN_1378 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1325; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2382:29]
  wire [31:0] _GEN_1379 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1326; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2383:28]
  wire [31:0] _GEN_1380 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1327; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2384:29]
  wire [31:0] _GEN_1381 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1328; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2385:28]
  wire [31:0] _GEN_1382 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1329; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2386:29]
  wire [31:0] _GEN_1383 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1330; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2387:29]
  wire [31:0] _GEN_1384 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1331; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2388:29]
  wire [31:0] _GEN_1385 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1332; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2389:28]
  wire [31:0] _GEN_1386 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1333; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2390:29]
  wire [31:0] _GEN_1387 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1334; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2391:28]
  wire [31:0] _GEN_1388 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1335; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2392:29]
  wire [31:0] _GEN_1389 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1336; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2393:28]
  wire [31:0] _GEN_1390 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1337; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2394:29]
  wire [31:0] _GEN_1391 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1338; // @[stackmanage_35.scala 2325:68 stackmanage_35.scala 2395:28]
  wire [31:0] _GEN_1392 = _T_105 & LUT_stack_io_pop_8 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2255:28]
  wire [31:0] _GEN_1393 = _T_105 & LUT_stack_io_pop_8 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2256:27]
  wire [31:0] _GEN_1395 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1339; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2273:28]
  wire [31:0] _GEN_1396 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1340; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2274:27]
  wire [31:0] _GEN_1397 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1342; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2275:29]
  wire [31:0] _GEN_1398 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1343; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2276:29]
  wire [31:0] _GEN_1399 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1344; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2277:29]
  wire [31:0] _GEN_1400 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1345; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2278:28]
  wire [31:0] _GEN_1401 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1346; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2279:29]
  wire [31:0] _GEN_1402 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1347; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2280:28]
  wire [31:0] _GEN_1403 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1348; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2281:29]
  wire [31:0] _GEN_1404 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1349; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2282:28]
  wire [31:0] _GEN_1405 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1350; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2283:29]
  wire [31:0] _GEN_1406 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1351; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2284:28]
  wire [31:0] _GEN_1407 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1352; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2285:29]
  wire [31:0] _GEN_1408 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1353; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2286:28]
  wire [31:0] _GEN_1409 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1354; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2287:29]
  wire [31:0] _GEN_1410 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1355; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2288:28]
  wire [31:0] _GEN_1411 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1356; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2289:29]
  wire [31:0] _GEN_1412 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1357; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2290:28]
  wire [31:0] _GEN_1413 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1358; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2291:29]
  wire [31:0] _GEN_1414 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1359; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2292:28]
  wire [31:0] _GEN_1415 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1360; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2293:29]
  wire [31:0] _GEN_1416 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1361; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2294:28]
  wire [31:0] _GEN_1417 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1362; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2295:29]
  wire [31:0] _GEN_1418 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1363; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2296:29]
  wire [31:0] _GEN_1419 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1364; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2297:29]
  wire [31:0] _GEN_1420 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1365; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2298:28]
  wire [31:0] _GEN_1421 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1366; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2299:29]
  wire [31:0] _GEN_1422 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1367; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2300:28]
  wire [31:0] _GEN_1423 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1368; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2301:29]
  wire [31:0] _GEN_1424 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1369; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2302:28]
  wire [31:0] _GEN_1425 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1370; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2303:29]
  wire [31:0] _GEN_1426 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1371; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2304:28]
  wire [31:0] _GEN_1427 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1372; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2305:29]
  wire [31:0] _GEN_1428 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1373; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2306:28]
  wire [31:0] _GEN_1429 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1374; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2307:29]
  wire [31:0] _GEN_1430 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1375; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2308:28]
  wire [31:0] _GEN_1431 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1376; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2309:29]
  wire [31:0] _GEN_1432 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1377; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2310:28]
  wire [31:0] _GEN_1433 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1378; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2311:29]
  wire [31:0] _GEN_1434 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1379; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2312:28]
  wire [31:0] _GEN_1435 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1380; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2313:29]
  wire [31:0] _GEN_1436 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1381; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2314:28]
  wire [31:0] _GEN_1437 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1382; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2315:29]
  wire [31:0] _GEN_1438 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1383; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2316:29]
  wire [31:0] _GEN_1439 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1384; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2317:29]
  wire [31:0] _GEN_1440 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1385; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2318:28]
  wire [31:0] _GEN_1441 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1386; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2319:29]
  wire [31:0] _GEN_1442 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1387; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2320:28]
  wire [31:0] _GEN_1443 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1388; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2321:29]
  wire [31:0] _GEN_1444 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1389; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2322:28]
  wire [31:0] _GEN_1445 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1390; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2323:29]
  wire [31:0] _GEN_1446 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1391; // @[stackmanage_35.scala 2254:68 stackmanage_35.scala 2324:28]
  wire [31:0] _GEN_1447 = _T_105 & LUT_stack_io_pop_7 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2184:28]
  wire [31:0] _GEN_1448 = _T_105 & LUT_stack_io_pop_7 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2185:27]
  wire [31:0] _GEN_1450 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1392; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2200:28]
  wire [31:0] _GEN_1451 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1393; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2201:27]
  wire [31:0] _GEN_1452 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1395; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2202:28]
  wire [31:0] _GEN_1453 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1396; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2203:27]
  wire [31:0] _GEN_1454 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1397; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2204:29]
  wire [31:0] _GEN_1455 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1398; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2205:29]
  wire [31:0] _GEN_1456 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1399; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2206:29]
  wire [31:0] _GEN_1457 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1400; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2207:28]
  wire [31:0] _GEN_1458 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1401; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2208:29]
  wire [31:0] _GEN_1459 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1402; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2209:28]
  wire [31:0] _GEN_1460 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1403; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2210:29]
  wire [31:0] _GEN_1461 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1404; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2211:28]
  wire [31:0] _GEN_1462 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1405; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2212:29]
  wire [31:0] _GEN_1463 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1406; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2213:28]
  wire [31:0] _GEN_1464 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1407; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2214:29]
  wire [31:0] _GEN_1465 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1408; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2215:28]
  wire [31:0] _GEN_1466 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1409; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2216:29]
  wire [31:0] _GEN_1467 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1410; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2217:28]
  wire [31:0] _GEN_1468 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1411; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2218:29]
  wire [31:0] _GEN_1469 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1412; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2219:28]
  wire [31:0] _GEN_1470 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1413; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2220:29]
  wire [31:0] _GEN_1471 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1414; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2221:28]
  wire [31:0] _GEN_1472 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1415; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2222:29]
  wire [31:0] _GEN_1473 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1416; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2223:28]
  wire [31:0] _GEN_1474 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1417; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2224:29]
  wire [31:0] _GEN_1475 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1418; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2225:29]
  wire [31:0] _GEN_1476 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1419; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2226:29]
  wire [31:0] _GEN_1477 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1420; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2227:28]
  wire [31:0] _GEN_1478 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1421; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2228:29]
  wire [31:0] _GEN_1479 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1422; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2229:28]
  wire [31:0] _GEN_1480 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1423; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2230:29]
  wire [31:0] _GEN_1481 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1424; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2231:28]
  wire [31:0] _GEN_1482 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1425; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2232:29]
  wire [31:0] _GEN_1483 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1426; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2233:28]
  wire [31:0] _GEN_1484 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1427; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2234:29]
  wire [31:0] _GEN_1485 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1428; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2235:28]
  wire [31:0] _GEN_1486 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1429; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2236:29]
  wire [31:0] _GEN_1487 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1430; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2237:28]
  wire [31:0] _GEN_1488 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1431; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2238:29]
  wire [31:0] _GEN_1489 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1432; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2239:28]
  wire [31:0] _GEN_1490 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1433; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2240:29]
  wire [31:0] _GEN_1491 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1434; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2241:28]
  wire [31:0] _GEN_1492 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1435; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2242:29]
  wire [31:0] _GEN_1493 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1436; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2243:28]
  wire [31:0] _GEN_1494 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1437; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2244:29]
  wire [31:0] _GEN_1495 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1438; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2245:29]
  wire [31:0] _GEN_1496 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1439; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2246:29]
  wire [31:0] _GEN_1497 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1440; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2247:28]
  wire [31:0] _GEN_1498 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1441; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2248:29]
  wire [31:0] _GEN_1499 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1442; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2249:28]
  wire [31:0] _GEN_1500 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1443; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2250:29]
  wire [31:0] _GEN_1501 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1444; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2251:28]
  wire [31:0] _GEN_1502 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1445; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2252:29]
  wire [31:0] _GEN_1503 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1446; // @[stackmanage_35.scala 2183:68 stackmanage_35.scala 2253:28]
  wire [31:0] _GEN_1504 = _T_105 & LUT_stack_io_pop_6 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2113:28]
  wire [31:0] _GEN_1505 = _T_105 & LUT_stack_io_pop_6 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2114:27]
  wire [31:0] _GEN_1507 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1447; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2127:28]
  wire [31:0] _GEN_1508 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1448; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2128:27]
  wire [31:0] _GEN_1509 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1450; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2129:28]
  wire [31:0] _GEN_1510 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1451; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2130:27]
  wire [31:0] _GEN_1511 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1452; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2131:28]
  wire [31:0] _GEN_1512 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1453; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2132:27]
  wire [31:0] _GEN_1513 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1454; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2133:29]
  wire [31:0] _GEN_1514 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1455; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2134:29]
  wire [31:0] _GEN_1515 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1456; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2135:29]
  wire [31:0] _GEN_1516 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1457; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2136:28]
  wire [31:0] _GEN_1517 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1458; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2137:29]
  wire [31:0] _GEN_1518 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1459; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2138:28]
  wire [31:0] _GEN_1519 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1460; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2139:29]
  wire [31:0] _GEN_1520 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1461; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2140:28]
  wire [31:0] _GEN_1521 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1462; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2141:29]
  wire [31:0] _GEN_1522 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1463; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2142:28]
  wire [31:0] _GEN_1523 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1464; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2143:29]
  wire [31:0] _GEN_1524 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1465; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2144:28]
  wire [31:0] _GEN_1525 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1466; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2145:29]
  wire [31:0] _GEN_1526 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1467; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2146:28]
  wire [31:0] _GEN_1527 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1468; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2147:29]
  wire [31:0] _GEN_1528 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1469; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2148:28]
  wire [31:0] _GEN_1529 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1470; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2149:29]
  wire [31:0] _GEN_1530 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1471; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2150:28]
  wire [31:0] _GEN_1531 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1472; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2151:29]
  wire [31:0] _GEN_1532 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1473; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2152:28]
  wire [31:0] _GEN_1533 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1474; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2153:29]
  wire [31:0] _GEN_1534 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1475; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2154:29]
  wire [31:0] _GEN_1535 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1476; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2155:29]
  wire [31:0] _GEN_1536 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1477; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2156:28]
  wire [31:0] _GEN_1537 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1478; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2157:29]
  wire [31:0] _GEN_1538 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1479; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2158:28]
  wire [31:0] _GEN_1539 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1480; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2159:29]
  wire [31:0] _GEN_1540 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1481; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2160:28]
  wire [31:0] _GEN_1541 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1482; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2161:29]
  wire [31:0] _GEN_1542 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1483; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2162:28]
  wire [31:0] _GEN_1543 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1484; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2163:29]
  wire [31:0] _GEN_1544 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1485; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2164:28]
  wire [31:0] _GEN_1545 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1486; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2165:29]
  wire [31:0] _GEN_1546 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1487; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2166:28]
  wire [31:0] _GEN_1547 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1488; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2167:29]
  wire [31:0] _GEN_1548 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1489; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2168:28]
  wire [31:0] _GEN_1549 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1490; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2169:29]
  wire [31:0] _GEN_1550 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1491; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2170:28]
  wire [31:0] _GEN_1551 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1492; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2171:29]
  wire [31:0] _GEN_1552 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1493; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2172:28]
  wire [31:0] _GEN_1553 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1494; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2173:29]
  wire [31:0] _GEN_1554 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1495; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2174:29]
  wire [31:0] _GEN_1555 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1496; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2175:29]
  wire [31:0] _GEN_1556 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1497; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2176:28]
  wire [31:0] _GEN_1557 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1498; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2177:29]
  wire [31:0] _GEN_1558 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1499; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2178:28]
  wire [31:0] _GEN_1559 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1500; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2179:29]
  wire [31:0] _GEN_1560 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1501; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2180:28]
  wire [31:0] _GEN_1561 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1502; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2181:29]
  wire [31:0] _GEN_1562 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1503; // @[stackmanage_35.scala 2112:68 stackmanage_35.scala 2182:28]
  wire [31:0] _GEN_1563 = _T_105 & LUT_stack_io_pop_5 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2042:28]
  wire [31:0] _GEN_1564 = _T_105 & LUT_stack_io_pop_5 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2043:27]
  wire [31:0] _GEN_1566 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1504; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2054:28]
  wire [31:0] _GEN_1567 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1505; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2055:27]
  wire [31:0] _GEN_1568 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1507; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2056:28]
  wire [31:0] _GEN_1569 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1508; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2057:27]
  wire [31:0] _GEN_1570 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1509; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2058:28]
  wire [31:0] _GEN_1571 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1510; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2059:27]
  wire [31:0] _GEN_1572 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1511; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2060:28]
  wire [31:0] _GEN_1573 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1512; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2061:27]
  wire [31:0] _GEN_1574 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1513; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2062:29]
  wire [31:0] _GEN_1575 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1514; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2063:29]
  wire [31:0] _GEN_1576 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1515; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2064:29]
  wire [31:0] _GEN_1577 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1516; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2065:28]
  wire [31:0] _GEN_1578 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1517; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2066:29]
  wire [31:0] _GEN_1579 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1518; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2067:28]
  wire [31:0] _GEN_1580 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1519; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2068:29]
  wire [31:0] _GEN_1581 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1520; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2069:28]
  wire [31:0] _GEN_1582 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1521; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2070:29]
  wire [31:0] _GEN_1583 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1522; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2071:28]
  wire [31:0] _GEN_1584 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1523; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2072:29]
  wire [31:0] _GEN_1585 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1524; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2073:28]
  wire [31:0] _GEN_1586 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1525; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2074:29]
  wire [31:0] _GEN_1587 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1526; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2075:28]
  wire [31:0] _GEN_1588 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1527; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2076:29]
  wire [31:0] _GEN_1589 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1528; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2077:28]
  wire [31:0] _GEN_1590 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1529; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2078:29]
  wire [31:0] _GEN_1591 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1530; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2079:28]
  wire [31:0] _GEN_1592 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1531; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2080:29]
  wire [31:0] _GEN_1593 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1532; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2081:28]
  wire [31:0] _GEN_1594 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1533; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2082:29]
  wire [31:0] _GEN_1595 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1534; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2083:29]
  wire [31:0] _GEN_1596 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1535; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2084:29]
  wire [31:0] _GEN_1597 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1536; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2085:28]
  wire [31:0] _GEN_1598 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1537; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2086:29]
  wire [31:0] _GEN_1599 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1538; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2087:28]
  wire [31:0] _GEN_1600 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1539; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2088:29]
  wire [31:0] _GEN_1601 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1540; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2089:28]
  wire [31:0] _GEN_1602 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1541; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2090:29]
  wire [31:0] _GEN_1603 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1542; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2091:28]
  wire [31:0] _GEN_1604 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1543; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2092:29]
  wire [31:0] _GEN_1605 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1544; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2093:28]
  wire [31:0] _GEN_1606 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1545; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2094:29]
  wire [31:0] _GEN_1607 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1546; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2095:28]
  wire [31:0] _GEN_1608 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1547; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2096:29]
  wire [31:0] _GEN_1609 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1548; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2097:28]
  wire [31:0] _GEN_1610 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1549; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2098:29]
  wire [31:0] _GEN_1611 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1550; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2099:28]
  wire [31:0] _GEN_1612 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1551; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2100:29]
  wire [31:0] _GEN_1613 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1552; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2101:28]
  wire [31:0] _GEN_1614 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1553; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2102:29]
  wire [31:0] _GEN_1615 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1554; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2103:29]
  wire [31:0] _GEN_1616 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1555; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2104:29]
  wire [31:0] _GEN_1617 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1556; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2105:28]
  wire [31:0] _GEN_1618 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1557; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2106:29]
  wire [31:0] _GEN_1619 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1558; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2107:28]
  wire [31:0] _GEN_1620 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1559; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2108:29]
  wire [31:0] _GEN_1621 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1560; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2109:28]
  wire [31:0] _GEN_1622 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1561; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2110:29]
  wire [31:0] _GEN_1623 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1562; // @[stackmanage_35.scala 2041:68 stackmanage_35.scala 2111:28]
  wire [31:0] _GEN_1624 = _T_105 & LUT_stack_io_pop_4 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 1971:28]
  wire [31:0] _GEN_1625 = _T_105 & LUT_stack_io_pop_4 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 1972:27]
  wire [31:0] _GEN_1627 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1563; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 1981:28]
  wire [31:0] _GEN_1628 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1564; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 1982:27]
  wire [31:0] _GEN_1629 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1566; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 1983:28]
  wire [31:0] _GEN_1630 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1567; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 1984:27]
  wire [31:0] _GEN_1631 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1568; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 1985:28]
  wire [31:0] _GEN_1632 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1569; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 1986:27]
  wire [31:0] _GEN_1633 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1570; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 1987:28]
  wire [31:0] _GEN_1634 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1571; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 1988:27]
  wire [31:0] _GEN_1635 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1572; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 1989:28]
  wire [31:0] _GEN_1636 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1573; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 1990:27]
  wire [31:0] _GEN_1637 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1574; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 1991:29]
  wire [31:0] _GEN_1638 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1575; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 1992:29]
  wire [31:0] _GEN_1639 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1576; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 1993:29]
  wire [31:0] _GEN_1640 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1577; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 1994:28]
  wire [31:0] _GEN_1641 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1578; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 1995:29]
  wire [31:0] _GEN_1642 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1579; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 1996:28]
  wire [31:0] _GEN_1643 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1580; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 1997:29]
  wire [31:0] _GEN_1644 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1581; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 1998:28]
  wire [31:0] _GEN_1645 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1582; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 1999:29]
  wire [31:0] _GEN_1646 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1583; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 2000:28]
  wire [31:0] _GEN_1647 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1584; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 2001:29]
  wire [31:0] _GEN_1648 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1585; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 2002:28]
  wire [31:0] _GEN_1649 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1586; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 2003:29]
  wire [31:0] _GEN_1650 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1587; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 2004:28]
  wire [31:0] _GEN_1651 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1588; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 2005:29]
  wire [31:0] _GEN_1652 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1589; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 2006:28]
  wire [31:0] _GEN_1653 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1590; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 2007:29]
  wire [31:0] _GEN_1654 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1591; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 2008:28]
  wire [31:0] _GEN_1655 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1592; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 2009:29]
  wire [31:0] _GEN_1656 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1593; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 2010:28]
  wire [31:0] _GEN_1657 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1594; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 2011:29]
  wire [31:0] _GEN_1658 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1595; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 2012:29]
  wire [31:0] _GEN_1659 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1596; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 2013:29]
  wire [31:0] _GEN_1660 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1597; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 2014:28]
  wire [31:0] _GEN_1661 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1598; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 2015:29]
  wire [31:0] _GEN_1662 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1599; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 2016:28]
  wire [31:0] _GEN_1663 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1600; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 2017:29]
  wire [31:0] _GEN_1664 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1601; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 2018:28]
  wire [31:0] _GEN_1665 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1602; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 2019:29]
  wire [31:0] _GEN_1666 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1603; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 2020:28]
  wire [31:0] _GEN_1667 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1604; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 2021:29]
  wire [31:0] _GEN_1668 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1605; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 2022:28]
  wire [31:0] _GEN_1669 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1606; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 2023:29]
  wire [31:0] _GEN_1670 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1607; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 2024:28]
  wire [31:0] _GEN_1671 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1608; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 2025:29]
  wire [31:0] _GEN_1672 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1609; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 2026:28]
  wire [31:0] _GEN_1673 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1610; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 2027:29]
  wire [31:0] _GEN_1674 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1611; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 2028:28]
  wire [31:0] _GEN_1675 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1612; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 2029:29]
  wire [31:0] _GEN_1676 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1613; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 2030:28]
  wire [31:0] _GEN_1677 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1614; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 2031:29]
  wire [31:0] _GEN_1678 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1615; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 2032:29]
  wire [31:0] _GEN_1679 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1616; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 2033:29]
  wire [31:0] _GEN_1680 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1617; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 2034:28]
  wire [31:0] _GEN_1681 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1618; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 2035:29]
  wire [31:0] _GEN_1682 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1619; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 2036:28]
  wire [31:0] _GEN_1683 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1620; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 2037:29]
  wire [31:0] _GEN_1684 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1621; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 2038:28]
  wire [31:0] _GEN_1685 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1622; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 2039:29]
  wire [31:0] _GEN_1686 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1623; // @[stackmanage_35.scala 1970:68 stackmanage_35.scala 2040:28]
  wire [31:0] _GEN_1687 = _T_105 & LUT_stack_io_pop_3 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1900:28]
  wire [31:0] _GEN_1688 = _T_105 & LUT_stack_io_pop_3 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1901:27]
  wire [31:0] _GEN_1690 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1624; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1908:28]
  wire [31:0] _GEN_1691 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1625; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1909:27]
  wire [31:0] _GEN_1692 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1627; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1910:28]
  wire [31:0] _GEN_1693 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1628; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1911:27]
  wire [31:0] _GEN_1694 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1629; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1912:28]
  wire [31:0] _GEN_1695 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1630; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1913:27]
  wire [31:0] _GEN_1696 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1631; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1914:28]
  wire [31:0] _GEN_1697 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1632; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1915:27]
  wire [31:0] _GEN_1698 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1633; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1916:28]
  wire [31:0] _GEN_1699 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1634; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1917:27]
  wire [31:0] _GEN_1700 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1635; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1918:28]
  wire [31:0] _GEN_1701 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1636; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1919:27]
  wire [31:0] _GEN_1702 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1637; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1920:29]
  wire [31:0] _GEN_1703 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1638; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1921:29]
  wire [31:0] _GEN_1704 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1639; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1922:29]
  wire [31:0] _GEN_1705 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1640; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1923:28]
  wire [31:0] _GEN_1706 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1641; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1924:29]
  wire [31:0] _GEN_1707 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1642; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1925:28]
  wire [31:0] _GEN_1708 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1643; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1926:29]
  wire [31:0] _GEN_1709 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1644; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1927:28]
  wire [31:0] _GEN_1710 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1645; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1928:29]
  wire [31:0] _GEN_1711 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1646; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1929:28]
  wire [31:0] _GEN_1712 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1647; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1930:29]
  wire [31:0] _GEN_1713 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1648; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1931:28]
  wire [31:0] _GEN_1714 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1649; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1932:29]
  wire [31:0] _GEN_1715 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1650; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1933:28]
  wire [31:0] _GEN_1716 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1651; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1934:29]
  wire [31:0] _GEN_1717 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1652; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1935:28]
  wire [31:0] _GEN_1718 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1653; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1936:29]
  wire [31:0] _GEN_1719 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1654; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1937:28]
  wire [31:0] _GEN_1720 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1655; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1938:29]
  wire [31:0] _GEN_1721 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1656; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1939:28]
  wire [31:0] _GEN_1722 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1657; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1940:29]
  wire [31:0] _GEN_1723 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1658; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1941:29]
  wire [31:0] _GEN_1724 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1659; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1942:29]
  wire [31:0] _GEN_1725 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1660; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1943:28]
  wire [31:0] _GEN_1726 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1661; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1944:29]
  wire [31:0] _GEN_1727 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1662; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1945:28]
  wire [31:0] _GEN_1728 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1663; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1946:29]
  wire [31:0] _GEN_1729 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1664; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1947:28]
  wire [31:0] _GEN_1730 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1665; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1948:29]
  wire [31:0] _GEN_1731 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1666; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1949:28]
  wire [31:0] _GEN_1732 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1667; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1950:29]
  wire [31:0] _GEN_1733 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1668; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1951:28]
  wire [31:0] _GEN_1734 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1669; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1952:29]
  wire [31:0] _GEN_1735 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1670; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1953:28]
  wire [31:0] _GEN_1736 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1671; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1954:29]
  wire [31:0] _GEN_1737 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1672; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1955:28]
  wire [31:0] _GEN_1738 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1673; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1956:29]
  wire [31:0] _GEN_1739 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1674; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1957:28]
  wire [31:0] _GEN_1740 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1675; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1958:29]
  wire [31:0] _GEN_1741 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1676; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1959:28]
  wire [31:0] _GEN_1742 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1677; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1960:29]
  wire [31:0] _GEN_1743 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1678; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1961:29]
  wire [31:0] _GEN_1744 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1679; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1962:29]
  wire [31:0] _GEN_1745 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1680; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1963:28]
  wire [31:0] _GEN_1746 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1681; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1964:29]
  wire [31:0] _GEN_1747 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1682; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1965:28]
  wire [31:0] _GEN_1748 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1683; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1966:29]
  wire [31:0] _GEN_1749 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1684; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1967:28]
  wire [31:0] _GEN_1750 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1685; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1968:29]
  wire [31:0] _GEN_1751 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1686; // @[stackmanage_35.scala 1899:68 stackmanage_35.scala 1969:28]
  wire [31:0] _GEN_1752 = _T_105 & LUT_stack_io_pop_2 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1829:28]
  wire [31:0] _GEN_1753 = _T_105 & LUT_stack_io_pop_2 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1830:27]
  wire [31:0] _GEN_1755 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1687; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1835:28]
  wire [31:0] _GEN_1756 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1688; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1836:27]
  wire [31:0] _GEN_1757 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1690; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1837:28]
  wire [31:0] _GEN_1758 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1691; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1838:27]
  wire [31:0] _GEN_1759 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1692; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1839:28]
  wire [31:0] _GEN_1760 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1693; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1840:27]
  wire [31:0] _GEN_1761 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1694; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1841:28]
  wire [31:0] _GEN_1762 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1695; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1842:27]
  wire [31:0] _GEN_1763 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1696; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1843:28]
  wire [31:0] _GEN_1764 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1697; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1844:27]
  wire [31:0] _GEN_1765 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1698; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1845:28]
  wire [31:0] _GEN_1766 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1699; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1846:27]
  wire [31:0] _GEN_1767 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1700; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1847:28]
  wire [31:0] _GEN_1768 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1701; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1848:27]
  wire [31:0] _GEN_1769 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1702; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1849:29]
  wire [31:0] _GEN_1770 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1703; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1850:29]
  wire [31:0] _GEN_1771 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1704; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1851:29]
  wire [31:0] _GEN_1772 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1705; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1852:28]
  wire [31:0] _GEN_1773 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1706; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1853:29]
  wire [31:0] _GEN_1774 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1707; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1854:28]
  wire [31:0] _GEN_1775 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1708; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1855:29]
  wire [31:0] _GEN_1776 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1709; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1856:28]
  wire [31:0] _GEN_1777 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1710; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1857:29]
  wire [31:0] _GEN_1778 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1711; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1858:28]
  wire [31:0] _GEN_1779 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1712; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1859:29]
  wire [31:0] _GEN_1780 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1713; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1860:28]
  wire [31:0] _GEN_1781 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1714; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1861:29]
  wire [31:0] _GEN_1782 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1715; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1862:28]
  wire [31:0] _GEN_1783 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1716; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1863:29]
  wire [31:0] _GEN_1784 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1717; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1864:28]
  wire [31:0] _GEN_1785 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1718; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1865:29]
  wire [31:0] _GEN_1786 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1719; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1866:28]
  wire [31:0] _GEN_1787 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1720; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1867:29]
  wire [31:0] _GEN_1788 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1721; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1868:28]
  wire [31:0] _GEN_1789 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1722; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1869:29]
  wire [31:0] _GEN_1790 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1723; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1870:29]
  wire [31:0] _GEN_1791 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1724; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1871:29]
  wire [31:0] _GEN_1792 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1725; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1872:28]
  wire [31:0] _GEN_1793 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1726; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1873:29]
  wire [31:0] _GEN_1794 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1727; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1874:28]
  wire [31:0] _GEN_1795 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1728; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1875:29]
  wire [31:0] _GEN_1796 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1729; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1876:28]
  wire [31:0] _GEN_1797 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1730; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1877:29]
  wire [31:0] _GEN_1798 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1731; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1878:28]
  wire [31:0] _GEN_1799 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1732; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1879:29]
  wire [31:0] _GEN_1800 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1733; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1880:28]
  wire [31:0] _GEN_1801 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1734; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1881:29]
  wire [31:0] _GEN_1802 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1735; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1882:28]
  wire [31:0] _GEN_1803 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1736; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1883:29]
  wire [31:0] _GEN_1804 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1737; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1884:28]
  wire [31:0] _GEN_1805 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1738; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1885:29]
  wire [31:0] _GEN_1806 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1739; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1886:28]
  wire [31:0] _GEN_1807 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1740; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1887:29]
  wire [31:0] _GEN_1808 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1741; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1888:28]
  wire [31:0] _GEN_1809 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1742; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1889:29]
  wire [31:0] _GEN_1810 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1743; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1890:29]
  wire [31:0] _GEN_1811 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1744; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1891:29]
  wire [31:0] _GEN_1812 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1745; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1892:28]
  wire [31:0] _GEN_1813 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1746; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1893:29]
  wire [31:0] _GEN_1814 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1747; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1894:28]
  wire [31:0] _GEN_1815 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1748; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1895:29]
  wire [31:0] _GEN_1816 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1749; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1896:28]
  wire [31:0] _GEN_1817 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1750; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1897:29]
  wire [31:0] _GEN_1818 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1751; // @[stackmanage_35.scala 1828:68 stackmanage_35.scala 1898:28]
  wire [31:0] _GEN_1819 = _T_105 & LUT_stack_io_pop_1 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1758:28]
  wire [31:0] _GEN_1820 = _T_105 & LUT_stack_io_pop_1 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1759:27]
  wire [31:0] _GEN_1822 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1752; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1762:28]
  wire [31:0] _GEN_1823 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1753; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1763:27]
  wire [31:0] _GEN_1824 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1755; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1764:28]
  wire [31:0] _GEN_1825 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1756; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1765:27]
  wire [31:0] _GEN_1826 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1757; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1766:28]
  wire [31:0] _GEN_1827 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1758; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1767:27]
  wire [31:0] _GEN_1828 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1759; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1768:28]
  wire [31:0] _GEN_1829 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1760; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1769:27]
  wire [31:0] _GEN_1830 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1761; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1770:28]
  wire [31:0] _GEN_1831 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1762; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1771:27]
  wire [31:0] _GEN_1832 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1763; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1772:28]
  wire [31:0] _GEN_1833 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1764; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1773:27]
  wire [31:0] _GEN_1834 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1765; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1774:28]
  wire [31:0] _GEN_1835 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1766; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1775:27]
  wire [31:0] _GEN_1836 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1767; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1776:28]
  wire [31:0] _GEN_1837 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1768; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1777:27]
  wire [31:0] _GEN_1838 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1769; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1778:29]
  wire [31:0] _GEN_1839 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1770; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1779:29]
  wire [31:0] _GEN_1840 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1771; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1780:29]
  wire [31:0] _GEN_1841 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1772; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1781:28]
  wire [31:0] _GEN_1842 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1773; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1782:29]
  wire [31:0] _GEN_1843 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1774; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1783:28]
  wire [31:0] _GEN_1844 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1775; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1784:29]
  wire [31:0] _GEN_1845 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1776; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1785:28]
  wire [31:0] _GEN_1846 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1777; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1786:29]
  wire [31:0] _GEN_1847 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1778; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1787:28]
  wire [31:0] _GEN_1848 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1779; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1788:29]
  wire [31:0] _GEN_1849 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1780; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1789:28]
  wire [31:0] _GEN_1850 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1781; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1790:29]
  wire [31:0] _GEN_1851 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1782; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1791:28]
  wire [31:0] _GEN_1852 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1783; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1792:29]
  wire [31:0] _GEN_1853 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1784; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1793:28]
  wire [31:0] _GEN_1854 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1785; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1794:29]
  wire [31:0] _GEN_1855 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1786; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1795:28]
  wire [31:0] _GEN_1856 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1787; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1796:29]
  wire [31:0] _GEN_1857 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1788; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1797:28]
  wire [31:0] _GEN_1858 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1789; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1798:29]
  wire [31:0] _GEN_1859 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1790; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1799:29]
  wire [31:0] _GEN_1860 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1791; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1800:29]
  wire [31:0] _GEN_1861 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1792; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1801:28]
  wire [31:0] _GEN_1862 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1793; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1802:29]
  wire [31:0] _GEN_1863 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1794; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1803:28]
  wire [31:0] _GEN_1864 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1795; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1804:29]
  wire [31:0] _GEN_1865 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1796; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1805:28]
  wire [31:0] _GEN_1866 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1797; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1806:29]
  wire [31:0] _GEN_1867 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1798; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1807:28]
  wire [31:0] _GEN_1868 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1799; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1808:29]
  wire [31:0] _GEN_1869 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1800; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1809:28]
  wire [31:0] _GEN_1870 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1801; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1810:29]
  wire [31:0] _GEN_1871 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1802; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1811:28]
  wire [31:0] _GEN_1872 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1803; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1812:29]
  wire [31:0] _GEN_1873 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1804; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1813:28]
  wire [31:0] _GEN_1874 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1805; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1814:29]
  wire [31:0] _GEN_1875 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1806; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1815:28]
  wire [31:0] _GEN_1876 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1807; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1816:29]
  wire [31:0] _GEN_1877 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1808; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1817:28]
  wire [31:0] _GEN_1878 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1809; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1818:29]
  wire [31:0] _GEN_1879 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1810; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1819:29]
  wire [31:0] _GEN_1880 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1811; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1820:29]
  wire [31:0] _GEN_1881 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1812; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1821:28]
  wire [31:0] _GEN_1882 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1813; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1822:29]
  wire [31:0] _GEN_1883 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1814; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1823:28]
  wire [31:0] _GEN_1884 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1815; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1824:29]
  wire [31:0] _GEN_1885 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1816; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1825:28]
  wire [31:0] _GEN_1886 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1817; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1826:29]
  wire [31:0] _GEN_1887 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1818; // @[stackmanage_35.scala 1757:68 stackmanage_35.scala 1827:28]
  reg  pop_0; // @[stackmanage_35.scala 4245:46]
  reg  pop_1; // @[stackmanage_35.scala 4246:46]
  reg  pop_2; // @[stackmanage_35.scala 4247:46]
  reg  pop_3; // @[stackmanage_35.scala 4248:46]
  reg  pop_4; // @[stackmanage_35.scala 4249:46]
  reg  pop_5; // @[stackmanage_35.scala 4250:46]
  reg  pop_6; // @[stackmanage_35.scala 4251:46]
  reg  pop_7; // @[stackmanage_35.scala 4252:46]
  reg  pop_8; // @[stackmanage_35.scala 4253:46]
  reg  pop_9; // @[stackmanage_35.scala 4254:46]
  reg  pop_10; // @[stackmanage_35.scala 4256:47]
  reg  pop_11; // @[stackmanage_35.scala 4257:47]
  reg  pop_12; // @[stackmanage_35.scala 4258:47]
  reg  pop_13; // @[stackmanage_35.scala 4259:47]
  reg  pop_14; // @[stackmanage_35.scala 4260:47]
  reg  pop_15; // @[stackmanage_35.scala 4261:47]
  reg  pop_16; // @[stackmanage_35.scala 4262:47]
  reg  pop_17; // @[stackmanage_35.scala 4263:47]
  reg  pop_18; // @[stackmanage_35.scala 4264:47]
  reg  pop_19; // @[stackmanage_35.scala 4265:47]
  reg  pop_20; // @[stackmanage_35.scala 4267:47]
  reg  pop_21; // @[stackmanage_35.scala 4268:47]
  reg  pop_22; // @[stackmanage_35.scala 4269:47]
  reg  pop_23; // @[stackmanage_35.scala 4270:47]
  reg  pop_24; // @[stackmanage_35.scala 4271:47]
  reg  pop_25; // @[stackmanage_35.scala 4272:47]
  reg  pop_26; // @[stackmanage_35.scala 4273:47]
  reg  pop_27; // @[stackmanage_35.scala 4274:47]
  reg  pop_28; // @[stackmanage_35.scala 4275:47]
  reg  pop_29; // @[stackmanage_35.scala 4276:47]
  reg  pop_30; // @[stackmanage_35.scala 4278:47]
  reg  pop_31; // @[stackmanage_35.scala 4279:47]
  reg  pop_32; // @[stackmanage_35.scala 4280:47]
  reg  pop_33; // @[stackmanage_35.scala 4281:47]
  reg  pop_34; // @[stackmanage_35.scala 4282:47]
  wire  _T_314 = pop_34 & Stack_34_io_enable; // @[stackmanage_35.scala 4503:28]
  wire [31:0] _GEN_1958 = pop_34 & Stack_34_io_enable ? Stack_34_io_hit_out : 32'h0; // @[stackmanage_35.scala 4503:55 stackmanage_35.scala 4504:27 stackmanage_35.scala 4510:27]
  wire [31:0] _GEN_1959 = pop_34 & Stack_34_io_enable ? Stack_34_io_ray_out : 32'h0; // @[stackmanage_35.scala 4503:55 stackmanage_35.scala 4505:28 stackmanage_35.scala 4511:28]
  wire [31:0] _GEN_1960 = pop_34 & Stack_34_io_enable ? $signed(Stack_34_io_dataOut) : $signed(32'sh0); // @[stackmanage_35.scala 4503:55 stackmanage_35.scala 4506:25 stackmanage_35.scala 4512:25]
  wire [31:0] _GEN_1962 = pop_33 & Stack_33_io_enable ? Stack_33_io_hit_out : _GEN_1958; // @[stackmanage_35.scala 4498:55 stackmanage_35.scala 4499:27]
  wire [31:0] _GEN_1963 = pop_33 & Stack_33_io_enable ? Stack_33_io_ray_out : _GEN_1959; // @[stackmanage_35.scala 4498:55 stackmanage_35.scala 4500:28]
  wire [31:0] _GEN_1964 = pop_33 & Stack_33_io_enable ? $signed(Stack_33_io_dataOut) : $signed(_GEN_1960); // @[stackmanage_35.scala 4498:55 stackmanage_35.scala 4501:25]
  wire  _GEN_1965 = pop_33 & Stack_33_io_enable | _T_314; // @[stackmanage_35.scala 4498:55 stackmanage_35.scala 4502:31]
  wire [31:0] _GEN_1966 = pop_32 & Stack_32_io_enable ? Stack_32_io_hit_out : _GEN_1962; // @[stackmanage_35.scala 4493:55 stackmanage_35.scala 4494:27]
  wire [31:0] _GEN_1967 = pop_32 & Stack_32_io_enable ? Stack_32_io_ray_out : _GEN_1963; // @[stackmanage_35.scala 4493:55 stackmanage_35.scala 4495:28]
  wire [31:0] _GEN_1968 = pop_32 & Stack_32_io_enable ? $signed(Stack_32_io_dataOut) : $signed(_GEN_1964); // @[stackmanage_35.scala 4493:55 stackmanage_35.scala 4496:25]
  wire  _GEN_1969 = pop_32 & Stack_32_io_enable | _GEN_1965; // @[stackmanage_35.scala 4493:55 stackmanage_35.scala 4497:31]
  wire [31:0] _GEN_1970 = pop_31 & Stack_31_io_enable ? Stack_31_io_hit_out : _GEN_1966; // @[stackmanage_35.scala 4488:55 stackmanage_35.scala 4489:27]
  wire [31:0] _GEN_1971 = pop_31 & Stack_31_io_enable ? Stack_31_io_ray_out : _GEN_1967; // @[stackmanage_35.scala 4488:55 stackmanage_35.scala 4490:28]
  wire [31:0] _GEN_1972 = pop_31 & Stack_31_io_enable ? $signed(Stack_31_io_dataOut) : $signed(_GEN_1968); // @[stackmanage_35.scala 4488:55 stackmanage_35.scala 4491:25]
  wire  _GEN_1973 = pop_31 & Stack_31_io_enable | _GEN_1969; // @[stackmanage_35.scala 4488:55 stackmanage_35.scala 4492:31]
  wire [31:0] _GEN_1974 = pop_30 & Stack_30_io_enable ? Stack_30_io_hit_out : _GEN_1970; // @[stackmanage_35.scala 4483:55 stackmanage_35.scala 4484:27]
  wire [31:0] _GEN_1975 = pop_30 & Stack_30_io_enable ? Stack_30_io_ray_out : _GEN_1971; // @[stackmanage_35.scala 4483:55 stackmanage_35.scala 4485:28]
  wire [31:0] _GEN_1976 = pop_30 & Stack_30_io_enable ? $signed(Stack_30_io_dataOut) : $signed(_GEN_1972); // @[stackmanage_35.scala 4483:55 stackmanage_35.scala 4486:25]
  wire  _GEN_1977 = pop_30 & Stack_30_io_enable | _GEN_1973; // @[stackmanage_35.scala 4483:55 stackmanage_35.scala 4487:31]
  wire [31:0] _GEN_1978 = pop_29 & Stack_29_io_enable ? Stack_29_io_hit_out : _GEN_1974; // @[stackmanage_35.scala 4478:55 stackmanage_35.scala 4479:27]
  wire [31:0] _GEN_1979 = pop_29 & Stack_29_io_enable ? Stack_29_io_ray_out : _GEN_1975; // @[stackmanage_35.scala 4478:55 stackmanage_35.scala 4480:28]
  wire [31:0] _GEN_1980 = pop_29 & Stack_29_io_enable ? $signed(Stack_29_io_dataOut) : $signed(_GEN_1976); // @[stackmanage_35.scala 4478:55 stackmanage_35.scala 4481:25]
  wire  _GEN_1981 = pop_29 & Stack_29_io_enable | _GEN_1977; // @[stackmanage_35.scala 4478:55 stackmanage_35.scala 4482:31]
  wire [31:0] _GEN_1982 = pop_28 & Stack_28_io_enable ? Stack_28_io_hit_out : _GEN_1978; // @[stackmanage_35.scala 4473:55 stackmanage_35.scala 4474:27]
  wire [31:0] _GEN_1983 = pop_28 & Stack_28_io_enable ? Stack_28_io_ray_out : _GEN_1979; // @[stackmanage_35.scala 4473:55 stackmanage_35.scala 4475:28]
  wire [31:0] _GEN_1984 = pop_28 & Stack_28_io_enable ? $signed(Stack_28_io_dataOut) : $signed(_GEN_1980); // @[stackmanage_35.scala 4473:55 stackmanage_35.scala 4476:25]
  wire  _GEN_1985 = pop_28 & Stack_28_io_enable | _GEN_1981; // @[stackmanage_35.scala 4473:55 stackmanage_35.scala 4477:31]
  wire [31:0] _GEN_1986 = pop_27 & Stack_27_io_enable ? Stack_27_io_hit_out : _GEN_1982; // @[stackmanage_35.scala 4468:55 stackmanage_35.scala 4469:27]
  wire [31:0] _GEN_1987 = pop_27 & Stack_27_io_enable ? Stack_27_io_ray_out : _GEN_1983; // @[stackmanage_35.scala 4468:55 stackmanage_35.scala 4470:28]
  wire [31:0] _GEN_1988 = pop_27 & Stack_27_io_enable ? $signed(Stack_27_io_dataOut) : $signed(_GEN_1984); // @[stackmanage_35.scala 4468:55 stackmanage_35.scala 4471:25]
  wire  _GEN_1989 = pop_27 & Stack_27_io_enable | _GEN_1985; // @[stackmanage_35.scala 4468:55 stackmanage_35.scala 4472:31]
  wire [31:0] _GEN_1990 = pop_26 & Stack_26_io_enable ? Stack_26_io_hit_out : _GEN_1986; // @[stackmanage_35.scala 4463:55 stackmanage_35.scala 4464:27]
  wire [31:0] _GEN_1991 = pop_26 & Stack_26_io_enable ? Stack_26_io_ray_out : _GEN_1987; // @[stackmanage_35.scala 4463:55 stackmanage_35.scala 4465:28]
  wire [31:0] _GEN_1992 = pop_26 & Stack_26_io_enable ? $signed(Stack_26_io_dataOut) : $signed(_GEN_1988); // @[stackmanage_35.scala 4463:55 stackmanage_35.scala 4466:25]
  wire  _GEN_1993 = pop_26 & Stack_26_io_enable | _GEN_1989; // @[stackmanage_35.scala 4463:55 stackmanage_35.scala 4467:31]
  wire [31:0] _GEN_1994 = pop_25 & Stack_25_io_enable ? Stack_25_io_hit_out : _GEN_1990; // @[stackmanage_35.scala 4458:56 stackmanage_35.scala 4459:27]
  wire [31:0] _GEN_1995 = pop_25 & Stack_25_io_enable ? Stack_25_io_ray_out : _GEN_1991; // @[stackmanage_35.scala 4458:56 stackmanage_35.scala 4460:28]
  wire [31:0] _GEN_1996 = pop_25 & Stack_25_io_enable ? $signed(Stack_25_io_dataOut) : $signed(_GEN_1992); // @[stackmanage_35.scala 4458:56 stackmanage_35.scala 4461:25]
  wire  _GEN_1997 = pop_25 & Stack_25_io_enable | _GEN_1993; // @[stackmanage_35.scala 4458:56 stackmanage_35.scala 4462:31]
  wire [31:0] _GEN_1998 = pop_24 & Stack_24_io_enable ? Stack_24_io_hit_out : _GEN_1994; // @[stackmanage_35.scala 4453:55 stackmanage_35.scala 4454:27]
  wire [31:0] _GEN_1999 = pop_24 & Stack_24_io_enable ? Stack_24_io_ray_out : _GEN_1995; // @[stackmanage_35.scala 4453:55 stackmanage_35.scala 4455:28]
  wire [31:0] _GEN_2000 = pop_24 & Stack_24_io_enable ? $signed(Stack_24_io_dataOut) : $signed(_GEN_1996); // @[stackmanage_35.scala 4453:55 stackmanage_35.scala 4456:25]
  wire  _GEN_2001 = pop_24 & Stack_24_io_enable | _GEN_1997; // @[stackmanage_35.scala 4453:55 stackmanage_35.scala 4457:31]
  wire [31:0] _GEN_2002 = pop_23 & Stack_23_io_enable ? Stack_23_io_hit_out : _GEN_1998; // @[stackmanage_35.scala 4448:55 stackmanage_35.scala 4449:27]
  wire [31:0] _GEN_2003 = pop_23 & Stack_23_io_enable ? Stack_23_io_ray_out : _GEN_1999; // @[stackmanage_35.scala 4448:55 stackmanage_35.scala 4450:28]
  wire [31:0] _GEN_2004 = pop_23 & Stack_23_io_enable ? $signed(Stack_23_io_dataOut) : $signed(_GEN_2000); // @[stackmanage_35.scala 4448:55 stackmanage_35.scala 4451:25]
  wire  _GEN_2005 = pop_23 & Stack_23_io_enable | _GEN_2001; // @[stackmanage_35.scala 4448:55 stackmanage_35.scala 4452:31]
  wire [31:0] _GEN_2006 = pop_22 & Stack_22_io_enable ? Stack_22_io_hit_out : _GEN_2002; // @[stackmanage_35.scala 4443:55 stackmanage_35.scala 4444:27]
  wire [31:0] _GEN_2007 = pop_22 & Stack_22_io_enable ? Stack_22_io_ray_out : _GEN_2003; // @[stackmanage_35.scala 4443:55 stackmanage_35.scala 4445:28]
  wire [31:0] _GEN_2008 = pop_22 & Stack_22_io_enable ? $signed(Stack_22_io_dataOut) : $signed(_GEN_2004); // @[stackmanage_35.scala 4443:55 stackmanage_35.scala 4446:25]
  wire  _GEN_2009 = pop_22 & Stack_22_io_enable | _GEN_2005; // @[stackmanage_35.scala 4443:55 stackmanage_35.scala 4447:31]
  wire [31:0] _GEN_2010 = pop_21 & Stack_21_io_enable ? Stack_21_io_hit_out : _GEN_2006; // @[stackmanage_35.scala 4438:55 stackmanage_35.scala 4439:27]
  wire [31:0] _GEN_2011 = pop_21 & Stack_21_io_enable ? Stack_21_io_ray_out : _GEN_2007; // @[stackmanage_35.scala 4438:55 stackmanage_35.scala 4440:28]
  wire [31:0] _GEN_2012 = pop_21 & Stack_21_io_enable ? $signed(Stack_21_io_dataOut) : $signed(_GEN_2008); // @[stackmanage_35.scala 4438:55 stackmanage_35.scala 4441:25]
  wire  _GEN_2013 = pop_21 & Stack_21_io_enable | _GEN_2009; // @[stackmanage_35.scala 4438:55 stackmanage_35.scala 4442:31]
  wire [31:0] _GEN_2014 = pop_20 & Stack_20_io_enable ? Stack_20_io_hit_out : _GEN_2010; // @[stackmanage_35.scala 4433:55 stackmanage_35.scala 4434:27]
  wire [31:0] _GEN_2015 = pop_20 & Stack_20_io_enable ? Stack_20_io_ray_out : _GEN_2011; // @[stackmanage_35.scala 4433:55 stackmanage_35.scala 4435:28]
  wire [31:0] _GEN_2016 = pop_20 & Stack_20_io_enable ? $signed(Stack_20_io_dataOut) : $signed(_GEN_2012); // @[stackmanage_35.scala 4433:55 stackmanage_35.scala 4436:25]
  wire  _GEN_2017 = pop_20 & Stack_20_io_enable | _GEN_2013; // @[stackmanage_35.scala 4433:55 stackmanage_35.scala 4437:31]
  wire [31:0] _GEN_2018 = pop_19 & Stack_19_io_enable ? Stack_19_io_hit_out : _GEN_2014; // @[stackmanage_35.scala 4428:55 stackmanage_35.scala 4429:27]
  wire [31:0] _GEN_2019 = pop_19 & Stack_19_io_enable ? Stack_19_io_ray_out : _GEN_2015; // @[stackmanage_35.scala 4428:55 stackmanage_35.scala 4430:28]
  wire [31:0] _GEN_2020 = pop_19 & Stack_19_io_enable ? $signed(Stack_19_io_dataOut) : $signed(_GEN_2016); // @[stackmanage_35.scala 4428:55 stackmanage_35.scala 4431:25]
  wire  _GEN_2021 = pop_19 & Stack_19_io_enable | _GEN_2017; // @[stackmanage_35.scala 4428:55 stackmanage_35.scala 4432:31]
  wire [31:0] _GEN_2022 = pop_18 & Stack_18_io_enable ? Stack_18_io_hit_out : _GEN_2018; // @[stackmanage_35.scala 4423:55 stackmanage_35.scala 4424:27]
  wire [31:0] _GEN_2023 = pop_18 & Stack_18_io_enable ? Stack_18_io_ray_out : _GEN_2019; // @[stackmanage_35.scala 4423:55 stackmanage_35.scala 4425:28]
  wire [31:0] _GEN_2024 = pop_18 & Stack_18_io_enable ? $signed(Stack_18_io_dataOut) : $signed(_GEN_2020); // @[stackmanage_35.scala 4423:55 stackmanage_35.scala 4426:25]
  wire  _GEN_2025 = pop_18 & Stack_18_io_enable | _GEN_2021; // @[stackmanage_35.scala 4423:55 stackmanage_35.scala 4427:31]
  wire [31:0] _GEN_2026 = pop_17 & Stack_17_io_enable ? Stack_17_io_hit_out : _GEN_2022; // @[stackmanage_35.scala 4418:55 stackmanage_35.scala 4419:27]
  wire [31:0] _GEN_2027 = pop_17 & Stack_17_io_enable ? Stack_17_io_ray_out : _GEN_2023; // @[stackmanage_35.scala 4418:55 stackmanage_35.scala 4420:28]
  wire [31:0] _GEN_2028 = pop_17 & Stack_17_io_enable ? $signed(Stack_17_io_dataOut) : $signed(_GEN_2024); // @[stackmanage_35.scala 4418:55 stackmanage_35.scala 4421:25]
  wire  _GEN_2029 = pop_17 & Stack_17_io_enable | _GEN_2025; // @[stackmanage_35.scala 4418:55 stackmanage_35.scala 4422:31]
  wire [31:0] _GEN_2030 = pop_16 & Stack_16_io_enable ? Stack_16_io_hit_out : _GEN_2026; // @[stackmanage_35.scala 4413:55 stackmanage_35.scala 4414:27]
  wire [31:0] _GEN_2031 = pop_16 & Stack_16_io_enable ? Stack_16_io_ray_out : _GEN_2027; // @[stackmanage_35.scala 4413:55 stackmanage_35.scala 4415:28]
  wire [31:0] _GEN_2032 = pop_16 & Stack_16_io_enable ? $signed(Stack_16_io_dataOut) : $signed(_GEN_2028); // @[stackmanage_35.scala 4413:55 stackmanage_35.scala 4416:25]
  wire  _GEN_2033 = pop_16 & Stack_16_io_enable | _GEN_2029; // @[stackmanage_35.scala 4413:55 stackmanage_35.scala 4417:31]
  wire [31:0] _GEN_2034 = pop_15 & Stack_15_io_enable ? Stack_15_io_hit_out : _GEN_2030; // @[stackmanage_35.scala 4408:55 stackmanage_35.scala 4409:27]
  wire [31:0] _GEN_2035 = pop_15 & Stack_15_io_enable ? Stack_15_io_ray_out : _GEN_2031; // @[stackmanage_35.scala 4408:55 stackmanage_35.scala 4410:28]
  wire [31:0] _GEN_2036 = pop_15 & Stack_15_io_enable ? $signed(Stack_15_io_dataOut) : $signed(_GEN_2032); // @[stackmanage_35.scala 4408:55 stackmanage_35.scala 4411:25]
  wire  _GEN_2037 = pop_15 & Stack_15_io_enable | _GEN_2033; // @[stackmanage_35.scala 4408:55 stackmanage_35.scala 4412:31]
  wire [31:0] _GEN_2038 = pop_14 & Stack_14_io_enable ? Stack_14_io_hit_out : _GEN_2034; // @[stackmanage_35.scala 4403:55 stackmanage_35.scala 4404:27]
  wire [31:0] _GEN_2039 = pop_14 & Stack_14_io_enable ? Stack_14_io_ray_out : _GEN_2035; // @[stackmanage_35.scala 4403:55 stackmanage_35.scala 4405:28]
  wire [31:0] _GEN_2040 = pop_14 & Stack_14_io_enable ? $signed(Stack_14_io_dataOut) : $signed(_GEN_2036); // @[stackmanage_35.scala 4403:55 stackmanage_35.scala 4406:25]
  wire  _GEN_2041 = pop_14 & Stack_14_io_enable | _GEN_2037; // @[stackmanage_35.scala 4403:55 stackmanage_35.scala 4407:31]
  wire [31:0] _GEN_2042 = pop_13 & Stack_13_io_enable ? Stack_13_io_hit_out : _GEN_2038; // @[stackmanage_35.scala 4398:55 stackmanage_35.scala 4399:27]
  wire [31:0] _GEN_2043 = pop_13 & Stack_13_io_enable ? Stack_13_io_ray_out : _GEN_2039; // @[stackmanage_35.scala 4398:55 stackmanage_35.scala 4400:28]
  wire [31:0] _GEN_2044 = pop_13 & Stack_13_io_enable ? $signed(Stack_13_io_dataOut) : $signed(_GEN_2040); // @[stackmanage_35.scala 4398:55 stackmanage_35.scala 4401:25]
  wire  _GEN_2045 = pop_13 & Stack_13_io_enable | _GEN_2041; // @[stackmanage_35.scala 4398:55 stackmanage_35.scala 4402:31]
  wire [31:0] _GEN_2046 = pop_12 & Stack_12_io_enable ? Stack_12_io_hit_out : _GEN_2042; // @[stackmanage_35.scala 4393:55 stackmanage_35.scala 4394:27]
  wire [31:0] _GEN_2047 = pop_12 & Stack_12_io_enable ? Stack_12_io_ray_out : _GEN_2043; // @[stackmanage_35.scala 4393:55 stackmanage_35.scala 4395:28]
  wire [31:0] _GEN_2048 = pop_12 & Stack_12_io_enable ? $signed(Stack_12_io_dataOut) : $signed(_GEN_2044); // @[stackmanage_35.scala 4393:55 stackmanage_35.scala 4396:25]
  wire  _GEN_2049 = pop_12 & Stack_12_io_enable | _GEN_2045; // @[stackmanage_35.scala 4393:55 stackmanage_35.scala 4397:31]
  wire [31:0] _GEN_2050 = pop_11 & Stack_11_io_enable ? Stack_11_io_hit_out : _GEN_2046; // @[stackmanage_35.scala 4388:55 stackmanage_35.scala 4389:27]
  wire [31:0] _GEN_2051 = pop_11 & Stack_11_io_enable ? Stack_11_io_ray_out : _GEN_2047; // @[stackmanage_35.scala 4388:55 stackmanage_35.scala 4390:28]
  wire [31:0] _GEN_2052 = pop_11 & Stack_11_io_enable ? $signed(Stack_11_io_dataOut) : $signed(_GEN_2048); // @[stackmanage_35.scala 4388:55 stackmanage_35.scala 4391:25]
  wire  _GEN_2053 = pop_11 & Stack_11_io_enable | _GEN_2049; // @[stackmanage_35.scala 4388:55 stackmanage_35.scala 4392:31]
  wire [31:0] _GEN_2054 = pop_10 & Stack_10_io_enable ? Stack_10_io_hit_out : _GEN_2050; // @[stackmanage_35.scala 4383:55 stackmanage_35.scala 4384:27]
  wire [31:0] _GEN_2055 = pop_10 & Stack_10_io_enable ? Stack_10_io_ray_out : _GEN_2051; // @[stackmanage_35.scala 4383:55 stackmanage_35.scala 4385:28]
  wire [31:0] _GEN_2056 = pop_10 & Stack_10_io_enable ? $signed(Stack_10_io_dataOut) : $signed(_GEN_2052); // @[stackmanage_35.scala 4383:55 stackmanage_35.scala 4386:25]
  wire  _GEN_2057 = pop_10 & Stack_10_io_enable | _GEN_2053; // @[stackmanage_35.scala 4383:55 stackmanage_35.scala 4387:31]
  wire [31:0] _GEN_2058 = pop_9 & Stack_9_io_enable ? Stack_9_io_hit_out : _GEN_2054; // @[stackmanage_35.scala 4378:53 stackmanage_35.scala 4379:27]
  wire [31:0] _GEN_2059 = pop_9 & Stack_9_io_enable ? Stack_9_io_ray_out : _GEN_2055; // @[stackmanage_35.scala 4378:53 stackmanage_35.scala 4380:28]
  wire [31:0] _GEN_2060 = pop_9 & Stack_9_io_enable ? $signed(Stack_9_io_dataOut) : $signed(_GEN_2056); // @[stackmanage_35.scala 4378:53 stackmanage_35.scala 4381:25]
  wire  _GEN_2061 = pop_9 & Stack_9_io_enable | _GEN_2057; // @[stackmanage_35.scala 4378:53 stackmanage_35.scala 4382:31]
  wire [31:0] _GEN_2062 = pop_8 & Stack_8_io_enable ? Stack_8_io_hit_out : _GEN_2058; // @[stackmanage_35.scala 4373:53 stackmanage_35.scala 4374:27]
  wire [31:0] _GEN_2063 = pop_8 & Stack_8_io_enable ? Stack_8_io_ray_out : _GEN_2059; // @[stackmanage_35.scala 4373:53 stackmanage_35.scala 4375:28]
  wire [31:0] _GEN_2064 = pop_8 & Stack_8_io_enable ? $signed(Stack_8_io_dataOut) : $signed(_GEN_2060); // @[stackmanage_35.scala 4373:53 stackmanage_35.scala 4376:25]
  wire  _GEN_2065 = pop_8 & Stack_8_io_enable | _GEN_2061; // @[stackmanage_35.scala 4373:53 stackmanage_35.scala 4377:31]
  wire [31:0] _GEN_2066 = pop_7 & Stack_7_io_enable ? Stack_7_io_hit_out : _GEN_2062; // @[stackmanage_35.scala 4368:53 stackmanage_35.scala 4369:27]
  wire [31:0] _GEN_2067 = pop_7 & Stack_7_io_enable ? Stack_7_io_ray_out : _GEN_2063; // @[stackmanage_35.scala 4368:53 stackmanage_35.scala 4370:28]
  wire [31:0] _GEN_2068 = pop_7 & Stack_7_io_enable ? $signed(Stack_7_io_dataOut) : $signed(_GEN_2064); // @[stackmanage_35.scala 4368:53 stackmanage_35.scala 4371:25]
  wire  _GEN_2069 = pop_7 & Stack_7_io_enable | _GEN_2065; // @[stackmanage_35.scala 4368:53 stackmanage_35.scala 4372:31]
  wire [31:0] _GEN_2070 = pop_6 & Stack_6_io_enable ? Stack_6_io_hit_out : _GEN_2066; // @[stackmanage_35.scala 4363:53 stackmanage_35.scala 4364:27]
  wire [31:0] _GEN_2071 = pop_6 & Stack_6_io_enable ? Stack_6_io_ray_out : _GEN_2067; // @[stackmanage_35.scala 4363:53 stackmanage_35.scala 4365:28]
  wire [31:0] _GEN_2072 = pop_6 & Stack_6_io_enable ? $signed(Stack_6_io_dataOut) : $signed(_GEN_2068); // @[stackmanage_35.scala 4363:53 stackmanage_35.scala 4366:25]
  wire  _GEN_2073 = pop_6 & Stack_6_io_enable | _GEN_2069; // @[stackmanage_35.scala 4363:53 stackmanage_35.scala 4367:31]
  wire [31:0] _GEN_2074 = pop_5 & Stack_5_io_enable ? Stack_5_io_hit_out : _GEN_2070; // @[stackmanage_35.scala 4358:53 stackmanage_35.scala 4359:27]
  wire [31:0] _GEN_2075 = pop_5 & Stack_5_io_enable ? Stack_5_io_ray_out : _GEN_2071; // @[stackmanage_35.scala 4358:53 stackmanage_35.scala 4360:28]
  wire [31:0] _GEN_2076 = pop_5 & Stack_5_io_enable ? $signed(Stack_5_io_dataOut) : $signed(_GEN_2072); // @[stackmanage_35.scala 4358:53 stackmanage_35.scala 4361:25]
  wire  _GEN_2077 = pop_5 & Stack_5_io_enable | _GEN_2073; // @[stackmanage_35.scala 4358:53 stackmanage_35.scala 4362:31]
  wire [31:0] _GEN_2078 = pop_4 & Stack_4_io_enable ? Stack_4_io_hit_out : _GEN_2074; // @[stackmanage_35.scala 4353:53 stackmanage_35.scala 4354:27]
  wire [31:0] _GEN_2079 = pop_4 & Stack_4_io_enable ? Stack_4_io_ray_out : _GEN_2075; // @[stackmanage_35.scala 4353:53 stackmanage_35.scala 4355:28]
  wire [31:0] _GEN_2080 = pop_4 & Stack_4_io_enable ? $signed(Stack_4_io_dataOut) : $signed(_GEN_2076); // @[stackmanage_35.scala 4353:53 stackmanage_35.scala 4356:25]
  wire  _GEN_2081 = pop_4 & Stack_4_io_enable | _GEN_2077; // @[stackmanage_35.scala 4353:53 stackmanage_35.scala 4357:31]
  wire [31:0] _GEN_2082 = pop_3 & Stack_3_io_enable ? Stack_3_io_hit_out : _GEN_2078; // @[stackmanage_35.scala 4348:53 stackmanage_35.scala 4349:27]
  wire [31:0] _GEN_2083 = pop_3 & Stack_3_io_enable ? Stack_3_io_ray_out : _GEN_2079; // @[stackmanage_35.scala 4348:53 stackmanage_35.scala 4350:28]
  wire [31:0] _GEN_2084 = pop_3 & Stack_3_io_enable ? $signed(Stack_3_io_dataOut) : $signed(_GEN_2080); // @[stackmanage_35.scala 4348:53 stackmanage_35.scala 4351:25]
  wire  _GEN_2085 = pop_3 & Stack_3_io_enable | _GEN_2081; // @[stackmanage_35.scala 4348:53 stackmanage_35.scala 4352:31]
  wire  _GEN_2089 = pop_2 & Stack_2_io_enable | _GEN_2085; // @[stackmanage_35.scala 4343:53 stackmanage_35.scala 4347:31]
  wire  _GEN_2093 = pop_1 & Stack_1_io_enable | _GEN_2089; // @[stackmanage_35.scala 4338:53 stackmanage_35.scala 4342:31]
  wire  _GEN_2097 = pop_0 & Stack_0_io_enable | _GEN_2093; // @[stackmanage_35.scala 4332:48 stackmanage_35.scala 4337:31]
  reg  dispatch_0; // @[stackmanage_35.scala 4520:41]
  reg  dispatch_1; // @[stackmanage_35.scala 4521:41]
  reg  dispatch_2; // @[stackmanage_35.scala 4522:41]
  reg  dispatch_3; // @[stackmanage_35.scala 4523:41]
  reg  dispatch_4; // @[stackmanage_35.scala 4524:41]
  reg  dispatch_5; // @[stackmanage_35.scala 4525:41]
  reg  dispatch_6; // @[stackmanage_35.scala 4526:41]
  reg  dispatch_7; // @[stackmanage_35.scala 4527:41]
  reg  dispatch_8; // @[stackmanage_35.scala 4528:41]
  reg  dispatch_9; // @[stackmanage_35.scala 4529:41]
  reg  dispatch_10; // @[stackmanage_35.scala 4531:42]
  reg  dispatch_11; // @[stackmanage_35.scala 4532:42]
  reg  dispatch_12; // @[stackmanage_35.scala 4533:42]
  reg  dispatch_13; // @[stackmanage_35.scala 4534:42]
  reg  dispatch_14; // @[stackmanage_35.scala 4535:42]
  reg  dispatch_15; // @[stackmanage_35.scala 4536:42]
  reg  dispatch_16; // @[stackmanage_35.scala 4537:42]
  reg  dispatch_17; // @[stackmanage_35.scala 4538:42]
  reg  dispatch_18; // @[stackmanage_35.scala 4539:42]
  reg  dispatch_19; // @[stackmanage_35.scala 4540:42]
  reg  dispatch_20; // @[stackmanage_35.scala 4542:42]
  reg  dispatch_21; // @[stackmanage_35.scala 4543:42]
  reg  dispatch_22; // @[stackmanage_35.scala 4544:42]
  reg  dispatch_23; // @[stackmanage_35.scala 4545:42]
  reg  dispatch_24; // @[stackmanage_35.scala 4546:42]
  reg  dispatch_25; // @[stackmanage_35.scala 4547:42]
  reg  dispatch_26; // @[stackmanage_35.scala 4548:42]
  reg  dispatch_27; // @[stackmanage_35.scala 4549:42]
  reg  dispatch_28; // @[stackmanage_35.scala 4550:42]
  reg  dispatch_29; // @[stackmanage_35.scala 4551:42]
  reg  dispatch_30; // @[stackmanage_35.scala 4553:42]
  reg  dispatch_31; // @[stackmanage_35.scala 4554:42]
  reg  dispatch_32; // @[stackmanage_35.scala 4555:42]
  reg  dispatch_33; // @[stackmanage_35.scala 4556:42]
  reg  dispatch_34; // @[stackmanage_35.scala 4557:42]
  reg  dispatch_no_match; // @[stackmanage_35.scala 4558:42]
  reg  empty_0; // @[stackmanage_35.scala 4562:42]
  reg  empty_1; // @[stackmanage_35.scala 4563:42]
  reg  empty_2; // @[stackmanage_35.scala 4564:42]
  reg  empty_3; // @[stackmanage_35.scala 4565:42]
  reg  empty_4; // @[stackmanage_35.scala 4566:42]
  reg  empty_5; // @[stackmanage_35.scala 4567:42]
  reg  empty_6; // @[stackmanage_35.scala 4568:42]
  reg  empty_7; // @[stackmanage_35.scala 4569:42]
  reg  empty_8; // @[stackmanage_35.scala 4570:42]
  reg  empty_9; // @[stackmanage_35.scala 4571:42]
  reg  empty_10; // @[stackmanage_35.scala 4573:43]
  reg  empty_11; // @[stackmanage_35.scala 4574:43]
  reg  empty_12; // @[stackmanage_35.scala 4575:43]
  reg  empty_13; // @[stackmanage_35.scala 4576:43]
  reg  empty_14; // @[stackmanage_35.scala 4577:43]
  reg  empty_15; // @[stackmanage_35.scala 4578:43]
  reg  empty_16; // @[stackmanage_35.scala 4579:43]
  reg  empty_17; // @[stackmanage_35.scala 4580:43]
  reg  empty_18; // @[stackmanage_35.scala 4581:43]
  reg  empty_19; // @[stackmanage_35.scala 4582:43]
  reg  empty_20; // @[stackmanage_35.scala 4584:43]
  reg  empty_21; // @[stackmanage_35.scala 4585:43]
  reg  empty_22; // @[stackmanage_35.scala 4586:43]
  reg  empty_23; // @[stackmanage_35.scala 4587:43]
  reg  empty_24; // @[stackmanage_35.scala 4588:43]
  reg  empty_25; // @[stackmanage_35.scala 4589:43]
  reg  empty_26; // @[stackmanage_35.scala 4590:43]
  reg  empty_27; // @[stackmanage_35.scala 4591:43]
  reg  empty_28; // @[stackmanage_35.scala 4592:43]
  reg  empty_29; // @[stackmanage_35.scala 4593:43]
  reg  empty_30; // @[stackmanage_35.scala 4595:43]
  reg  empty_31; // @[stackmanage_35.scala 4596:43]
  reg  empty_32; // @[stackmanage_35.scala 4597:43]
  reg  empty_33; // @[stackmanage_35.scala 4598:43]
  reg  empty_34; // @[stackmanage_35.scala 4599:43]
  wire  _T_317 = pop_0 & empty_0; // @[stackmanage_35.scala 4643:22]
  wire  _T_320 = pop_1 & empty_1; // @[stackmanage_35.scala 4679:27]
  wire  _T_323 = pop_2 & empty_2; // @[stackmanage_35.scala 4716:27]
  wire  _T_326 = pop_3 & empty_3; // @[stackmanage_35.scala 4754:27]
  wire  _T_329 = pop_4 & empty_4; // @[stackmanage_35.scala 4792:27]
  wire  _T_332 = pop_5 & empty_5; // @[stackmanage_35.scala 4830:27]
  wire  _T_335 = pop_6 & empty_6; // @[stackmanage_35.scala 4868:27]
  wire  _T_338 = pop_7 & empty_7; // @[stackmanage_35.scala 4906:27]
  wire  _T_341 = pop_8 & empty_8; // @[stackmanage_35.scala 4944:27]
  wire  _T_344 = pop_9 & empty_9; // @[stackmanage_35.scala 4981:27]
  wire  _T_347 = pop_10 & empty_10; // @[stackmanage_35.scala 5019:28]
  wire  _T_350 = pop_11 & empty_11; // @[stackmanage_35.scala 5056:28]
  wire  _T_353 = pop_12 & empty_12; // @[stackmanage_35.scala 5093:28]
  wire  _T_356 = pop_13 & empty_13; // @[stackmanage_35.scala 5130:28]
  wire  _T_359 = pop_14 & empty_14; // @[stackmanage_35.scala 5167:28]
  wire  _T_362 = pop_15 & empty_15; // @[stackmanage_35.scala 5204:28]
  wire  _T_365 = pop_16 & empty_16; // @[stackmanage_35.scala 5241:28]
  wire  _T_368 = pop_17 & empty_17; // @[stackmanage_35.scala 5278:28]
  wire  _T_371 = pop_18 & empty_18; // @[stackmanage_35.scala 5315:28]
  wire  _T_374 = pop_19 & empty_19; // @[stackmanage_35.scala 5352:28]
  wire  _T_377 = pop_20 & empty_20; // @[stackmanage_35.scala 5389:28]
  wire  _T_380 = pop_21 & empty_21; // @[stackmanage_35.scala 5426:28]
  wire  _T_383 = pop_22 & empty_22; // @[stackmanage_35.scala 5463:28]
  wire  _T_386 = pop_23 & empty_23; // @[stackmanage_35.scala 5500:28]
  wire  _T_389 = pop_24 & empty_24; // @[stackmanage_35.scala 5537:28]
  wire  _T_392 = pop_25 & empty_25; // @[stackmanage_35.scala 5574:28]
  wire  _T_395 = pop_26 & empty_26; // @[stackmanage_35.scala 5611:30]
  wire  _T_398 = pop_27 & empty_27; // @[stackmanage_35.scala 5648:28]
  wire  _T_401 = pop_28 & empty_28; // @[stackmanage_35.scala 5685:28]
  wire  _T_404 = pop_29 & empty_29; // @[stackmanage_35.scala 5722:28]
  wire  _T_407 = pop_30 & empty_30; // @[stackmanage_35.scala 5759:29]
  wire  _T_410 = pop_31 & empty_31; // @[stackmanage_35.scala 5796:29]
  wire  _T_413 = pop_32 & empty_32; // @[stackmanage_35.scala 5833:29]
  wire  _T_416 = pop_33 & empty_33; // @[stackmanage_35.scala 5871:29]
  wire  _T_419 = pop_34 & empty_34; // @[stackmanage_35.scala 5908:29]
  wire  _GEN_2102 = pop_33 & empty_33 ? 1'h0 : _T_419; // @[stackmanage_35.scala 5871:46 stackmanage_35.scala 5907:34]
  wire  _GEN_2105 = pop_32 & empty_32 ? 1'h0 : _T_416; // @[stackmanage_35.scala 5833:46 stackmanage_35.scala 5868:34]
  wire  _GEN_2106 = pop_32 & empty_32 ? 1'h0 : _GEN_2102; // @[stackmanage_35.scala 5833:46 stackmanage_35.scala 5869:34]
  wire  _GEN_2109 = pop_31 & empty_31 ? 1'h0 : _T_413; // @[stackmanage_35.scala 5796:46 stackmanage_35.scala 5830:34]
  wire  _GEN_2110 = pop_31 & empty_31 ? 1'h0 : _GEN_2105; // @[stackmanage_35.scala 5796:46 stackmanage_35.scala 5831:34]
  wire  _GEN_2111 = pop_31 & empty_31 ? 1'h0 : _GEN_2106; // @[stackmanage_35.scala 5796:46 stackmanage_35.scala 5832:34]
  wire  _GEN_2114 = pop_30 & empty_30 ? 1'h0 : _T_410; // @[stackmanage_35.scala 5759:46 stackmanage_35.scala 5792:34]
  wire  _GEN_2115 = pop_30 & empty_30 ? 1'h0 : _GEN_2109; // @[stackmanage_35.scala 5759:46 stackmanage_35.scala 5793:34]
  wire  _GEN_2116 = pop_30 & empty_30 ? 1'h0 : _GEN_2110; // @[stackmanage_35.scala 5759:46 stackmanage_35.scala 5794:34]
  wire  _GEN_2117 = pop_30 & empty_30 ? 1'h0 : _GEN_2111; // @[stackmanage_35.scala 5759:46 stackmanage_35.scala 5795:34]
  wire  _GEN_2120 = pop_29 & empty_29 ? 1'h0 : _T_407; // @[stackmanage_35.scala 5722:45 stackmanage_35.scala 5754:34]
  wire  _GEN_2121 = pop_29 & empty_29 ? 1'h0 : _GEN_2114; // @[stackmanage_35.scala 5722:45 stackmanage_35.scala 5755:34]
  wire  _GEN_2122 = pop_29 & empty_29 ? 1'h0 : _GEN_2115; // @[stackmanage_35.scala 5722:45 stackmanage_35.scala 5756:34]
  wire  _GEN_2123 = pop_29 & empty_29 ? 1'h0 : _GEN_2116; // @[stackmanage_35.scala 5722:45 stackmanage_35.scala 5757:34]
  wire  _GEN_2124 = pop_29 & empty_29 ? 1'h0 : _GEN_2117; // @[stackmanage_35.scala 5722:45 stackmanage_35.scala 5758:34]
  wire  _GEN_2127 = pop_28 & empty_28 ? 1'h0 : _T_404; // @[stackmanage_35.scala 5685:45 stackmanage_35.scala 5716:34]
  wire  _GEN_2128 = pop_28 & empty_28 ? 1'h0 : _GEN_2120; // @[stackmanage_35.scala 5685:45 stackmanage_35.scala 5717:34]
  wire  _GEN_2129 = pop_28 & empty_28 ? 1'h0 : _GEN_2121; // @[stackmanage_35.scala 5685:45 stackmanage_35.scala 5718:34]
  wire  _GEN_2130 = pop_28 & empty_28 ? 1'h0 : _GEN_2122; // @[stackmanage_35.scala 5685:45 stackmanage_35.scala 5719:34]
  wire  _GEN_2131 = pop_28 & empty_28 ? 1'h0 : _GEN_2123; // @[stackmanage_35.scala 5685:45 stackmanage_35.scala 5720:34]
  wire  _GEN_2132 = pop_28 & empty_28 ? 1'h0 : _GEN_2124; // @[stackmanage_35.scala 5685:45 stackmanage_35.scala 5721:34]
  wire  _GEN_2135 = pop_27 & empty_27 ? 1'h0 : _T_401; // @[stackmanage_35.scala 5648:45 stackmanage_35.scala 5678:34]
  wire  _GEN_2136 = pop_27 & empty_27 ? 1'h0 : _GEN_2127; // @[stackmanage_35.scala 5648:45 stackmanage_35.scala 5679:34]
  wire  _GEN_2137 = pop_27 & empty_27 ? 1'h0 : _GEN_2128; // @[stackmanage_35.scala 5648:45 stackmanage_35.scala 5680:34]
  wire  _GEN_2138 = pop_27 & empty_27 ? 1'h0 : _GEN_2129; // @[stackmanage_35.scala 5648:45 stackmanage_35.scala 5681:34]
  wire  _GEN_2139 = pop_27 & empty_27 ? 1'h0 : _GEN_2130; // @[stackmanage_35.scala 5648:45 stackmanage_35.scala 5682:34]
  wire  _GEN_2140 = pop_27 & empty_27 ? 1'h0 : _GEN_2131; // @[stackmanage_35.scala 5648:45 stackmanage_35.scala 5683:34]
  wire  _GEN_2141 = pop_27 & empty_27 ? 1'h0 : _GEN_2132; // @[stackmanage_35.scala 5648:45 stackmanage_35.scala 5684:34]
  wire  _GEN_2144 = pop_26 & empty_26 ? 1'h0 : _T_398; // @[stackmanage_35.scala 5611:47 stackmanage_35.scala 5640:34]
  wire  _GEN_2145 = pop_26 & empty_26 ? 1'h0 : _GEN_2135; // @[stackmanage_35.scala 5611:47 stackmanage_35.scala 5641:34]
  wire  _GEN_2146 = pop_26 & empty_26 ? 1'h0 : _GEN_2136; // @[stackmanage_35.scala 5611:47 stackmanage_35.scala 5642:34]
  wire  _GEN_2147 = pop_26 & empty_26 ? 1'h0 : _GEN_2137; // @[stackmanage_35.scala 5611:47 stackmanage_35.scala 5643:34]
  wire  _GEN_2148 = pop_26 & empty_26 ? 1'h0 : _GEN_2138; // @[stackmanage_35.scala 5611:47 stackmanage_35.scala 5644:34]
  wire  _GEN_2149 = pop_26 & empty_26 ? 1'h0 : _GEN_2139; // @[stackmanage_35.scala 5611:47 stackmanage_35.scala 5645:34]
  wire  _GEN_2150 = pop_26 & empty_26 ? 1'h0 : _GEN_2140; // @[stackmanage_35.scala 5611:47 stackmanage_35.scala 5646:34]
  wire  _GEN_2151 = pop_26 & empty_26 ? 1'h0 : _GEN_2141; // @[stackmanage_35.scala 5611:47 stackmanage_35.scala 5647:34]
  wire  _GEN_2154 = pop_25 & empty_25 ? 1'h0 : _T_395; // @[stackmanage_35.scala 5574:45 stackmanage_35.scala 5602:34]
  wire  _GEN_2155 = pop_25 & empty_25 ? 1'h0 : _GEN_2144; // @[stackmanage_35.scala 5574:45 stackmanage_35.scala 5603:34]
  wire  _GEN_2156 = pop_25 & empty_25 ? 1'h0 : _GEN_2145; // @[stackmanage_35.scala 5574:45 stackmanage_35.scala 5604:34]
  wire  _GEN_2157 = pop_25 & empty_25 ? 1'h0 : _GEN_2146; // @[stackmanage_35.scala 5574:45 stackmanage_35.scala 5605:34]
  wire  _GEN_2158 = pop_25 & empty_25 ? 1'h0 : _GEN_2147; // @[stackmanage_35.scala 5574:45 stackmanage_35.scala 5606:34]
  wire  _GEN_2159 = pop_25 & empty_25 ? 1'h0 : _GEN_2148; // @[stackmanage_35.scala 5574:45 stackmanage_35.scala 5607:34]
  wire  _GEN_2160 = pop_25 & empty_25 ? 1'h0 : _GEN_2149; // @[stackmanage_35.scala 5574:45 stackmanage_35.scala 5608:34]
  wire  _GEN_2161 = pop_25 & empty_25 ? 1'h0 : _GEN_2150; // @[stackmanage_35.scala 5574:45 stackmanage_35.scala 5609:34]
  wire  _GEN_2162 = pop_25 & empty_25 ? 1'h0 : _GEN_2151; // @[stackmanage_35.scala 5574:45 stackmanage_35.scala 5610:34]
  wire  _GEN_2165 = pop_24 & empty_24 ? 1'h0 : _T_392; // @[stackmanage_35.scala 5537:45 stackmanage_35.scala 5564:34]
  wire  _GEN_2166 = pop_24 & empty_24 ? 1'h0 : _GEN_2154; // @[stackmanage_35.scala 5537:45 stackmanage_35.scala 5565:34]
  wire  _GEN_2167 = pop_24 & empty_24 ? 1'h0 : _GEN_2155; // @[stackmanage_35.scala 5537:45 stackmanage_35.scala 5566:34]
  wire  _GEN_2168 = pop_24 & empty_24 ? 1'h0 : _GEN_2156; // @[stackmanage_35.scala 5537:45 stackmanage_35.scala 5567:34]
  wire  _GEN_2169 = pop_24 & empty_24 ? 1'h0 : _GEN_2157; // @[stackmanage_35.scala 5537:45 stackmanage_35.scala 5568:34]
  wire  _GEN_2170 = pop_24 & empty_24 ? 1'h0 : _GEN_2158; // @[stackmanage_35.scala 5537:45 stackmanage_35.scala 5569:34]
  wire  _GEN_2171 = pop_24 & empty_24 ? 1'h0 : _GEN_2159; // @[stackmanage_35.scala 5537:45 stackmanage_35.scala 5570:34]
  wire  _GEN_2172 = pop_24 & empty_24 ? 1'h0 : _GEN_2160; // @[stackmanage_35.scala 5537:45 stackmanage_35.scala 5571:34]
  wire  _GEN_2173 = pop_24 & empty_24 ? 1'h0 : _GEN_2161; // @[stackmanage_35.scala 5537:45 stackmanage_35.scala 5572:34]
  wire  _GEN_2174 = pop_24 & empty_24 ? 1'h0 : _GEN_2162; // @[stackmanage_35.scala 5537:45 stackmanage_35.scala 5573:34]
  wire  _GEN_2177 = pop_23 & empty_23 ? 1'h0 : _T_389; // @[stackmanage_35.scala 5500:45 stackmanage_35.scala 5526:34]
  wire  _GEN_2178 = pop_23 & empty_23 ? 1'h0 : _GEN_2165; // @[stackmanage_35.scala 5500:45 stackmanage_35.scala 5527:34]
  wire  _GEN_2179 = pop_23 & empty_23 ? 1'h0 : _GEN_2166; // @[stackmanage_35.scala 5500:45 stackmanage_35.scala 5528:34]
  wire  _GEN_2180 = pop_23 & empty_23 ? 1'h0 : _GEN_2167; // @[stackmanage_35.scala 5500:45 stackmanage_35.scala 5529:34]
  wire  _GEN_2181 = pop_23 & empty_23 ? 1'h0 : _GEN_2168; // @[stackmanage_35.scala 5500:45 stackmanage_35.scala 5530:34]
  wire  _GEN_2182 = pop_23 & empty_23 ? 1'h0 : _GEN_2169; // @[stackmanage_35.scala 5500:45 stackmanage_35.scala 5531:34]
  wire  _GEN_2183 = pop_23 & empty_23 ? 1'h0 : _GEN_2170; // @[stackmanage_35.scala 5500:45 stackmanage_35.scala 5532:34]
  wire  _GEN_2184 = pop_23 & empty_23 ? 1'h0 : _GEN_2171; // @[stackmanage_35.scala 5500:45 stackmanage_35.scala 5533:34]
  wire  _GEN_2185 = pop_23 & empty_23 ? 1'h0 : _GEN_2172; // @[stackmanage_35.scala 5500:45 stackmanage_35.scala 5534:34]
  wire  _GEN_2186 = pop_23 & empty_23 ? 1'h0 : _GEN_2173; // @[stackmanage_35.scala 5500:45 stackmanage_35.scala 5535:34]
  wire  _GEN_2187 = pop_23 & empty_23 ? 1'h0 : _GEN_2174; // @[stackmanage_35.scala 5500:45 stackmanage_35.scala 5536:34]
  wire  _GEN_2190 = pop_22 & empty_22 ? 1'h0 : _T_386; // @[stackmanage_35.scala 5463:45 stackmanage_35.scala 5488:34]
  wire  _GEN_2191 = pop_22 & empty_22 ? 1'h0 : _GEN_2177; // @[stackmanage_35.scala 5463:45 stackmanage_35.scala 5489:34]
  wire  _GEN_2192 = pop_22 & empty_22 ? 1'h0 : _GEN_2178; // @[stackmanage_35.scala 5463:45 stackmanage_35.scala 5490:34]
  wire  _GEN_2193 = pop_22 & empty_22 ? 1'h0 : _GEN_2179; // @[stackmanage_35.scala 5463:45 stackmanage_35.scala 5491:34]
  wire  _GEN_2194 = pop_22 & empty_22 ? 1'h0 : _GEN_2180; // @[stackmanage_35.scala 5463:45 stackmanage_35.scala 5492:34]
  wire  _GEN_2195 = pop_22 & empty_22 ? 1'h0 : _GEN_2181; // @[stackmanage_35.scala 5463:45 stackmanage_35.scala 5493:34]
  wire  _GEN_2196 = pop_22 & empty_22 ? 1'h0 : _GEN_2182; // @[stackmanage_35.scala 5463:45 stackmanage_35.scala 5494:34]
  wire  _GEN_2197 = pop_22 & empty_22 ? 1'h0 : _GEN_2183; // @[stackmanage_35.scala 5463:45 stackmanage_35.scala 5495:34]
  wire  _GEN_2198 = pop_22 & empty_22 ? 1'h0 : _GEN_2184; // @[stackmanage_35.scala 5463:45 stackmanage_35.scala 5496:34]
  wire  _GEN_2199 = pop_22 & empty_22 ? 1'h0 : _GEN_2185; // @[stackmanage_35.scala 5463:45 stackmanage_35.scala 5497:34]
  wire  _GEN_2200 = pop_22 & empty_22 ? 1'h0 : _GEN_2186; // @[stackmanage_35.scala 5463:45 stackmanage_35.scala 5498:34]
  wire  _GEN_2201 = pop_22 & empty_22 ? 1'h0 : _GEN_2187; // @[stackmanage_35.scala 5463:45 stackmanage_35.scala 5499:34]
  wire  _GEN_2204 = pop_21 & empty_21 ? 1'h0 : _T_383; // @[stackmanage_35.scala 5426:45 stackmanage_35.scala 5450:34]
  wire  _GEN_2205 = pop_21 & empty_21 ? 1'h0 : _GEN_2190; // @[stackmanage_35.scala 5426:45 stackmanage_35.scala 5451:34]
  wire  _GEN_2206 = pop_21 & empty_21 ? 1'h0 : _GEN_2191; // @[stackmanage_35.scala 5426:45 stackmanage_35.scala 5452:34]
  wire  _GEN_2207 = pop_21 & empty_21 ? 1'h0 : _GEN_2192; // @[stackmanage_35.scala 5426:45 stackmanage_35.scala 5453:34]
  wire  _GEN_2208 = pop_21 & empty_21 ? 1'h0 : _GEN_2193; // @[stackmanage_35.scala 5426:45 stackmanage_35.scala 5454:34]
  wire  _GEN_2209 = pop_21 & empty_21 ? 1'h0 : _GEN_2194; // @[stackmanage_35.scala 5426:45 stackmanage_35.scala 5455:34]
  wire  _GEN_2210 = pop_21 & empty_21 ? 1'h0 : _GEN_2195; // @[stackmanage_35.scala 5426:45 stackmanage_35.scala 5456:34]
  wire  _GEN_2211 = pop_21 & empty_21 ? 1'h0 : _GEN_2196; // @[stackmanage_35.scala 5426:45 stackmanage_35.scala 5457:34]
  wire  _GEN_2212 = pop_21 & empty_21 ? 1'h0 : _GEN_2197; // @[stackmanage_35.scala 5426:45 stackmanage_35.scala 5458:34]
  wire  _GEN_2213 = pop_21 & empty_21 ? 1'h0 : _GEN_2198; // @[stackmanage_35.scala 5426:45 stackmanage_35.scala 5459:34]
  wire  _GEN_2214 = pop_21 & empty_21 ? 1'h0 : _GEN_2199; // @[stackmanage_35.scala 5426:45 stackmanage_35.scala 5460:34]
  wire  _GEN_2215 = pop_21 & empty_21 ? 1'h0 : _GEN_2200; // @[stackmanage_35.scala 5426:45 stackmanage_35.scala 5461:34]
  wire  _GEN_2216 = pop_21 & empty_21 ? 1'h0 : _GEN_2201; // @[stackmanage_35.scala 5426:45 stackmanage_35.scala 5462:34]
  wire  _GEN_2219 = pop_20 & empty_20 ? 1'h0 : _T_380; // @[stackmanage_35.scala 5389:45 stackmanage_35.scala 5412:34]
  wire  _GEN_2220 = pop_20 & empty_20 ? 1'h0 : _GEN_2204; // @[stackmanage_35.scala 5389:45 stackmanage_35.scala 5413:34]
  wire  _GEN_2221 = pop_20 & empty_20 ? 1'h0 : _GEN_2205; // @[stackmanage_35.scala 5389:45 stackmanage_35.scala 5414:34]
  wire  _GEN_2222 = pop_20 & empty_20 ? 1'h0 : _GEN_2206; // @[stackmanage_35.scala 5389:45 stackmanage_35.scala 5415:34]
  wire  _GEN_2223 = pop_20 & empty_20 ? 1'h0 : _GEN_2207; // @[stackmanage_35.scala 5389:45 stackmanage_35.scala 5416:34]
  wire  _GEN_2224 = pop_20 & empty_20 ? 1'h0 : _GEN_2208; // @[stackmanage_35.scala 5389:45 stackmanage_35.scala 5417:34]
  wire  _GEN_2225 = pop_20 & empty_20 ? 1'h0 : _GEN_2209; // @[stackmanage_35.scala 5389:45 stackmanage_35.scala 5418:34]
  wire  _GEN_2226 = pop_20 & empty_20 ? 1'h0 : _GEN_2210; // @[stackmanage_35.scala 5389:45 stackmanage_35.scala 5419:34]
  wire  _GEN_2227 = pop_20 & empty_20 ? 1'h0 : _GEN_2211; // @[stackmanage_35.scala 5389:45 stackmanage_35.scala 5420:34]
  wire  _GEN_2228 = pop_20 & empty_20 ? 1'h0 : _GEN_2212; // @[stackmanage_35.scala 5389:45 stackmanage_35.scala 5421:34]
  wire  _GEN_2229 = pop_20 & empty_20 ? 1'h0 : _GEN_2213; // @[stackmanage_35.scala 5389:45 stackmanage_35.scala 5422:34]
  wire  _GEN_2230 = pop_20 & empty_20 ? 1'h0 : _GEN_2214; // @[stackmanage_35.scala 5389:45 stackmanage_35.scala 5423:34]
  wire  _GEN_2231 = pop_20 & empty_20 ? 1'h0 : _GEN_2215; // @[stackmanage_35.scala 5389:45 stackmanage_35.scala 5424:34]
  wire  _GEN_2232 = pop_20 & empty_20 ? 1'h0 : _GEN_2216; // @[stackmanage_35.scala 5389:45 stackmanage_35.scala 5425:34]
  wire  _GEN_2235 = pop_19 & empty_19 ? 1'h0 : _T_377; // @[stackmanage_35.scala 5352:45 stackmanage_35.scala 5374:34]
  wire  _GEN_2236 = pop_19 & empty_19 ? 1'h0 : _GEN_2219; // @[stackmanage_35.scala 5352:45 stackmanage_35.scala 5375:34]
  wire  _GEN_2237 = pop_19 & empty_19 ? 1'h0 : _GEN_2220; // @[stackmanage_35.scala 5352:45 stackmanage_35.scala 5376:34]
  wire  _GEN_2238 = pop_19 & empty_19 ? 1'h0 : _GEN_2221; // @[stackmanage_35.scala 5352:45 stackmanage_35.scala 5377:34]
  wire  _GEN_2239 = pop_19 & empty_19 ? 1'h0 : _GEN_2222; // @[stackmanage_35.scala 5352:45 stackmanage_35.scala 5378:34]
  wire  _GEN_2240 = pop_19 & empty_19 ? 1'h0 : _GEN_2223; // @[stackmanage_35.scala 5352:45 stackmanage_35.scala 5379:34]
  wire  _GEN_2241 = pop_19 & empty_19 ? 1'h0 : _GEN_2224; // @[stackmanage_35.scala 5352:45 stackmanage_35.scala 5380:34]
  wire  _GEN_2242 = pop_19 & empty_19 ? 1'h0 : _GEN_2225; // @[stackmanage_35.scala 5352:45 stackmanage_35.scala 5381:34]
  wire  _GEN_2243 = pop_19 & empty_19 ? 1'h0 : _GEN_2226; // @[stackmanage_35.scala 5352:45 stackmanage_35.scala 5382:34]
  wire  _GEN_2244 = pop_19 & empty_19 ? 1'h0 : _GEN_2227; // @[stackmanage_35.scala 5352:45 stackmanage_35.scala 5383:34]
  wire  _GEN_2245 = pop_19 & empty_19 ? 1'h0 : _GEN_2228; // @[stackmanage_35.scala 5352:45 stackmanage_35.scala 5384:34]
  wire  _GEN_2246 = pop_19 & empty_19 ? 1'h0 : _GEN_2229; // @[stackmanage_35.scala 5352:45 stackmanage_35.scala 5385:34]
  wire  _GEN_2247 = pop_19 & empty_19 ? 1'h0 : _GEN_2230; // @[stackmanage_35.scala 5352:45 stackmanage_35.scala 5386:34]
  wire  _GEN_2248 = pop_19 & empty_19 ? 1'h0 : _GEN_2231; // @[stackmanage_35.scala 5352:45 stackmanage_35.scala 5387:34]
  wire  _GEN_2249 = pop_19 & empty_19 ? 1'h0 : _GEN_2232; // @[stackmanage_35.scala 5352:45 stackmanage_35.scala 5388:34]
  wire  _GEN_2252 = pop_18 & empty_18 ? 1'h0 : _T_374; // @[stackmanage_35.scala 5315:45 stackmanage_35.scala 5336:34]
  wire  _GEN_2253 = pop_18 & empty_18 ? 1'h0 : _GEN_2235; // @[stackmanage_35.scala 5315:45 stackmanage_35.scala 5337:34]
  wire  _GEN_2254 = pop_18 & empty_18 ? 1'h0 : _GEN_2236; // @[stackmanage_35.scala 5315:45 stackmanage_35.scala 5338:34]
  wire  _GEN_2255 = pop_18 & empty_18 ? 1'h0 : _GEN_2237; // @[stackmanage_35.scala 5315:45 stackmanage_35.scala 5339:34]
  wire  _GEN_2256 = pop_18 & empty_18 ? 1'h0 : _GEN_2238; // @[stackmanage_35.scala 5315:45 stackmanage_35.scala 5340:34]
  wire  _GEN_2257 = pop_18 & empty_18 ? 1'h0 : _GEN_2239; // @[stackmanage_35.scala 5315:45 stackmanage_35.scala 5341:34]
  wire  _GEN_2258 = pop_18 & empty_18 ? 1'h0 : _GEN_2240; // @[stackmanage_35.scala 5315:45 stackmanage_35.scala 5342:34]
  wire  _GEN_2259 = pop_18 & empty_18 ? 1'h0 : _GEN_2241; // @[stackmanage_35.scala 5315:45 stackmanage_35.scala 5343:34]
  wire  _GEN_2260 = pop_18 & empty_18 ? 1'h0 : _GEN_2242; // @[stackmanage_35.scala 5315:45 stackmanage_35.scala 5344:34]
  wire  _GEN_2261 = pop_18 & empty_18 ? 1'h0 : _GEN_2243; // @[stackmanage_35.scala 5315:45 stackmanage_35.scala 5345:34]
  wire  _GEN_2262 = pop_18 & empty_18 ? 1'h0 : _GEN_2244; // @[stackmanage_35.scala 5315:45 stackmanage_35.scala 5346:34]
  wire  _GEN_2263 = pop_18 & empty_18 ? 1'h0 : _GEN_2245; // @[stackmanage_35.scala 5315:45 stackmanage_35.scala 5347:34]
  wire  _GEN_2264 = pop_18 & empty_18 ? 1'h0 : _GEN_2246; // @[stackmanage_35.scala 5315:45 stackmanage_35.scala 5348:34]
  wire  _GEN_2265 = pop_18 & empty_18 ? 1'h0 : _GEN_2247; // @[stackmanage_35.scala 5315:45 stackmanage_35.scala 5349:34]
  wire  _GEN_2266 = pop_18 & empty_18 ? 1'h0 : _GEN_2248; // @[stackmanage_35.scala 5315:45 stackmanage_35.scala 5350:34]
  wire  _GEN_2267 = pop_18 & empty_18 ? 1'h0 : _GEN_2249; // @[stackmanage_35.scala 5315:45 stackmanage_35.scala 5351:34]
  wire  _GEN_2270 = pop_17 & empty_17 ? 1'h0 : _T_371; // @[stackmanage_35.scala 5278:45 stackmanage_35.scala 5298:34]
  wire  _GEN_2271 = pop_17 & empty_17 ? 1'h0 : _GEN_2252; // @[stackmanage_35.scala 5278:45 stackmanage_35.scala 5299:34]
  wire  _GEN_2272 = pop_17 & empty_17 ? 1'h0 : _GEN_2253; // @[stackmanage_35.scala 5278:45 stackmanage_35.scala 5300:34]
  wire  _GEN_2273 = pop_17 & empty_17 ? 1'h0 : _GEN_2254; // @[stackmanage_35.scala 5278:45 stackmanage_35.scala 5301:34]
  wire  _GEN_2274 = pop_17 & empty_17 ? 1'h0 : _GEN_2255; // @[stackmanage_35.scala 5278:45 stackmanage_35.scala 5302:34]
  wire  _GEN_2275 = pop_17 & empty_17 ? 1'h0 : _GEN_2256; // @[stackmanage_35.scala 5278:45 stackmanage_35.scala 5303:34]
  wire  _GEN_2276 = pop_17 & empty_17 ? 1'h0 : _GEN_2257; // @[stackmanage_35.scala 5278:45 stackmanage_35.scala 5304:34]
  wire  _GEN_2277 = pop_17 & empty_17 ? 1'h0 : _GEN_2258; // @[stackmanage_35.scala 5278:45 stackmanage_35.scala 5305:34]
  wire  _GEN_2278 = pop_17 & empty_17 ? 1'h0 : _GEN_2259; // @[stackmanage_35.scala 5278:45 stackmanage_35.scala 5306:34]
  wire  _GEN_2279 = pop_17 & empty_17 ? 1'h0 : _GEN_2260; // @[stackmanage_35.scala 5278:45 stackmanage_35.scala 5307:34]
  wire  _GEN_2280 = pop_17 & empty_17 ? 1'h0 : _GEN_2261; // @[stackmanage_35.scala 5278:45 stackmanage_35.scala 5308:34]
  wire  _GEN_2281 = pop_17 & empty_17 ? 1'h0 : _GEN_2262; // @[stackmanage_35.scala 5278:45 stackmanage_35.scala 5309:34]
  wire  _GEN_2282 = pop_17 & empty_17 ? 1'h0 : _GEN_2263; // @[stackmanage_35.scala 5278:45 stackmanage_35.scala 5310:34]
  wire  _GEN_2283 = pop_17 & empty_17 ? 1'h0 : _GEN_2264; // @[stackmanage_35.scala 5278:45 stackmanage_35.scala 5311:34]
  wire  _GEN_2284 = pop_17 & empty_17 ? 1'h0 : _GEN_2265; // @[stackmanage_35.scala 5278:45 stackmanage_35.scala 5312:34]
  wire  _GEN_2285 = pop_17 & empty_17 ? 1'h0 : _GEN_2266; // @[stackmanage_35.scala 5278:45 stackmanage_35.scala 5313:34]
  wire  _GEN_2286 = pop_17 & empty_17 ? 1'h0 : _GEN_2267; // @[stackmanage_35.scala 5278:45 stackmanage_35.scala 5314:34]
  wire  _GEN_2289 = pop_16 & empty_16 ? 1'h0 : _T_368; // @[stackmanage_35.scala 5241:45 stackmanage_35.scala 5260:34]
  wire  _GEN_2290 = pop_16 & empty_16 ? 1'h0 : _GEN_2270; // @[stackmanage_35.scala 5241:45 stackmanage_35.scala 5261:34]
  wire  _GEN_2291 = pop_16 & empty_16 ? 1'h0 : _GEN_2271; // @[stackmanage_35.scala 5241:45 stackmanage_35.scala 5262:34]
  wire  _GEN_2292 = pop_16 & empty_16 ? 1'h0 : _GEN_2272; // @[stackmanage_35.scala 5241:45 stackmanage_35.scala 5263:34]
  wire  _GEN_2293 = pop_16 & empty_16 ? 1'h0 : _GEN_2273; // @[stackmanage_35.scala 5241:45 stackmanage_35.scala 5264:34]
  wire  _GEN_2294 = pop_16 & empty_16 ? 1'h0 : _GEN_2274; // @[stackmanage_35.scala 5241:45 stackmanage_35.scala 5265:34]
  wire  _GEN_2295 = pop_16 & empty_16 ? 1'h0 : _GEN_2275; // @[stackmanage_35.scala 5241:45 stackmanage_35.scala 5266:34]
  wire  _GEN_2296 = pop_16 & empty_16 ? 1'h0 : _GEN_2276; // @[stackmanage_35.scala 5241:45 stackmanage_35.scala 5267:34]
  wire  _GEN_2297 = pop_16 & empty_16 ? 1'h0 : _GEN_2277; // @[stackmanage_35.scala 5241:45 stackmanage_35.scala 5268:34]
  wire  _GEN_2298 = pop_16 & empty_16 ? 1'h0 : _GEN_2278; // @[stackmanage_35.scala 5241:45 stackmanage_35.scala 5269:34]
  wire  _GEN_2299 = pop_16 & empty_16 ? 1'h0 : _GEN_2279; // @[stackmanage_35.scala 5241:45 stackmanage_35.scala 5270:34]
  wire  _GEN_2300 = pop_16 & empty_16 ? 1'h0 : _GEN_2280; // @[stackmanage_35.scala 5241:45 stackmanage_35.scala 5271:34]
  wire  _GEN_2301 = pop_16 & empty_16 ? 1'h0 : _GEN_2281; // @[stackmanage_35.scala 5241:45 stackmanage_35.scala 5272:34]
  wire  _GEN_2302 = pop_16 & empty_16 ? 1'h0 : _GEN_2282; // @[stackmanage_35.scala 5241:45 stackmanage_35.scala 5273:34]
  wire  _GEN_2303 = pop_16 & empty_16 ? 1'h0 : _GEN_2283; // @[stackmanage_35.scala 5241:45 stackmanage_35.scala 5274:34]
  wire  _GEN_2304 = pop_16 & empty_16 ? 1'h0 : _GEN_2284; // @[stackmanage_35.scala 5241:45 stackmanage_35.scala 5275:34]
  wire  _GEN_2305 = pop_16 & empty_16 ? 1'h0 : _GEN_2285; // @[stackmanage_35.scala 5241:45 stackmanage_35.scala 5276:34]
  wire  _GEN_2306 = pop_16 & empty_16 ? 1'h0 : _GEN_2286; // @[stackmanage_35.scala 5241:45 stackmanage_35.scala 5277:34]
  wire  _GEN_2309 = pop_15 & empty_15 ? 1'h0 : _T_365; // @[stackmanage_35.scala 5204:45 stackmanage_35.scala 5222:34]
  wire  _GEN_2310 = pop_15 & empty_15 ? 1'h0 : _GEN_2289; // @[stackmanage_35.scala 5204:45 stackmanage_35.scala 5223:34]
  wire  _GEN_2311 = pop_15 & empty_15 ? 1'h0 : _GEN_2290; // @[stackmanage_35.scala 5204:45 stackmanage_35.scala 5224:34]
  wire  _GEN_2312 = pop_15 & empty_15 ? 1'h0 : _GEN_2291; // @[stackmanage_35.scala 5204:45 stackmanage_35.scala 5225:34]
  wire  _GEN_2313 = pop_15 & empty_15 ? 1'h0 : _GEN_2292; // @[stackmanage_35.scala 5204:45 stackmanage_35.scala 5226:34]
  wire  _GEN_2314 = pop_15 & empty_15 ? 1'h0 : _GEN_2293; // @[stackmanage_35.scala 5204:45 stackmanage_35.scala 5227:34]
  wire  _GEN_2315 = pop_15 & empty_15 ? 1'h0 : _GEN_2294; // @[stackmanage_35.scala 5204:45 stackmanage_35.scala 5228:34]
  wire  _GEN_2316 = pop_15 & empty_15 ? 1'h0 : _GEN_2295; // @[stackmanage_35.scala 5204:45 stackmanage_35.scala 5229:34]
  wire  _GEN_2317 = pop_15 & empty_15 ? 1'h0 : _GEN_2296; // @[stackmanage_35.scala 5204:45 stackmanage_35.scala 5230:34]
  wire  _GEN_2318 = pop_15 & empty_15 ? 1'h0 : _GEN_2297; // @[stackmanage_35.scala 5204:45 stackmanage_35.scala 5231:34]
  wire  _GEN_2319 = pop_15 & empty_15 ? 1'h0 : _GEN_2298; // @[stackmanage_35.scala 5204:45 stackmanage_35.scala 5232:34]
  wire  _GEN_2320 = pop_15 & empty_15 ? 1'h0 : _GEN_2299; // @[stackmanage_35.scala 5204:45 stackmanage_35.scala 5233:34]
  wire  _GEN_2321 = pop_15 & empty_15 ? 1'h0 : _GEN_2300; // @[stackmanage_35.scala 5204:45 stackmanage_35.scala 5234:34]
  wire  _GEN_2322 = pop_15 & empty_15 ? 1'h0 : _GEN_2301; // @[stackmanage_35.scala 5204:45 stackmanage_35.scala 5235:34]
  wire  _GEN_2323 = pop_15 & empty_15 ? 1'h0 : _GEN_2302; // @[stackmanage_35.scala 5204:45 stackmanage_35.scala 5236:34]
  wire  _GEN_2324 = pop_15 & empty_15 ? 1'h0 : _GEN_2303; // @[stackmanage_35.scala 5204:45 stackmanage_35.scala 5237:34]
  wire  _GEN_2325 = pop_15 & empty_15 ? 1'h0 : _GEN_2304; // @[stackmanage_35.scala 5204:45 stackmanage_35.scala 5238:34]
  wire  _GEN_2326 = pop_15 & empty_15 ? 1'h0 : _GEN_2305; // @[stackmanage_35.scala 5204:45 stackmanage_35.scala 5239:34]
  wire  _GEN_2327 = pop_15 & empty_15 ? 1'h0 : _GEN_2306; // @[stackmanage_35.scala 5204:45 stackmanage_35.scala 5240:34]
  wire  _GEN_2330 = pop_14 & empty_14 ? 1'h0 : _T_362; // @[stackmanage_35.scala 5167:45 stackmanage_35.scala 5184:34]
  wire  _GEN_2331 = pop_14 & empty_14 ? 1'h0 : _GEN_2309; // @[stackmanage_35.scala 5167:45 stackmanage_35.scala 5185:34]
  wire  _GEN_2332 = pop_14 & empty_14 ? 1'h0 : _GEN_2310; // @[stackmanage_35.scala 5167:45 stackmanage_35.scala 5186:34]
  wire  _GEN_2333 = pop_14 & empty_14 ? 1'h0 : _GEN_2311; // @[stackmanage_35.scala 5167:45 stackmanage_35.scala 5187:34]
  wire  _GEN_2334 = pop_14 & empty_14 ? 1'h0 : _GEN_2312; // @[stackmanage_35.scala 5167:45 stackmanage_35.scala 5188:34]
  wire  _GEN_2335 = pop_14 & empty_14 ? 1'h0 : _GEN_2313; // @[stackmanage_35.scala 5167:45 stackmanage_35.scala 5189:34]
  wire  _GEN_2336 = pop_14 & empty_14 ? 1'h0 : _GEN_2314; // @[stackmanage_35.scala 5167:45 stackmanage_35.scala 5190:34]
  wire  _GEN_2337 = pop_14 & empty_14 ? 1'h0 : _GEN_2315; // @[stackmanage_35.scala 5167:45 stackmanage_35.scala 5191:34]
  wire  _GEN_2338 = pop_14 & empty_14 ? 1'h0 : _GEN_2316; // @[stackmanage_35.scala 5167:45 stackmanage_35.scala 5192:34]
  wire  _GEN_2339 = pop_14 & empty_14 ? 1'h0 : _GEN_2317; // @[stackmanage_35.scala 5167:45 stackmanage_35.scala 5193:34]
  wire  _GEN_2340 = pop_14 & empty_14 ? 1'h0 : _GEN_2318; // @[stackmanage_35.scala 5167:45 stackmanage_35.scala 5194:34]
  wire  _GEN_2341 = pop_14 & empty_14 ? 1'h0 : _GEN_2319; // @[stackmanage_35.scala 5167:45 stackmanage_35.scala 5195:34]
  wire  _GEN_2342 = pop_14 & empty_14 ? 1'h0 : _GEN_2320; // @[stackmanage_35.scala 5167:45 stackmanage_35.scala 5196:34]
  wire  _GEN_2343 = pop_14 & empty_14 ? 1'h0 : _GEN_2321; // @[stackmanage_35.scala 5167:45 stackmanage_35.scala 5197:34]
  wire  _GEN_2344 = pop_14 & empty_14 ? 1'h0 : _GEN_2322; // @[stackmanage_35.scala 5167:45 stackmanage_35.scala 5198:34]
  wire  _GEN_2345 = pop_14 & empty_14 ? 1'h0 : _GEN_2323; // @[stackmanage_35.scala 5167:45 stackmanage_35.scala 5199:34]
  wire  _GEN_2346 = pop_14 & empty_14 ? 1'h0 : _GEN_2324; // @[stackmanage_35.scala 5167:45 stackmanage_35.scala 5200:34]
  wire  _GEN_2347 = pop_14 & empty_14 ? 1'h0 : _GEN_2325; // @[stackmanage_35.scala 5167:45 stackmanage_35.scala 5201:34]
  wire  _GEN_2348 = pop_14 & empty_14 ? 1'h0 : _GEN_2326; // @[stackmanage_35.scala 5167:45 stackmanage_35.scala 5202:34]
  wire  _GEN_2349 = pop_14 & empty_14 ? 1'h0 : _GEN_2327; // @[stackmanage_35.scala 5167:45 stackmanage_35.scala 5203:34]
  wire  _GEN_2352 = pop_13 & empty_13 ? 1'h0 : _T_359; // @[stackmanage_35.scala 5130:45 stackmanage_35.scala 5146:34]
  wire  _GEN_2353 = pop_13 & empty_13 ? 1'h0 : _GEN_2330; // @[stackmanage_35.scala 5130:45 stackmanage_35.scala 5147:34]
  wire  _GEN_2354 = pop_13 & empty_13 ? 1'h0 : _GEN_2331; // @[stackmanage_35.scala 5130:45 stackmanage_35.scala 5148:34]
  wire  _GEN_2355 = pop_13 & empty_13 ? 1'h0 : _GEN_2332; // @[stackmanage_35.scala 5130:45 stackmanage_35.scala 5149:34]
  wire  _GEN_2356 = pop_13 & empty_13 ? 1'h0 : _GEN_2333; // @[stackmanage_35.scala 5130:45 stackmanage_35.scala 5150:34]
  wire  _GEN_2357 = pop_13 & empty_13 ? 1'h0 : _GEN_2334; // @[stackmanage_35.scala 5130:45 stackmanage_35.scala 5151:34]
  wire  _GEN_2358 = pop_13 & empty_13 ? 1'h0 : _GEN_2335; // @[stackmanage_35.scala 5130:45 stackmanage_35.scala 5152:34]
  wire  _GEN_2359 = pop_13 & empty_13 ? 1'h0 : _GEN_2336; // @[stackmanage_35.scala 5130:45 stackmanage_35.scala 5153:34]
  wire  _GEN_2360 = pop_13 & empty_13 ? 1'h0 : _GEN_2337; // @[stackmanage_35.scala 5130:45 stackmanage_35.scala 5154:34]
  wire  _GEN_2361 = pop_13 & empty_13 ? 1'h0 : _GEN_2338; // @[stackmanage_35.scala 5130:45 stackmanage_35.scala 5155:34]
  wire  _GEN_2362 = pop_13 & empty_13 ? 1'h0 : _GEN_2339; // @[stackmanage_35.scala 5130:45 stackmanage_35.scala 5156:34]
  wire  _GEN_2363 = pop_13 & empty_13 ? 1'h0 : _GEN_2340; // @[stackmanage_35.scala 5130:45 stackmanage_35.scala 5157:34]
  wire  _GEN_2364 = pop_13 & empty_13 ? 1'h0 : _GEN_2341; // @[stackmanage_35.scala 5130:45 stackmanage_35.scala 5158:34]
  wire  _GEN_2365 = pop_13 & empty_13 ? 1'h0 : _GEN_2342; // @[stackmanage_35.scala 5130:45 stackmanage_35.scala 5159:34]
  wire  _GEN_2366 = pop_13 & empty_13 ? 1'h0 : _GEN_2343; // @[stackmanage_35.scala 5130:45 stackmanage_35.scala 5160:34]
  wire  _GEN_2367 = pop_13 & empty_13 ? 1'h0 : _GEN_2344; // @[stackmanage_35.scala 5130:45 stackmanage_35.scala 5161:34]
  wire  _GEN_2368 = pop_13 & empty_13 ? 1'h0 : _GEN_2345; // @[stackmanage_35.scala 5130:45 stackmanage_35.scala 5162:34]
  wire  _GEN_2369 = pop_13 & empty_13 ? 1'h0 : _GEN_2346; // @[stackmanage_35.scala 5130:45 stackmanage_35.scala 5163:34]
  wire  _GEN_2370 = pop_13 & empty_13 ? 1'h0 : _GEN_2347; // @[stackmanage_35.scala 5130:45 stackmanage_35.scala 5164:34]
  wire  _GEN_2371 = pop_13 & empty_13 ? 1'h0 : _GEN_2348; // @[stackmanage_35.scala 5130:45 stackmanage_35.scala 5165:34]
  wire  _GEN_2372 = pop_13 & empty_13 ? 1'h0 : _GEN_2349; // @[stackmanage_35.scala 5130:45 stackmanage_35.scala 5166:34]
  wire  _GEN_2375 = pop_12 & empty_12 ? 1'h0 : _T_356; // @[stackmanage_35.scala 5093:45 stackmanage_35.scala 5108:34]
  wire  _GEN_2376 = pop_12 & empty_12 ? 1'h0 : _GEN_2352; // @[stackmanage_35.scala 5093:45 stackmanage_35.scala 5109:34]
  wire  _GEN_2377 = pop_12 & empty_12 ? 1'h0 : _GEN_2353; // @[stackmanage_35.scala 5093:45 stackmanage_35.scala 5110:34]
  wire  _GEN_2378 = pop_12 & empty_12 ? 1'h0 : _GEN_2354; // @[stackmanage_35.scala 5093:45 stackmanage_35.scala 5111:34]
  wire  _GEN_2379 = pop_12 & empty_12 ? 1'h0 : _GEN_2355; // @[stackmanage_35.scala 5093:45 stackmanage_35.scala 5112:34]
  wire  _GEN_2380 = pop_12 & empty_12 ? 1'h0 : _GEN_2356; // @[stackmanage_35.scala 5093:45 stackmanage_35.scala 5113:34]
  wire  _GEN_2381 = pop_12 & empty_12 ? 1'h0 : _GEN_2357; // @[stackmanage_35.scala 5093:45 stackmanage_35.scala 5114:34]
  wire  _GEN_2382 = pop_12 & empty_12 ? 1'h0 : _GEN_2358; // @[stackmanage_35.scala 5093:45 stackmanage_35.scala 5115:34]
  wire  _GEN_2383 = pop_12 & empty_12 ? 1'h0 : _GEN_2359; // @[stackmanage_35.scala 5093:45 stackmanage_35.scala 5116:34]
  wire  _GEN_2384 = pop_12 & empty_12 ? 1'h0 : _GEN_2360; // @[stackmanage_35.scala 5093:45 stackmanage_35.scala 5117:34]
  wire  _GEN_2385 = pop_12 & empty_12 ? 1'h0 : _GEN_2361; // @[stackmanage_35.scala 5093:45 stackmanage_35.scala 5118:34]
  wire  _GEN_2386 = pop_12 & empty_12 ? 1'h0 : _GEN_2362; // @[stackmanage_35.scala 5093:45 stackmanage_35.scala 5119:34]
  wire  _GEN_2387 = pop_12 & empty_12 ? 1'h0 : _GEN_2363; // @[stackmanage_35.scala 5093:45 stackmanage_35.scala 5120:34]
  wire  _GEN_2388 = pop_12 & empty_12 ? 1'h0 : _GEN_2364; // @[stackmanage_35.scala 5093:45 stackmanage_35.scala 5121:34]
  wire  _GEN_2389 = pop_12 & empty_12 ? 1'h0 : _GEN_2365; // @[stackmanage_35.scala 5093:45 stackmanage_35.scala 5122:34]
  wire  _GEN_2390 = pop_12 & empty_12 ? 1'h0 : _GEN_2366; // @[stackmanage_35.scala 5093:45 stackmanage_35.scala 5123:34]
  wire  _GEN_2391 = pop_12 & empty_12 ? 1'h0 : _GEN_2367; // @[stackmanage_35.scala 5093:45 stackmanage_35.scala 5124:34]
  wire  _GEN_2392 = pop_12 & empty_12 ? 1'h0 : _GEN_2368; // @[stackmanage_35.scala 5093:45 stackmanage_35.scala 5125:34]
  wire  _GEN_2393 = pop_12 & empty_12 ? 1'h0 : _GEN_2369; // @[stackmanage_35.scala 5093:45 stackmanage_35.scala 5126:34]
  wire  _GEN_2394 = pop_12 & empty_12 ? 1'h0 : _GEN_2370; // @[stackmanage_35.scala 5093:45 stackmanage_35.scala 5127:34]
  wire  _GEN_2395 = pop_12 & empty_12 ? 1'h0 : _GEN_2371; // @[stackmanage_35.scala 5093:45 stackmanage_35.scala 5128:34]
  wire  _GEN_2396 = pop_12 & empty_12 ? 1'h0 : _GEN_2372; // @[stackmanage_35.scala 5093:45 stackmanage_35.scala 5129:34]
  wire  _GEN_2399 = pop_11 & empty_11 ? 1'h0 : _T_353; // @[stackmanage_35.scala 5056:45 stackmanage_35.scala 5070:34]
  wire  _GEN_2400 = pop_11 & empty_11 ? 1'h0 : _GEN_2375; // @[stackmanage_35.scala 5056:45 stackmanage_35.scala 5071:34]
  wire  _GEN_2401 = pop_11 & empty_11 ? 1'h0 : _GEN_2376; // @[stackmanage_35.scala 5056:45 stackmanage_35.scala 5072:34]
  wire  _GEN_2402 = pop_11 & empty_11 ? 1'h0 : _GEN_2377; // @[stackmanage_35.scala 5056:45 stackmanage_35.scala 5073:34]
  wire  _GEN_2403 = pop_11 & empty_11 ? 1'h0 : _GEN_2378; // @[stackmanage_35.scala 5056:45 stackmanage_35.scala 5074:34]
  wire  _GEN_2404 = pop_11 & empty_11 ? 1'h0 : _GEN_2379; // @[stackmanage_35.scala 5056:45 stackmanage_35.scala 5075:34]
  wire  _GEN_2405 = pop_11 & empty_11 ? 1'h0 : _GEN_2380; // @[stackmanage_35.scala 5056:45 stackmanage_35.scala 5076:34]
  wire  _GEN_2406 = pop_11 & empty_11 ? 1'h0 : _GEN_2381; // @[stackmanage_35.scala 5056:45 stackmanage_35.scala 5077:34]
  wire  _GEN_2407 = pop_11 & empty_11 ? 1'h0 : _GEN_2382; // @[stackmanage_35.scala 5056:45 stackmanage_35.scala 5078:34]
  wire  _GEN_2408 = pop_11 & empty_11 ? 1'h0 : _GEN_2383; // @[stackmanage_35.scala 5056:45 stackmanage_35.scala 5079:34]
  wire  _GEN_2409 = pop_11 & empty_11 ? 1'h0 : _GEN_2384; // @[stackmanage_35.scala 5056:45 stackmanage_35.scala 5080:34]
  wire  _GEN_2410 = pop_11 & empty_11 ? 1'h0 : _GEN_2385; // @[stackmanage_35.scala 5056:45 stackmanage_35.scala 5081:34]
  wire  _GEN_2411 = pop_11 & empty_11 ? 1'h0 : _GEN_2386; // @[stackmanage_35.scala 5056:45 stackmanage_35.scala 5082:34]
  wire  _GEN_2412 = pop_11 & empty_11 ? 1'h0 : _GEN_2387; // @[stackmanage_35.scala 5056:45 stackmanage_35.scala 5083:34]
  wire  _GEN_2413 = pop_11 & empty_11 ? 1'h0 : _GEN_2388; // @[stackmanage_35.scala 5056:45 stackmanage_35.scala 5084:34]
  wire  _GEN_2414 = pop_11 & empty_11 ? 1'h0 : _GEN_2389; // @[stackmanage_35.scala 5056:45 stackmanage_35.scala 5085:34]
  wire  _GEN_2415 = pop_11 & empty_11 ? 1'h0 : _GEN_2390; // @[stackmanage_35.scala 5056:45 stackmanage_35.scala 5086:34]
  wire  _GEN_2416 = pop_11 & empty_11 ? 1'h0 : _GEN_2391; // @[stackmanage_35.scala 5056:45 stackmanage_35.scala 5087:34]
  wire  _GEN_2417 = pop_11 & empty_11 ? 1'h0 : _GEN_2392; // @[stackmanage_35.scala 5056:45 stackmanage_35.scala 5088:34]
  wire  _GEN_2418 = pop_11 & empty_11 ? 1'h0 : _GEN_2393; // @[stackmanage_35.scala 5056:45 stackmanage_35.scala 5089:34]
  wire  _GEN_2419 = pop_11 & empty_11 ? 1'h0 : _GEN_2394; // @[stackmanage_35.scala 5056:45 stackmanage_35.scala 5090:34]
  wire  _GEN_2420 = pop_11 & empty_11 ? 1'h0 : _GEN_2395; // @[stackmanage_35.scala 5056:45 stackmanage_35.scala 5091:34]
  wire  _GEN_2421 = pop_11 & empty_11 ? 1'h0 : _GEN_2396; // @[stackmanage_35.scala 5056:45 stackmanage_35.scala 5092:34]
  wire  _GEN_2424 = pop_10 & empty_10 ? 1'h0 : _T_350; // @[stackmanage_35.scala 5019:45 stackmanage_35.scala 5032:34]
  wire  _GEN_2425 = pop_10 & empty_10 ? 1'h0 : _GEN_2399; // @[stackmanage_35.scala 5019:45 stackmanage_35.scala 5033:34]
  wire  _GEN_2426 = pop_10 & empty_10 ? 1'h0 : _GEN_2400; // @[stackmanage_35.scala 5019:45 stackmanage_35.scala 5034:34]
  wire  _GEN_2427 = pop_10 & empty_10 ? 1'h0 : _GEN_2401; // @[stackmanage_35.scala 5019:45 stackmanage_35.scala 5035:34]
  wire  _GEN_2428 = pop_10 & empty_10 ? 1'h0 : _GEN_2402; // @[stackmanage_35.scala 5019:45 stackmanage_35.scala 5036:34]
  wire  _GEN_2429 = pop_10 & empty_10 ? 1'h0 : _GEN_2403; // @[stackmanage_35.scala 5019:45 stackmanage_35.scala 5037:34]
  wire  _GEN_2430 = pop_10 & empty_10 ? 1'h0 : _GEN_2404; // @[stackmanage_35.scala 5019:45 stackmanage_35.scala 5038:34]
  wire  _GEN_2431 = pop_10 & empty_10 ? 1'h0 : _GEN_2405; // @[stackmanage_35.scala 5019:45 stackmanage_35.scala 5039:34]
  wire  _GEN_2432 = pop_10 & empty_10 ? 1'h0 : _GEN_2406; // @[stackmanage_35.scala 5019:45 stackmanage_35.scala 5040:34]
  wire  _GEN_2433 = pop_10 & empty_10 ? 1'h0 : _GEN_2407; // @[stackmanage_35.scala 5019:45 stackmanage_35.scala 5041:34]
  wire  _GEN_2434 = pop_10 & empty_10 ? 1'h0 : _GEN_2408; // @[stackmanage_35.scala 5019:45 stackmanage_35.scala 5042:34]
  wire  _GEN_2435 = pop_10 & empty_10 ? 1'h0 : _GEN_2409; // @[stackmanage_35.scala 5019:45 stackmanage_35.scala 5043:34]
  wire  _GEN_2436 = pop_10 & empty_10 ? 1'h0 : _GEN_2410; // @[stackmanage_35.scala 5019:45 stackmanage_35.scala 5044:34]
  wire  _GEN_2437 = pop_10 & empty_10 ? 1'h0 : _GEN_2411; // @[stackmanage_35.scala 5019:45 stackmanage_35.scala 5045:34]
  wire  _GEN_2438 = pop_10 & empty_10 ? 1'h0 : _GEN_2412; // @[stackmanage_35.scala 5019:45 stackmanage_35.scala 5046:34]
  wire  _GEN_2439 = pop_10 & empty_10 ? 1'h0 : _GEN_2413; // @[stackmanage_35.scala 5019:45 stackmanage_35.scala 5047:34]
  wire  _GEN_2440 = pop_10 & empty_10 ? 1'h0 : _GEN_2414; // @[stackmanage_35.scala 5019:45 stackmanage_35.scala 5048:34]
  wire  _GEN_2441 = pop_10 & empty_10 ? 1'h0 : _GEN_2415; // @[stackmanage_35.scala 5019:45 stackmanage_35.scala 5049:34]
  wire  _GEN_2442 = pop_10 & empty_10 ? 1'h0 : _GEN_2416; // @[stackmanage_35.scala 5019:45 stackmanage_35.scala 5050:34]
  wire  _GEN_2443 = pop_10 & empty_10 ? 1'h0 : _GEN_2417; // @[stackmanage_35.scala 5019:45 stackmanage_35.scala 5051:34]
  wire  _GEN_2444 = pop_10 & empty_10 ? 1'h0 : _GEN_2418; // @[stackmanage_35.scala 5019:45 stackmanage_35.scala 5052:34]
  wire  _GEN_2445 = pop_10 & empty_10 ? 1'h0 : _GEN_2419; // @[stackmanage_35.scala 5019:45 stackmanage_35.scala 5053:34]
  wire  _GEN_2446 = pop_10 & empty_10 ? 1'h0 : _GEN_2420; // @[stackmanage_35.scala 5019:45 stackmanage_35.scala 5054:34]
  wire  _GEN_2447 = pop_10 & empty_10 ? 1'h0 : _GEN_2421; // @[stackmanage_35.scala 5019:45 stackmanage_35.scala 5055:34]
  wire  _GEN_2450 = pop_9 & empty_9 ? 1'h0 : _T_347; // @[stackmanage_35.scala 4981:43 stackmanage_35.scala 4993:34]
  wire  _GEN_2451 = pop_9 & empty_9 ? 1'h0 : _GEN_2424; // @[stackmanage_35.scala 4981:43 stackmanage_35.scala 4994:34]
  wire  _GEN_2452 = pop_9 & empty_9 ? 1'h0 : _GEN_2425; // @[stackmanage_35.scala 4981:43 stackmanage_35.scala 4995:34]
  wire  _GEN_2453 = pop_9 & empty_9 ? 1'h0 : _GEN_2426; // @[stackmanage_35.scala 4981:43 stackmanage_35.scala 4996:34]
  wire  _GEN_2454 = pop_9 & empty_9 ? 1'h0 : _GEN_2427; // @[stackmanage_35.scala 4981:43 stackmanage_35.scala 4997:34]
  wire  _GEN_2455 = pop_9 & empty_9 ? 1'h0 : _GEN_2428; // @[stackmanage_35.scala 4981:43 stackmanage_35.scala 4998:34]
  wire  _GEN_2456 = pop_9 & empty_9 ? 1'h0 : _GEN_2429; // @[stackmanage_35.scala 4981:43 stackmanage_35.scala 4999:34]
  wire  _GEN_2457 = pop_9 & empty_9 ? 1'h0 : _GEN_2430; // @[stackmanage_35.scala 4981:43 stackmanage_35.scala 5000:34]
  wire  _GEN_2458 = pop_9 & empty_9 ? 1'h0 : _GEN_2431; // @[stackmanage_35.scala 4981:43 stackmanage_35.scala 5001:34]
  wire  _GEN_2459 = pop_9 & empty_9 ? 1'h0 : _GEN_2432; // @[stackmanage_35.scala 4981:43 stackmanage_35.scala 5002:34]
  wire  _GEN_2460 = pop_9 & empty_9 ? 1'h0 : _GEN_2433; // @[stackmanage_35.scala 4981:43 stackmanage_35.scala 5003:34]
  wire  _GEN_2461 = pop_9 & empty_9 ? 1'h0 : _GEN_2434; // @[stackmanage_35.scala 4981:43 stackmanage_35.scala 5004:34]
  wire  _GEN_2462 = pop_9 & empty_9 ? 1'h0 : _GEN_2435; // @[stackmanage_35.scala 4981:43 stackmanage_35.scala 5005:34]
  wire  _GEN_2463 = pop_9 & empty_9 ? 1'h0 : _GEN_2436; // @[stackmanage_35.scala 4981:43 stackmanage_35.scala 5006:34]
  wire  _GEN_2464 = pop_9 & empty_9 ? 1'h0 : _GEN_2437; // @[stackmanage_35.scala 4981:43 stackmanage_35.scala 5007:34]
  wire  _GEN_2465 = pop_9 & empty_9 ? 1'h0 : _GEN_2438; // @[stackmanage_35.scala 4981:43 stackmanage_35.scala 5008:34]
  wire  _GEN_2466 = pop_9 & empty_9 ? 1'h0 : _GEN_2439; // @[stackmanage_35.scala 4981:43 stackmanage_35.scala 5009:34]
  wire  _GEN_2467 = pop_9 & empty_9 ? 1'h0 : _GEN_2440; // @[stackmanage_35.scala 4981:43 stackmanage_35.scala 5010:34]
  wire  _GEN_2468 = pop_9 & empty_9 ? 1'h0 : _GEN_2441; // @[stackmanage_35.scala 4981:43 stackmanage_35.scala 5011:34]
  wire  _GEN_2469 = pop_9 & empty_9 ? 1'h0 : _GEN_2442; // @[stackmanage_35.scala 4981:43 stackmanage_35.scala 5012:34]
  wire  _GEN_2470 = pop_9 & empty_9 ? 1'h0 : _GEN_2443; // @[stackmanage_35.scala 4981:43 stackmanage_35.scala 5013:34]
  wire  _GEN_2471 = pop_9 & empty_9 ? 1'h0 : _GEN_2444; // @[stackmanage_35.scala 4981:43 stackmanage_35.scala 5014:34]
  wire  _GEN_2472 = pop_9 & empty_9 ? 1'h0 : _GEN_2445; // @[stackmanage_35.scala 4981:43 stackmanage_35.scala 5015:34]
  wire  _GEN_2473 = pop_9 & empty_9 ? 1'h0 : _GEN_2446; // @[stackmanage_35.scala 4981:43 stackmanage_35.scala 5016:34]
  wire  _GEN_2474 = pop_9 & empty_9 ? 1'h0 : _GEN_2447; // @[stackmanage_35.scala 4981:43 stackmanage_35.scala 5017:34]
  wire  _GEN_2477 = pop_8 & empty_8 ? 1'h0 : _T_344; // @[stackmanage_35.scala 4944:43 stackmanage_35.scala 4955:33]
  wire  _GEN_2478 = pop_8 & empty_8 ? 1'h0 : _GEN_2450; // @[stackmanage_35.scala 4944:43 stackmanage_35.scala 4956:34]
  wire  _GEN_2479 = pop_8 & empty_8 ? 1'h0 : _GEN_2451; // @[stackmanage_35.scala 4944:43 stackmanage_35.scala 4957:34]
  wire  _GEN_2480 = pop_8 & empty_8 ? 1'h0 : _GEN_2452; // @[stackmanage_35.scala 4944:43 stackmanage_35.scala 4958:34]
  wire  _GEN_2481 = pop_8 & empty_8 ? 1'h0 : _GEN_2453; // @[stackmanage_35.scala 4944:43 stackmanage_35.scala 4959:34]
  wire  _GEN_2482 = pop_8 & empty_8 ? 1'h0 : _GEN_2454; // @[stackmanage_35.scala 4944:43 stackmanage_35.scala 4960:34]
  wire  _GEN_2483 = pop_8 & empty_8 ? 1'h0 : _GEN_2455; // @[stackmanage_35.scala 4944:43 stackmanage_35.scala 4961:34]
  wire  _GEN_2484 = pop_8 & empty_8 ? 1'h0 : _GEN_2456; // @[stackmanage_35.scala 4944:43 stackmanage_35.scala 4962:34]
  wire  _GEN_2485 = pop_8 & empty_8 ? 1'h0 : _GEN_2457; // @[stackmanage_35.scala 4944:43 stackmanage_35.scala 4963:34]
  wire  _GEN_2486 = pop_8 & empty_8 ? 1'h0 : _GEN_2458; // @[stackmanage_35.scala 4944:43 stackmanage_35.scala 4964:34]
  wire  _GEN_2487 = pop_8 & empty_8 ? 1'h0 : _GEN_2459; // @[stackmanage_35.scala 4944:43 stackmanage_35.scala 4965:34]
  wire  _GEN_2488 = pop_8 & empty_8 ? 1'h0 : _GEN_2460; // @[stackmanage_35.scala 4944:43 stackmanage_35.scala 4966:34]
  wire  _GEN_2489 = pop_8 & empty_8 ? 1'h0 : _GEN_2461; // @[stackmanage_35.scala 4944:43 stackmanage_35.scala 4967:34]
  wire  _GEN_2490 = pop_8 & empty_8 ? 1'h0 : _GEN_2462; // @[stackmanage_35.scala 4944:43 stackmanage_35.scala 4968:34]
  wire  _GEN_2491 = pop_8 & empty_8 ? 1'h0 : _GEN_2463; // @[stackmanage_35.scala 4944:43 stackmanage_35.scala 4969:34]
  wire  _GEN_2492 = pop_8 & empty_8 ? 1'h0 : _GEN_2464; // @[stackmanage_35.scala 4944:43 stackmanage_35.scala 4970:34]
  wire  _GEN_2493 = pop_8 & empty_8 ? 1'h0 : _GEN_2465; // @[stackmanage_35.scala 4944:43 stackmanage_35.scala 4971:34]
  wire  _GEN_2494 = pop_8 & empty_8 ? 1'h0 : _GEN_2466; // @[stackmanage_35.scala 4944:43 stackmanage_35.scala 4972:34]
  wire  _GEN_2495 = pop_8 & empty_8 ? 1'h0 : _GEN_2467; // @[stackmanage_35.scala 4944:43 stackmanage_35.scala 4973:34]
  wire  _GEN_2496 = pop_8 & empty_8 ? 1'h0 : _GEN_2468; // @[stackmanage_35.scala 4944:43 stackmanage_35.scala 4974:34]
  wire  _GEN_2497 = pop_8 & empty_8 ? 1'h0 : _GEN_2469; // @[stackmanage_35.scala 4944:43 stackmanage_35.scala 4975:34]
  wire  _GEN_2498 = pop_8 & empty_8 ? 1'h0 : _GEN_2470; // @[stackmanage_35.scala 4944:43 stackmanage_35.scala 4976:34]
  wire  _GEN_2499 = pop_8 & empty_8 ? 1'h0 : _GEN_2471; // @[stackmanage_35.scala 4944:43 stackmanage_35.scala 4977:34]
  wire  _GEN_2500 = pop_8 & empty_8 ? 1'h0 : _GEN_2472; // @[stackmanage_35.scala 4944:43 stackmanage_35.scala 4978:34]
  wire  _GEN_2501 = pop_8 & empty_8 ? 1'h0 : _GEN_2473; // @[stackmanage_35.scala 4944:43 stackmanage_35.scala 4979:34]
  wire  _GEN_2502 = pop_8 & empty_8 ? 1'h0 : _GEN_2474; // @[stackmanage_35.scala 4944:43 stackmanage_35.scala 4980:34]
  wire  _GEN_2505 = pop_7 & empty_7 ? 1'h0 : _T_341; // @[stackmanage_35.scala 4906:43 stackmanage_35.scala 4916:33]
  wire  _GEN_2506 = pop_7 & empty_7 ? 1'h0 : _GEN_2477; // @[stackmanage_35.scala 4906:43 stackmanage_35.scala 4917:33]
  wire  _GEN_2507 = pop_7 & empty_7 ? 1'h0 : _GEN_2478; // @[stackmanage_35.scala 4906:43 stackmanage_35.scala 4918:34]
  wire  _GEN_2508 = pop_7 & empty_7 ? 1'h0 : _GEN_2479; // @[stackmanage_35.scala 4906:43 stackmanage_35.scala 4919:34]
  wire  _GEN_2509 = pop_7 & empty_7 ? 1'h0 : _GEN_2480; // @[stackmanage_35.scala 4906:43 stackmanage_35.scala 4920:34]
  wire  _GEN_2510 = pop_7 & empty_7 ? 1'h0 : _GEN_2481; // @[stackmanage_35.scala 4906:43 stackmanage_35.scala 4921:34]
  wire  _GEN_2511 = pop_7 & empty_7 ? 1'h0 : _GEN_2482; // @[stackmanage_35.scala 4906:43 stackmanage_35.scala 4922:34]
  wire  _GEN_2512 = pop_7 & empty_7 ? 1'h0 : _GEN_2483; // @[stackmanage_35.scala 4906:43 stackmanage_35.scala 4923:34]
  wire  _GEN_2513 = pop_7 & empty_7 ? 1'h0 : _GEN_2484; // @[stackmanage_35.scala 4906:43 stackmanage_35.scala 4924:34]
  wire  _GEN_2514 = pop_7 & empty_7 ? 1'h0 : _GEN_2485; // @[stackmanage_35.scala 4906:43 stackmanage_35.scala 4925:34]
  wire  _GEN_2515 = pop_7 & empty_7 ? 1'h0 : _GEN_2486; // @[stackmanage_35.scala 4906:43 stackmanage_35.scala 4926:34]
  wire  _GEN_2516 = pop_7 & empty_7 ? 1'h0 : _GEN_2487; // @[stackmanage_35.scala 4906:43 stackmanage_35.scala 4927:34]
  wire  _GEN_2517 = pop_7 & empty_7 ? 1'h0 : _GEN_2488; // @[stackmanage_35.scala 4906:43 stackmanage_35.scala 4928:34]
  wire  _GEN_2518 = pop_7 & empty_7 ? 1'h0 : _GEN_2489; // @[stackmanage_35.scala 4906:43 stackmanage_35.scala 4929:34]
  wire  _GEN_2519 = pop_7 & empty_7 ? 1'h0 : _GEN_2490; // @[stackmanage_35.scala 4906:43 stackmanage_35.scala 4930:34]
  wire  _GEN_2520 = pop_7 & empty_7 ? 1'h0 : _GEN_2491; // @[stackmanage_35.scala 4906:43 stackmanage_35.scala 4931:34]
  wire  _GEN_2521 = pop_7 & empty_7 ? 1'h0 : _GEN_2492; // @[stackmanage_35.scala 4906:43 stackmanage_35.scala 4932:34]
  wire  _GEN_2522 = pop_7 & empty_7 ? 1'h0 : _GEN_2493; // @[stackmanage_35.scala 4906:43 stackmanage_35.scala 4933:34]
  wire  _GEN_2523 = pop_7 & empty_7 ? 1'h0 : _GEN_2494; // @[stackmanage_35.scala 4906:43 stackmanage_35.scala 4934:34]
  wire  _GEN_2524 = pop_7 & empty_7 ? 1'h0 : _GEN_2495; // @[stackmanage_35.scala 4906:43 stackmanage_35.scala 4935:34]
  wire  _GEN_2525 = pop_7 & empty_7 ? 1'h0 : _GEN_2496; // @[stackmanage_35.scala 4906:43 stackmanage_35.scala 4936:34]
  wire  _GEN_2526 = pop_7 & empty_7 ? 1'h0 : _GEN_2497; // @[stackmanage_35.scala 4906:43 stackmanage_35.scala 4937:34]
  wire  _GEN_2527 = pop_7 & empty_7 ? 1'h0 : _GEN_2498; // @[stackmanage_35.scala 4906:43 stackmanage_35.scala 4938:34]
  wire  _GEN_2528 = pop_7 & empty_7 ? 1'h0 : _GEN_2499; // @[stackmanage_35.scala 4906:43 stackmanage_35.scala 4939:34]
  wire  _GEN_2529 = pop_7 & empty_7 ? 1'h0 : _GEN_2500; // @[stackmanage_35.scala 4906:43 stackmanage_35.scala 4940:34]
  wire  _GEN_2530 = pop_7 & empty_7 ? 1'h0 : _GEN_2501; // @[stackmanage_35.scala 4906:43 stackmanage_35.scala 4941:34]
  wire  _GEN_2531 = pop_7 & empty_7 ? 1'h0 : _GEN_2502; // @[stackmanage_35.scala 4906:43 stackmanage_35.scala 4942:34]
  wire  _GEN_2534 = pop_6 & empty_6 ? 1'h0 : _T_338; // @[stackmanage_35.scala 4868:43 stackmanage_35.scala 4877:33]
  wire  _GEN_2535 = pop_6 & empty_6 ? 1'h0 : _GEN_2505; // @[stackmanage_35.scala 4868:43 stackmanage_35.scala 4878:33]
  wire  _GEN_2536 = pop_6 & empty_6 ? 1'h0 : _GEN_2506; // @[stackmanage_35.scala 4868:43 stackmanage_35.scala 4879:33]
  wire  _GEN_2537 = pop_6 & empty_6 ? 1'h0 : _GEN_2507; // @[stackmanage_35.scala 4868:43 stackmanage_35.scala 4880:34]
  wire  _GEN_2538 = pop_6 & empty_6 ? 1'h0 : _GEN_2508; // @[stackmanage_35.scala 4868:43 stackmanage_35.scala 4881:34]
  wire  _GEN_2539 = pop_6 & empty_6 ? 1'h0 : _GEN_2509; // @[stackmanage_35.scala 4868:43 stackmanage_35.scala 4882:34]
  wire  _GEN_2540 = pop_6 & empty_6 ? 1'h0 : _GEN_2510; // @[stackmanage_35.scala 4868:43 stackmanage_35.scala 4883:34]
  wire  _GEN_2541 = pop_6 & empty_6 ? 1'h0 : _GEN_2511; // @[stackmanage_35.scala 4868:43 stackmanage_35.scala 4884:34]
  wire  _GEN_2542 = pop_6 & empty_6 ? 1'h0 : _GEN_2512; // @[stackmanage_35.scala 4868:43 stackmanage_35.scala 4885:34]
  wire  _GEN_2543 = pop_6 & empty_6 ? 1'h0 : _GEN_2513; // @[stackmanage_35.scala 4868:43 stackmanage_35.scala 4886:34]
  wire  _GEN_2544 = pop_6 & empty_6 ? 1'h0 : _GEN_2514; // @[stackmanage_35.scala 4868:43 stackmanage_35.scala 4887:34]
  wire  _GEN_2545 = pop_6 & empty_6 ? 1'h0 : _GEN_2515; // @[stackmanage_35.scala 4868:43 stackmanage_35.scala 4888:34]
  wire  _GEN_2546 = pop_6 & empty_6 ? 1'h0 : _GEN_2516; // @[stackmanage_35.scala 4868:43 stackmanage_35.scala 4889:34]
  wire  _GEN_2547 = pop_6 & empty_6 ? 1'h0 : _GEN_2517; // @[stackmanage_35.scala 4868:43 stackmanage_35.scala 4890:34]
  wire  _GEN_2548 = pop_6 & empty_6 ? 1'h0 : _GEN_2518; // @[stackmanage_35.scala 4868:43 stackmanage_35.scala 4891:34]
  wire  _GEN_2549 = pop_6 & empty_6 ? 1'h0 : _GEN_2519; // @[stackmanage_35.scala 4868:43 stackmanage_35.scala 4892:34]
  wire  _GEN_2550 = pop_6 & empty_6 ? 1'h0 : _GEN_2520; // @[stackmanage_35.scala 4868:43 stackmanage_35.scala 4893:34]
  wire  _GEN_2551 = pop_6 & empty_6 ? 1'h0 : _GEN_2521; // @[stackmanage_35.scala 4868:43 stackmanage_35.scala 4894:34]
  wire  _GEN_2552 = pop_6 & empty_6 ? 1'h0 : _GEN_2522; // @[stackmanage_35.scala 4868:43 stackmanage_35.scala 4895:34]
  wire  _GEN_2553 = pop_6 & empty_6 ? 1'h0 : _GEN_2523; // @[stackmanage_35.scala 4868:43 stackmanage_35.scala 4896:34]
  wire  _GEN_2554 = pop_6 & empty_6 ? 1'h0 : _GEN_2524; // @[stackmanage_35.scala 4868:43 stackmanage_35.scala 4897:34]
  wire  _GEN_2555 = pop_6 & empty_6 ? 1'h0 : _GEN_2525; // @[stackmanage_35.scala 4868:43 stackmanage_35.scala 4898:34]
  wire  _GEN_2556 = pop_6 & empty_6 ? 1'h0 : _GEN_2526; // @[stackmanage_35.scala 4868:43 stackmanage_35.scala 4899:34]
  wire  _GEN_2557 = pop_6 & empty_6 ? 1'h0 : _GEN_2527; // @[stackmanage_35.scala 4868:43 stackmanage_35.scala 4900:34]
  wire  _GEN_2558 = pop_6 & empty_6 ? 1'h0 : _GEN_2528; // @[stackmanage_35.scala 4868:43 stackmanage_35.scala 4901:34]
  wire  _GEN_2559 = pop_6 & empty_6 ? 1'h0 : _GEN_2529; // @[stackmanage_35.scala 4868:43 stackmanage_35.scala 4902:34]
  wire  _GEN_2560 = pop_6 & empty_6 ? 1'h0 : _GEN_2530; // @[stackmanage_35.scala 4868:43 stackmanage_35.scala 4903:34]
  wire  _GEN_2561 = pop_6 & empty_6 ? 1'h0 : _GEN_2531; // @[stackmanage_35.scala 4868:43 stackmanage_35.scala 4904:34]
  wire  _GEN_2564 = pop_5 & empty_5 ? 1'h0 : _T_335; // @[stackmanage_35.scala 4830:43 stackmanage_35.scala 4838:33]
  wire  _GEN_2565 = pop_5 & empty_5 ? 1'h0 : _GEN_2534; // @[stackmanage_35.scala 4830:43 stackmanage_35.scala 4839:33]
  wire  _GEN_2566 = pop_5 & empty_5 ? 1'h0 : _GEN_2535; // @[stackmanage_35.scala 4830:43 stackmanage_35.scala 4840:33]
  wire  _GEN_2567 = pop_5 & empty_5 ? 1'h0 : _GEN_2536; // @[stackmanage_35.scala 4830:43 stackmanage_35.scala 4841:33]
  wire  _GEN_2568 = pop_5 & empty_5 ? 1'h0 : _GEN_2537; // @[stackmanage_35.scala 4830:43 stackmanage_35.scala 4842:34]
  wire  _GEN_2569 = pop_5 & empty_5 ? 1'h0 : _GEN_2538; // @[stackmanage_35.scala 4830:43 stackmanage_35.scala 4843:34]
  wire  _GEN_2570 = pop_5 & empty_5 ? 1'h0 : _GEN_2539; // @[stackmanage_35.scala 4830:43 stackmanage_35.scala 4844:34]
  wire  _GEN_2571 = pop_5 & empty_5 ? 1'h0 : _GEN_2540; // @[stackmanage_35.scala 4830:43 stackmanage_35.scala 4845:34]
  wire  _GEN_2572 = pop_5 & empty_5 ? 1'h0 : _GEN_2541; // @[stackmanage_35.scala 4830:43 stackmanage_35.scala 4846:34]
  wire  _GEN_2573 = pop_5 & empty_5 ? 1'h0 : _GEN_2542; // @[stackmanage_35.scala 4830:43 stackmanage_35.scala 4847:34]
  wire  _GEN_2574 = pop_5 & empty_5 ? 1'h0 : _GEN_2543; // @[stackmanage_35.scala 4830:43 stackmanage_35.scala 4848:34]
  wire  _GEN_2575 = pop_5 & empty_5 ? 1'h0 : _GEN_2544; // @[stackmanage_35.scala 4830:43 stackmanage_35.scala 4849:34]
  wire  _GEN_2576 = pop_5 & empty_5 ? 1'h0 : _GEN_2545; // @[stackmanage_35.scala 4830:43 stackmanage_35.scala 4850:34]
  wire  _GEN_2577 = pop_5 & empty_5 ? 1'h0 : _GEN_2546; // @[stackmanage_35.scala 4830:43 stackmanage_35.scala 4851:34]
  wire  _GEN_2578 = pop_5 & empty_5 ? 1'h0 : _GEN_2547; // @[stackmanage_35.scala 4830:43 stackmanage_35.scala 4852:34]
  wire  _GEN_2579 = pop_5 & empty_5 ? 1'h0 : _GEN_2548; // @[stackmanage_35.scala 4830:43 stackmanage_35.scala 4853:34]
  wire  _GEN_2580 = pop_5 & empty_5 ? 1'h0 : _GEN_2549; // @[stackmanage_35.scala 4830:43 stackmanage_35.scala 4854:34]
  wire  _GEN_2581 = pop_5 & empty_5 ? 1'h0 : _GEN_2550; // @[stackmanage_35.scala 4830:43 stackmanage_35.scala 4855:34]
  wire  _GEN_2582 = pop_5 & empty_5 ? 1'h0 : _GEN_2551; // @[stackmanage_35.scala 4830:43 stackmanage_35.scala 4856:34]
  wire  _GEN_2583 = pop_5 & empty_5 ? 1'h0 : _GEN_2552; // @[stackmanage_35.scala 4830:43 stackmanage_35.scala 4857:34]
  wire  _GEN_2584 = pop_5 & empty_5 ? 1'h0 : _GEN_2553; // @[stackmanage_35.scala 4830:43 stackmanage_35.scala 4858:34]
  wire  _GEN_2585 = pop_5 & empty_5 ? 1'h0 : _GEN_2554; // @[stackmanage_35.scala 4830:43 stackmanage_35.scala 4859:34]
  wire  _GEN_2586 = pop_5 & empty_5 ? 1'h0 : _GEN_2555; // @[stackmanage_35.scala 4830:43 stackmanage_35.scala 4860:34]
  wire  _GEN_2587 = pop_5 & empty_5 ? 1'h0 : _GEN_2556; // @[stackmanage_35.scala 4830:43 stackmanage_35.scala 4861:34]
  wire  _GEN_2588 = pop_5 & empty_5 ? 1'h0 : _GEN_2557; // @[stackmanage_35.scala 4830:43 stackmanage_35.scala 4862:34]
  wire  _GEN_2589 = pop_5 & empty_5 ? 1'h0 : _GEN_2558; // @[stackmanage_35.scala 4830:43 stackmanage_35.scala 4863:34]
  wire  _GEN_2590 = pop_5 & empty_5 ? 1'h0 : _GEN_2559; // @[stackmanage_35.scala 4830:43 stackmanage_35.scala 4864:34]
  wire  _GEN_2591 = pop_5 & empty_5 ? 1'h0 : _GEN_2560; // @[stackmanage_35.scala 4830:43 stackmanage_35.scala 4865:34]
  wire  _GEN_2592 = pop_5 & empty_5 ? 1'h0 : _GEN_2561; // @[stackmanage_35.scala 4830:43 stackmanage_35.scala 4866:34]
  wire  _GEN_2595 = pop_4 & empty_4 ? 1'h0 : _T_332; // @[stackmanage_35.scala 4792:43 stackmanage_35.scala 4799:33]
  wire  _GEN_2596 = pop_4 & empty_4 ? 1'h0 : _GEN_2564; // @[stackmanage_35.scala 4792:43 stackmanage_35.scala 4800:33]
  wire  _GEN_2597 = pop_4 & empty_4 ? 1'h0 : _GEN_2565; // @[stackmanage_35.scala 4792:43 stackmanage_35.scala 4801:33]
  wire  _GEN_2598 = pop_4 & empty_4 ? 1'h0 : _GEN_2566; // @[stackmanage_35.scala 4792:43 stackmanage_35.scala 4802:33]
  wire  _GEN_2599 = pop_4 & empty_4 ? 1'h0 : _GEN_2567; // @[stackmanage_35.scala 4792:43 stackmanage_35.scala 4803:33]
  wire  _GEN_2600 = pop_4 & empty_4 ? 1'h0 : _GEN_2568; // @[stackmanage_35.scala 4792:43 stackmanage_35.scala 4804:34]
  wire  _GEN_2601 = pop_4 & empty_4 ? 1'h0 : _GEN_2569; // @[stackmanage_35.scala 4792:43 stackmanage_35.scala 4805:34]
  wire  _GEN_2602 = pop_4 & empty_4 ? 1'h0 : _GEN_2570; // @[stackmanage_35.scala 4792:43 stackmanage_35.scala 4806:34]
  wire  _GEN_2603 = pop_4 & empty_4 ? 1'h0 : _GEN_2571; // @[stackmanage_35.scala 4792:43 stackmanage_35.scala 4807:34]
  wire  _GEN_2604 = pop_4 & empty_4 ? 1'h0 : _GEN_2572; // @[stackmanage_35.scala 4792:43 stackmanage_35.scala 4808:34]
  wire  _GEN_2605 = pop_4 & empty_4 ? 1'h0 : _GEN_2573; // @[stackmanage_35.scala 4792:43 stackmanage_35.scala 4809:34]
  wire  _GEN_2606 = pop_4 & empty_4 ? 1'h0 : _GEN_2574; // @[stackmanage_35.scala 4792:43 stackmanage_35.scala 4810:34]
  wire  _GEN_2607 = pop_4 & empty_4 ? 1'h0 : _GEN_2575; // @[stackmanage_35.scala 4792:43 stackmanage_35.scala 4811:34]
  wire  _GEN_2608 = pop_4 & empty_4 ? 1'h0 : _GEN_2576; // @[stackmanage_35.scala 4792:43 stackmanage_35.scala 4812:34]
  wire  _GEN_2609 = pop_4 & empty_4 ? 1'h0 : _GEN_2577; // @[stackmanage_35.scala 4792:43 stackmanage_35.scala 4813:34]
  wire  _GEN_2610 = pop_4 & empty_4 ? 1'h0 : _GEN_2578; // @[stackmanage_35.scala 4792:43 stackmanage_35.scala 4814:34]
  wire  _GEN_2611 = pop_4 & empty_4 ? 1'h0 : _GEN_2579; // @[stackmanage_35.scala 4792:43 stackmanage_35.scala 4815:34]
  wire  _GEN_2612 = pop_4 & empty_4 ? 1'h0 : _GEN_2580; // @[stackmanage_35.scala 4792:43 stackmanage_35.scala 4816:34]
  wire  _GEN_2613 = pop_4 & empty_4 ? 1'h0 : _GEN_2581; // @[stackmanage_35.scala 4792:43 stackmanage_35.scala 4817:34]
  wire  _GEN_2614 = pop_4 & empty_4 ? 1'h0 : _GEN_2582; // @[stackmanage_35.scala 4792:43 stackmanage_35.scala 4818:34]
  wire  _GEN_2615 = pop_4 & empty_4 ? 1'h0 : _GEN_2583; // @[stackmanage_35.scala 4792:43 stackmanage_35.scala 4819:34]
  wire  _GEN_2616 = pop_4 & empty_4 ? 1'h0 : _GEN_2584; // @[stackmanage_35.scala 4792:43 stackmanage_35.scala 4820:34]
  wire  _GEN_2617 = pop_4 & empty_4 ? 1'h0 : _GEN_2585; // @[stackmanage_35.scala 4792:43 stackmanage_35.scala 4821:34]
  wire  _GEN_2618 = pop_4 & empty_4 ? 1'h0 : _GEN_2586; // @[stackmanage_35.scala 4792:43 stackmanage_35.scala 4822:34]
  wire  _GEN_2619 = pop_4 & empty_4 ? 1'h0 : _GEN_2587; // @[stackmanage_35.scala 4792:43 stackmanage_35.scala 4823:34]
  wire  _GEN_2620 = pop_4 & empty_4 ? 1'h0 : _GEN_2588; // @[stackmanage_35.scala 4792:43 stackmanage_35.scala 4824:34]
  wire  _GEN_2621 = pop_4 & empty_4 ? 1'h0 : _GEN_2589; // @[stackmanage_35.scala 4792:43 stackmanage_35.scala 4825:34]
  wire  _GEN_2622 = pop_4 & empty_4 ? 1'h0 : _GEN_2590; // @[stackmanage_35.scala 4792:43 stackmanage_35.scala 4826:34]
  wire  _GEN_2623 = pop_4 & empty_4 ? 1'h0 : _GEN_2591; // @[stackmanage_35.scala 4792:43 stackmanage_35.scala 4827:34]
  wire  _GEN_2624 = pop_4 & empty_4 ? 1'h0 : _GEN_2592; // @[stackmanage_35.scala 4792:43 stackmanage_35.scala 4828:34]
  wire  _GEN_2627 = pop_3 & empty_3 ? 1'h0 : _T_329; // @[stackmanage_35.scala 4754:43 stackmanage_35.scala 4760:33]
  wire  _GEN_2628 = pop_3 & empty_3 ? 1'h0 : _GEN_2595; // @[stackmanage_35.scala 4754:43 stackmanage_35.scala 4761:33]
  wire  _GEN_2629 = pop_3 & empty_3 ? 1'h0 : _GEN_2596; // @[stackmanage_35.scala 4754:43 stackmanage_35.scala 4762:33]
  wire  _GEN_2630 = pop_3 & empty_3 ? 1'h0 : _GEN_2597; // @[stackmanage_35.scala 4754:43 stackmanage_35.scala 4763:33]
  wire  _GEN_2631 = pop_3 & empty_3 ? 1'h0 : _GEN_2598; // @[stackmanage_35.scala 4754:43 stackmanage_35.scala 4764:33]
  wire  _GEN_2632 = pop_3 & empty_3 ? 1'h0 : _GEN_2599; // @[stackmanage_35.scala 4754:43 stackmanage_35.scala 4765:33]
  wire  _GEN_2633 = pop_3 & empty_3 ? 1'h0 : _GEN_2600; // @[stackmanage_35.scala 4754:43 stackmanage_35.scala 4766:34]
  wire  _GEN_2634 = pop_3 & empty_3 ? 1'h0 : _GEN_2601; // @[stackmanage_35.scala 4754:43 stackmanage_35.scala 4767:34]
  wire  _GEN_2635 = pop_3 & empty_3 ? 1'h0 : _GEN_2602; // @[stackmanage_35.scala 4754:43 stackmanage_35.scala 4768:34]
  wire  _GEN_2636 = pop_3 & empty_3 ? 1'h0 : _GEN_2603; // @[stackmanage_35.scala 4754:43 stackmanage_35.scala 4769:34]
  wire  _GEN_2637 = pop_3 & empty_3 ? 1'h0 : _GEN_2604; // @[stackmanage_35.scala 4754:43 stackmanage_35.scala 4770:34]
  wire  _GEN_2638 = pop_3 & empty_3 ? 1'h0 : _GEN_2605; // @[stackmanage_35.scala 4754:43 stackmanage_35.scala 4771:34]
  wire  _GEN_2639 = pop_3 & empty_3 ? 1'h0 : _GEN_2606; // @[stackmanage_35.scala 4754:43 stackmanage_35.scala 4772:34]
  wire  _GEN_2640 = pop_3 & empty_3 ? 1'h0 : _GEN_2607; // @[stackmanage_35.scala 4754:43 stackmanage_35.scala 4773:34]
  wire  _GEN_2641 = pop_3 & empty_3 ? 1'h0 : _GEN_2608; // @[stackmanage_35.scala 4754:43 stackmanage_35.scala 4774:34]
  wire  _GEN_2642 = pop_3 & empty_3 ? 1'h0 : _GEN_2609; // @[stackmanage_35.scala 4754:43 stackmanage_35.scala 4775:34]
  wire  _GEN_2643 = pop_3 & empty_3 ? 1'h0 : _GEN_2610; // @[stackmanage_35.scala 4754:43 stackmanage_35.scala 4776:34]
  wire  _GEN_2644 = pop_3 & empty_3 ? 1'h0 : _GEN_2611; // @[stackmanage_35.scala 4754:43 stackmanage_35.scala 4777:34]
  wire  _GEN_2645 = pop_3 & empty_3 ? 1'h0 : _GEN_2612; // @[stackmanage_35.scala 4754:43 stackmanage_35.scala 4778:34]
  wire  _GEN_2646 = pop_3 & empty_3 ? 1'h0 : _GEN_2613; // @[stackmanage_35.scala 4754:43 stackmanage_35.scala 4779:34]
  wire  _GEN_2647 = pop_3 & empty_3 ? 1'h0 : _GEN_2614; // @[stackmanage_35.scala 4754:43 stackmanage_35.scala 4780:34]
  wire  _GEN_2648 = pop_3 & empty_3 ? 1'h0 : _GEN_2615; // @[stackmanage_35.scala 4754:43 stackmanage_35.scala 4781:34]
  wire  _GEN_2649 = pop_3 & empty_3 ? 1'h0 : _GEN_2616; // @[stackmanage_35.scala 4754:43 stackmanage_35.scala 4782:34]
  wire  _GEN_2650 = pop_3 & empty_3 ? 1'h0 : _GEN_2617; // @[stackmanage_35.scala 4754:43 stackmanage_35.scala 4783:34]
  wire  _GEN_2651 = pop_3 & empty_3 ? 1'h0 : _GEN_2618; // @[stackmanage_35.scala 4754:43 stackmanage_35.scala 4784:34]
  wire  _GEN_2652 = pop_3 & empty_3 ? 1'h0 : _GEN_2619; // @[stackmanage_35.scala 4754:43 stackmanage_35.scala 4785:34]
  wire  _GEN_2653 = pop_3 & empty_3 ? 1'h0 : _GEN_2620; // @[stackmanage_35.scala 4754:43 stackmanage_35.scala 4786:34]
  wire  _GEN_2654 = pop_3 & empty_3 ? 1'h0 : _GEN_2621; // @[stackmanage_35.scala 4754:43 stackmanage_35.scala 4787:34]
  wire  _GEN_2655 = pop_3 & empty_3 ? 1'h0 : _GEN_2622; // @[stackmanage_35.scala 4754:43 stackmanage_35.scala 4788:34]
  wire  _GEN_2656 = pop_3 & empty_3 ? 1'h0 : _GEN_2623; // @[stackmanage_35.scala 4754:43 stackmanage_35.scala 4789:34]
  wire  _GEN_2657 = pop_3 & empty_3 ? 1'h0 : _GEN_2624; // @[stackmanage_35.scala 4754:43 stackmanage_35.scala 4790:34]
  wire  _T_468 = dispatch_0 | dispatch_1 | dispatch_2 | dispatch_3 | dispatch_4 | dispatch_5 | dispatch_6 | dispatch_7
     | dispatch_8 | dispatch_9 | dispatch_10 | dispatch_11 | dispatch_12 | dispatch_13 | dispatch_14 | dispatch_15 |
    dispatch_16 | dispatch_17 | dispatch_18 | dispatch_19 | dispatch_20 | dispatch_21 | dispatch_22 | dispatch_23 |
    dispatch_24; // @[stackmanage_35.scala 5988:538]
  wire  _T_514 = Stack_0_io_empty & Stack_1_io_empty & Stack_2_io_empty & Stack_3_io_empty & Stack_4_io_empty &
    Stack_5_io_empty & Stack_6_io_empty & Stack_7_io_empty & Stack_8_io_empty & Stack_9_io_empty & Stack_10_io_empty &
    Stack_11_io_empty & Stack_12_io_empty & Stack_13_io_empty & Stack_14_io_empty & Stack_15_io_empty &
    Stack_16_io_empty & Stack_17_io_empty & Stack_18_io_empty & Stack_19_io_empty & Stack_20_io_empty &
    Stack_21_io_empty & Stack_22_io_empty & Stack_23_io_empty & Stack_24_io_empty; // @[stackmanage_35.scala 5990:496]
  LUT LUT_stack ( // @[stackmanage_35.scala 35:45]
    .clock(LUT_stack_clock),
    .reset(LUT_stack_reset),
    .io_push(LUT_stack_io_push),
    .io_push_valid(LUT_stack_io_push_valid),
    .io_pop(LUT_stack_io_pop),
    .io_pop_valid(LUT_stack_io_pop_valid),
    .io_clear(LUT_stack_io_clear),
    .io_empty_0(LUT_stack_io_empty_0),
    .io_empty_1(LUT_stack_io_empty_1),
    .io_empty_2(LUT_stack_io_empty_2),
    .io_empty_3(LUT_stack_io_empty_3),
    .io_empty_4(LUT_stack_io_empty_4),
    .io_empty_5(LUT_stack_io_empty_5),
    .io_empty_6(LUT_stack_io_empty_6),
    .io_empty_7(LUT_stack_io_empty_7),
    .io_empty_8(LUT_stack_io_empty_8),
    .io_empty_9(LUT_stack_io_empty_9),
    .io_empty_10(LUT_stack_io_empty_10),
    .io_empty_11(LUT_stack_io_empty_11),
    .io_empty_12(LUT_stack_io_empty_12),
    .io_empty_13(LUT_stack_io_empty_13),
    .io_empty_14(LUT_stack_io_empty_14),
    .io_empty_15(LUT_stack_io_empty_15),
    .io_empty_16(LUT_stack_io_empty_16),
    .io_empty_17(LUT_stack_io_empty_17),
    .io_empty_18(LUT_stack_io_empty_18),
    .io_empty_19(LUT_stack_io_empty_19),
    .io_empty_20(LUT_stack_io_empty_20),
    .io_empty_21(LUT_stack_io_empty_21),
    .io_empty_22(LUT_stack_io_empty_22),
    .io_empty_23(LUT_stack_io_empty_23),
    .io_empty_24(LUT_stack_io_empty_24),
    .io_empty_25(LUT_stack_io_empty_25),
    .io_empty_26(LUT_stack_io_empty_26),
    .io_empty_27(LUT_stack_io_empty_27),
    .io_empty_28(LUT_stack_io_empty_28),
    .io_empty_29(LUT_stack_io_empty_29),
    .io_empty_30(LUT_stack_io_empty_30),
    .io_empty_31(LUT_stack_io_empty_31),
    .io_empty_32(LUT_stack_io_empty_32),
    .io_empty_33(LUT_stack_io_empty_33),
    .io_empty_34(LUT_stack_io_empty_34),
    .io_dispatch_0(LUT_stack_io_dispatch_0),
    .io_dispatch_1(LUT_stack_io_dispatch_1),
    .io_dispatch_2(LUT_stack_io_dispatch_2),
    .io_dispatch_3(LUT_stack_io_dispatch_3),
    .io_dispatch_4(LUT_stack_io_dispatch_4),
    .io_dispatch_5(LUT_stack_io_dispatch_5),
    .io_dispatch_6(LUT_stack_io_dispatch_6),
    .io_dispatch_7(LUT_stack_io_dispatch_7),
    .io_dispatch_8(LUT_stack_io_dispatch_8),
    .io_dispatch_9(LUT_stack_io_dispatch_9),
    .io_dispatch_10(LUT_stack_io_dispatch_10),
    .io_dispatch_11(LUT_stack_io_dispatch_11),
    .io_dispatch_12(LUT_stack_io_dispatch_12),
    .io_dispatch_13(LUT_stack_io_dispatch_13),
    .io_dispatch_14(LUT_stack_io_dispatch_14),
    .io_dispatch_15(LUT_stack_io_dispatch_15),
    .io_dispatch_16(LUT_stack_io_dispatch_16),
    .io_dispatch_17(LUT_stack_io_dispatch_17),
    .io_dispatch_18(LUT_stack_io_dispatch_18),
    .io_dispatch_19(LUT_stack_io_dispatch_19),
    .io_dispatch_20(LUT_stack_io_dispatch_20),
    .io_dispatch_21(LUT_stack_io_dispatch_21),
    .io_dispatch_22(LUT_stack_io_dispatch_22),
    .io_dispatch_23(LUT_stack_io_dispatch_23),
    .io_dispatch_24(LUT_stack_io_dispatch_24),
    .io_dispatch_25(LUT_stack_io_dispatch_25),
    .io_dispatch_26(LUT_stack_io_dispatch_26),
    .io_dispatch_27(LUT_stack_io_dispatch_27),
    .io_dispatch_28(LUT_stack_io_dispatch_28),
    .io_dispatch_29(LUT_stack_io_dispatch_29),
    .io_dispatch_30(LUT_stack_io_dispatch_30),
    .io_dispatch_31(LUT_stack_io_dispatch_31),
    .io_dispatch_32(LUT_stack_io_dispatch_32),
    .io_dispatch_33(LUT_stack_io_dispatch_33),
    .io_dispatch_34(LUT_stack_io_dispatch_34),
    .io_ray_id_push(LUT_stack_io_ray_id_push),
    .io_ray_id_pop(LUT_stack_io_ray_id_pop),
    .io_node_id_push_in(LUT_stack_io_node_id_push_in),
    .io_hitT_in(LUT_stack_io_hitT_in),
    .io_ray_id_pop_out(LUT_stack_io_ray_id_pop_out),
    .io_hitT_out(LUT_stack_io_hitT_out),
    .io_pop_0(LUT_stack_io_pop_0),
    .io_pop_1(LUT_stack_io_pop_1),
    .io_pop_2(LUT_stack_io_pop_2),
    .io_pop_3(LUT_stack_io_pop_3),
    .io_pop_4(LUT_stack_io_pop_4),
    .io_pop_5(LUT_stack_io_pop_5),
    .io_pop_6(LUT_stack_io_pop_6),
    .io_pop_7(LUT_stack_io_pop_7),
    .io_pop_8(LUT_stack_io_pop_8),
    .io_pop_9(LUT_stack_io_pop_9),
    .io_pop_10(LUT_stack_io_pop_10),
    .io_pop_11(LUT_stack_io_pop_11),
    .io_pop_12(LUT_stack_io_pop_12),
    .io_pop_13(LUT_stack_io_pop_13),
    .io_pop_14(LUT_stack_io_pop_14),
    .io_pop_15(LUT_stack_io_pop_15),
    .io_pop_16(LUT_stack_io_pop_16),
    .io_pop_17(LUT_stack_io_pop_17),
    .io_pop_18(LUT_stack_io_pop_18),
    .io_pop_19(LUT_stack_io_pop_19),
    .io_pop_20(LUT_stack_io_pop_20),
    .io_pop_21(LUT_stack_io_pop_21),
    .io_pop_22(LUT_stack_io_pop_22),
    .io_pop_23(LUT_stack_io_pop_23),
    .io_pop_24(LUT_stack_io_pop_24),
    .io_pop_25(LUT_stack_io_pop_25),
    .io_pop_26(LUT_stack_io_pop_26),
    .io_pop_27(LUT_stack_io_pop_27),
    .io_pop_28(LUT_stack_io_pop_28),
    .io_pop_29(LUT_stack_io_pop_29),
    .io_pop_30(LUT_stack_io_pop_30),
    .io_pop_31(LUT_stack_io_pop_31),
    .io_pop_32(LUT_stack_io_pop_32),
    .io_pop_33(LUT_stack_io_pop_33),
    .io_pop_34(LUT_stack_io_pop_34),
    .io_pop_en(LUT_stack_io_pop_en),
    .io_push_0(LUT_stack_io_push_0),
    .io_push_1(LUT_stack_io_push_1),
    .io_push_2(LUT_stack_io_push_2),
    .io_push_3(LUT_stack_io_push_3),
    .io_push_4(LUT_stack_io_push_4),
    .io_push_5(LUT_stack_io_push_5),
    .io_push_6(LUT_stack_io_push_6),
    .io_push_7(LUT_stack_io_push_7),
    .io_push_8(LUT_stack_io_push_8),
    .io_push_9(LUT_stack_io_push_9),
    .io_push_10(LUT_stack_io_push_10),
    .io_push_11(LUT_stack_io_push_11),
    .io_push_12(LUT_stack_io_push_12),
    .io_push_13(LUT_stack_io_push_13),
    .io_push_14(LUT_stack_io_push_14),
    .io_push_15(LUT_stack_io_push_15),
    .io_push_16(LUT_stack_io_push_16),
    .io_push_17(LUT_stack_io_push_17),
    .io_push_18(LUT_stack_io_push_18),
    .io_push_19(LUT_stack_io_push_19),
    .io_push_20(LUT_stack_io_push_20),
    .io_push_21(LUT_stack_io_push_21),
    .io_push_22(LUT_stack_io_push_22),
    .io_push_23(LUT_stack_io_push_23),
    .io_push_24(LUT_stack_io_push_24),
    .io_push_25(LUT_stack_io_push_25),
    .io_push_26(LUT_stack_io_push_26),
    .io_push_27(LUT_stack_io_push_27),
    .io_push_28(LUT_stack_io_push_28),
    .io_push_29(LUT_stack_io_push_29),
    .io_push_30(LUT_stack_io_push_30),
    .io_push_31(LUT_stack_io_push_31),
    .io_push_32(LUT_stack_io_push_32),
    .io_push_33(LUT_stack_io_push_33),
    .io_push_34(LUT_stack_io_push_34),
    .io_clear_0(LUT_stack_io_clear_0),
    .io_clear_1(LUT_stack_io_clear_1),
    .io_clear_2(LUT_stack_io_clear_2),
    .io_clear_3(LUT_stack_io_clear_3),
    .io_clear_4(LUT_stack_io_clear_4),
    .io_clear_5(LUT_stack_io_clear_5),
    .io_clear_6(LUT_stack_io_clear_6),
    .io_clear_7(LUT_stack_io_clear_7),
    .io_clear_8(LUT_stack_io_clear_8),
    .io_clear_9(LUT_stack_io_clear_9),
    .io_clear_10(LUT_stack_io_clear_10),
    .io_clear_11(LUT_stack_io_clear_11),
    .io_clear_12(LUT_stack_io_clear_12),
    .io_clear_13(LUT_stack_io_clear_13),
    .io_clear_14(LUT_stack_io_clear_14),
    .io_clear_15(LUT_stack_io_clear_15),
    .io_clear_16(LUT_stack_io_clear_16),
    .io_clear_17(LUT_stack_io_clear_17),
    .io_clear_18(LUT_stack_io_clear_18),
    .io_clear_19(LUT_stack_io_clear_19),
    .io_clear_20(LUT_stack_io_clear_20),
    .io_clear_21(LUT_stack_io_clear_21),
    .io_clear_22(LUT_stack_io_clear_22),
    .io_clear_23(LUT_stack_io_clear_23),
    .io_clear_24(LUT_stack_io_clear_24),
    .io_clear_25(LUT_stack_io_clear_25),
    .io_clear_26(LUT_stack_io_clear_26),
    .io_clear_27(LUT_stack_io_clear_27),
    .io_clear_28(LUT_stack_io_clear_28),
    .io_clear_29(LUT_stack_io_clear_29),
    .io_clear_30(LUT_stack_io_clear_30),
    .io_clear_31(LUT_stack_io_clear_31),
    .io_clear_32(LUT_stack_io_clear_32),
    .io_clear_33(LUT_stack_io_clear_33),
    .io_clear_34(LUT_stack_io_clear_34),
    .io_push_en(LUT_stack_io_push_en),
    .io_no_match(LUT_stack_io_no_match)
  );
  Stack Stack_0 ( // @[stackmanage_35.scala 36:48]
    .clock(Stack_0_clock),
    .reset(Stack_0_reset),
    .io_push(Stack_0_io_push),
    .io_pop(Stack_0_io_pop),
    .io_dataIn(Stack_0_io_dataIn),
    .io_clear(Stack_0_io_clear),
    .io_ray_id(Stack_0_io_ray_id),
    .io_dataOut(Stack_0_io_dataOut),
    .io_empty(Stack_0_io_empty),
    .io_hit_in(Stack_0_io_hit_in),
    .io_hit_out(Stack_0_io_hit_out),
    .io_ray_out(Stack_0_io_ray_out),
    .io_enable(Stack_0_io_enable)
  );
  Stack Stack_1 ( // @[stackmanage_35.scala 37:48]
    .clock(Stack_1_clock),
    .reset(Stack_1_reset),
    .io_push(Stack_1_io_push),
    .io_pop(Stack_1_io_pop),
    .io_dataIn(Stack_1_io_dataIn),
    .io_clear(Stack_1_io_clear),
    .io_ray_id(Stack_1_io_ray_id),
    .io_dataOut(Stack_1_io_dataOut),
    .io_empty(Stack_1_io_empty),
    .io_hit_in(Stack_1_io_hit_in),
    .io_hit_out(Stack_1_io_hit_out),
    .io_ray_out(Stack_1_io_ray_out),
    .io_enable(Stack_1_io_enable)
  );
  Stack Stack_2 ( // @[stackmanage_35.scala 38:48]
    .clock(Stack_2_clock),
    .reset(Stack_2_reset),
    .io_push(Stack_2_io_push),
    .io_pop(Stack_2_io_pop),
    .io_dataIn(Stack_2_io_dataIn),
    .io_clear(Stack_2_io_clear),
    .io_ray_id(Stack_2_io_ray_id),
    .io_dataOut(Stack_2_io_dataOut),
    .io_empty(Stack_2_io_empty),
    .io_hit_in(Stack_2_io_hit_in),
    .io_hit_out(Stack_2_io_hit_out),
    .io_ray_out(Stack_2_io_ray_out),
    .io_enable(Stack_2_io_enable)
  );
  Stack Stack_3 ( // @[stackmanage_35.scala 39:48]
    .clock(Stack_3_clock),
    .reset(Stack_3_reset),
    .io_push(Stack_3_io_push),
    .io_pop(Stack_3_io_pop),
    .io_dataIn(Stack_3_io_dataIn),
    .io_clear(Stack_3_io_clear),
    .io_ray_id(Stack_3_io_ray_id),
    .io_dataOut(Stack_3_io_dataOut),
    .io_empty(Stack_3_io_empty),
    .io_hit_in(Stack_3_io_hit_in),
    .io_hit_out(Stack_3_io_hit_out),
    .io_ray_out(Stack_3_io_ray_out),
    .io_enable(Stack_3_io_enable)
  );
  Stack Stack_4 ( // @[stackmanage_35.scala 40:48]
    .clock(Stack_4_clock),
    .reset(Stack_4_reset),
    .io_push(Stack_4_io_push),
    .io_pop(Stack_4_io_pop),
    .io_dataIn(Stack_4_io_dataIn),
    .io_clear(Stack_4_io_clear),
    .io_ray_id(Stack_4_io_ray_id),
    .io_dataOut(Stack_4_io_dataOut),
    .io_empty(Stack_4_io_empty),
    .io_hit_in(Stack_4_io_hit_in),
    .io_hit_out(Stack_4_io_hit_out),
    .io_ray_out(Stack_4_io_ray_out),
    .io_enable(Stack_4_io_enable)
  );
  Stack Stack_5 ( // @[stackmanage_35.scala 41:48]
    .clock(Stack_5_clock),
    .reset(Stack_5_reset),
    .io_push(Stack_5_io_push),
    .io_pop(Stack_5_io_pop),
    .io_dataIn(Stack_5_io_dataIn),
    .io_clear(Stack_5_io_clear),
    .io_ray_id(Stack_5_io_ray_id),
    .io_dataOut(Stack_5_io_dataOut),
    .io_empty(Stack_5_io_empty),
    .io_hit_in(Stack_5_io_hit_in),
    .io_hit_out(Stack_5_io_hit_out),
    .io_ray_out(Stack_5_io_ray_out),
    .io_enable(Stack_5_io_enable)
  );
  Stack Stack_6 ( // @[stackmanage_35.scala 42:48]
    .clock(Stack_6_clock),
    .reset(Stack_6_reset),
    .io_push(Stack_6_io_push),
    .io_pop(Stack_6_io_pop),
    .io_dataIn(Stack_6_io_dataIn),
    .io_clear(Stack_6_io_clear),
    .io_ray_id(Stack_6_io_ray_id),
    .io_dataOut(Stack_6_io_dataOut),
    .io_empty(Stack_6_io_empty),
    .io_hit_in(Stack_6_io_hit_in),
    .io_hit_out(Stack_6_io_hit_out),
    .io_ray_out(Stack_6_io_ray_out),
    .io_enable(Stack_6_io_enable)
  );
  Stack Stack_7 ( // @[stackmanage_35.scala 43:48]
    .clock(Stack_7_clock),
    .reset(Stack_7_reset),
    .io_push(Stack_7_io_push),
    .io_pop(Stack_7_io_pop),
    .io_dataIn(Stack_7_io_dataIn),
    .io_clear(Stack_7_io_clear),
    .io_ray_id(Stack_7_io_ray_id),
    .io_dataOut(Stack_7_io_dataOut),
    .io_empty(Stack_7_io_empty),
    .io_hit_in(Stack_7_io_hit_in),
    .io_hit_out(Stack_7_io_hit_out),
    .io_ray_out(Stack_7_io_ray_out),
    .io_enable(Stack_7_io_enable)
  );
  Stack Stack_8 ( // @[stackmanage_35.scala 44:48]
    .clock(Stack_8_clock),
    .reset(Stack_8_reset),
    .io_push(Stack_8_io_push),
    .io_pop(Stack_8_io_pop),
    .io_dataIn(Stack_8_io_dataIn),
    .io_clear(Stack_8_io_clear),
    .io_ray_id(Stack_8_io_ray_id),
    .io_dataOut(Stack_8_io_dataOut),
    .io_empty(Stack_8_io_empty),
    .io_hit_in(Stack_8_io_hit_in),
    .io_hit_out(Stack_8_io_hit_out),
    .io_ray_out(Stack_8_io_ray_out),
    .io_enable(Stack_8_io_enable)
  );
  Stack Stack_9 ( // @[stackmanage_35.scala 45:48]
    .clock(Stack_9_clock),
    .reset(Stack_9_reset),
    .io_push(Stack_9_io_push),
    .io_pop(Stack_9_io_pop),
    .io_dataIn(Stack_9_io_dataIn),
    .io_clear(Stack_9_io_clear),
    .io_ray_id(Stack_9_io_ray_id),
    .io_dataOut(Stack_9_io_dataOut),
    .io_empty(Stack_9_io_empty),
    .io_hit_in(Stack_9_io_hit_in),
    .io_hit_out(Stack_9_io_hit_out),
    .io_ray_out(Stack_9_io_ray_out),
    .io_enable(Stack_9_io_enable)
  );
  Stack Stack_10 ( // @[stackmanage_35.scala 46:47]
    .clock(Stack_10_clock),
    .reset(Stack_10_reset),
    .io_push(Stack_10_io_push),
    .io_pop(Stack_10_io_pop),
    .io_dataIn(Stack_10_io_dataIn),
    .io_clear(Stack_10_io_clear),
    .io_ray_id(Stack_10_io_ray_id),
    .io_dataOut(Stack_10_io_dataOut),
    .io_empty(Stack_10_io_empty),
    .io_hit_in(Stack_10_io_hit_in),
    .io_hit_out(Stack_10_io_hit_out),
    .io_ray_out(Stack_10_io_ray_out),
    .io_enable(Stack_10_io_enable)
  );
  Stack Stack_11 ( // @[stackmanage_35.scala 47:47]
    .clock(Stack_11_clock),
    .reset(Stack_11_reset),
    .io_push(Stack_11_io_push),
    .io_pop(Stack_11_io_pop),
    .io_dataIn(Stack_11_io_dataIn),
    .io_clear(Stack_11_io_clear),
    .io_ray_id(Stack_11_io_ray_id),
    .io_dataOut(Stack_11_io_dataOut),
    .io_empty(Stack_11_io_empty),
    .io_hit_in(Stack_11_io_hit_in),
    .io_hit_out(Stack_11_io_hit_out),
    .io_ray_out(Stack_11_io_ray_out),
    .io_enable(Stack_11_io_enable)
  );
  Stack Stack_12 ( // @[stackmanage_35.scala 48:47]
    .clock(Stack_12_clock),
    .reset(Stack_12_reset),
    .io_push(Stack_12_io_push),
    .io_pop(Stack_12_io_pop),
    .io_dataIn(Stack_12_io_dataIn),
    .io_clear(Stack_12_io_clear),
    .io_ray_id(Stack_12_io_ray_id),
    .io_dataOut(Stack_12_io_dataOut),
    .io_empty(Stack_12_io_empty),
    .io_hit_in(Stack_12_io_hit_in),
    .io_hit_out(Stack_12_io_hit_out),
    .io_ray_out(Stack_12_io_ray_out),
    .io_enable(Stack_12_io_enable)
  );
  Stack Stack_13 ( // @[stackmanage_35.scala 49:47]
    .clock(Stack_13_clock),
    .reset(Stack_13_reset),
    .io_push(Stack_13_io_push),
    .io_pop(Stack_13_io_pop),
    .io_dataIn(Stack_13_io_dataIn),
    .io_clear(Stack_13_io_clear),
    .io_ray_id(Stack_13_io_ray_id),
    .io_dataOut(Stack_13_io_dataOut),
    .io_empty(Stack_13_io_empty),
    .io_hit_in(Stack_13_io_hit_in),
    .io_hit_out(Stack_13_io_hit_out),
    .io_ray_out(Stack_13_io_ray_out),
    .io_enable(Stack_13_io_enable)
  );
  Stack Stack_14 ( // @[stackmanage_35.scala 50:47]
    .clock(Stack_14_clock),
    .reset(Stack_14_reset),
    .io_push(Stack_14_io_push),
    .io_pop(Stack_14_io_pop),
    .io_dataIn(Stack_14_io_dataIn),
    .io_clear(Stack_14_io_clear),
    .io_ray_id(Stack_14_io_ray_id),
    .io_dataOut(Stack_14_io_dataOut),
    .io_empty(Stack_14_io_empty),
    .io_hit_in(Stack_14_io_hit_in),
    .io_hit_out(Stack_14_io_hit_out),
    .io_ray_out(Stack_14_io_ray_out),
    .io_enable(Stack_14_io_enable)
  );
  Stack Stack_15 ( // @[stackmanage_35.scala 51:47]
    .clock(Stack_15_clock),
    .reset(Stack_15_reset),
    .io_push(Stack_15_io_push),
    .io_pop(Stack_15_io_pop),
    .io_dataIn(Stack_15_io_dataIn),
    .io_clear(Stack_15_io_clear),
    .io_ray_id(Stack_15_io_ray_id),
    .io_dataOut(Stack_15_io_dataOut),
    .io_empty(Stack_15_io_empty),
    .io_hit_in(Stack_15_io_hit_in),
    .io_hit_out(Stack_15_io_hit_out),
    .io_ray_out(Stack_15_io_ray_out),
    .io_enable(Stack_15_io_enable)
  );
  Stack Stack_16 ( // @[stackmanage_35.scala 52:49]
    .clock(Stack_16_clock),
    .reset(Stack_16_reset),
    .io_push(Stack_16_io_push),
    .io_pop(Stack_16_io_pop),
    .io_dataIn(Stack_16_io_dataIn),
    .io_clear(Stack_16_io_clear),
    .io_ray_id(Stack_16_io_ray_id),
    .io_dataOut(Stack_16_io_dataOut),
    .io_empty(Stack_16_io_empty),
    .io_hit_in(Stack_16_io_hit_in),
    .io_hit_out(Stack_16_io_hit_out),
    .io_ray_out(Stack_16_io_ray_out),
    .io_enable(Stack_16_io_enable)
  );
  Stack Stack_17 ( // @[stackmanage_35.scala 53:49]
    .clock(Stack_17_clock),
    .reset(Stack_17_reset),
    .io_push(Stack_17_io_push),
    .io_pop(Stack_17_io_pop),
    .io_dataIn(Stack_17_io_dataIn),
    .io_clear(Stack_17_io_clear),
    .io_ray_id(Stack_17_io_ray_id),
    .io_dataOut(Stack_17_io_dataOut),
    .io_empty(Stack_17_io_empty),
    .io_hit_in(Stack_17_io_hit_in),
    .io_hit_out(Stack_17_io_hit_out),
    .io_ray_out(Stack_17_io_ray_out),
    .io_enable(Stack_17_io_enable)
  );
  Stack Stack_18 ( // @[stackmanage_35.scala 54:49]
    .clock(Stack_18_clock),
    .reset(Stack_18_reset),
    .io_push(Stack_18_io_push),
    .io_pop(Stack_18_io_pop),
    .io_dataIn(Stack_18_io_dataIn),
    .io_clear(Stack_18_io_clear),
    .io_ray_id(Stack_18_io_ray_id),
    .io_dataOut(Stack_18_io_dataOut),
    .io_empty(Stack_18_io_empty),
    .io_hit_in(Stack_18_io_hit_in),
    .io_hit_out(Stack_18_io_hit_out),
    .io_ray_out(Stack_18_io_ray_out),
    .io_enable(Stack_18_io_enable)
  );
  Stack Stack_19 ( // @[stackmanage_35.scala 55:49]
    .clock(Stack_19_clock),
    .reset(Stack_19_reset),
    .io_push(Stack_19_io_push),
    .io_pop(Stack_19_io_pop),
    .io_dataIn(Stack_19_io_dataIn),
    .io_clear(Stack_19_io_clear),
    .io_ray_id(Stack_19_io_ray_id),
    .io_dataOut(Stack_19_io_dataOut),
    .io_empty(Stack_19_io_empty),
    .io_hit_in(Stack_19_io_hit_in),
    .io_hit_out(Stack_19_io_hit_out),
    .io_ray_out(Stack_19_io_ray_out),
    .io_enable(Stack_19_io_enable)
  );
  Stack Stack_20 ( // @[stackmanage_35.scala 56:49]
    .clock(Stack_20_clock),
    .reset(Stack_20_reset),
    .io_push(Stack_20_io_push),
    .io_pop(Stack_20_io_pop),
    .io_dataIn(Stack_20_io_dataIn),
    .io_clear(Stack_20_io_clear),
    .io_ray_id(Stack_20_io_ray_id),
    .io_dataOut(Stack_20_io_dataOut),
    .io_empty(Stack_20_io_empty),
    .io_hit_in(Stack_20_io_hit_in),
    .io_hit_out(Stack_20_io_hit_out),
    .io_ray_out(Stack_20_io_ray_out),
    .io_enable(Stack_20_io_enable)
  );
  Stack Stack_21 ( // @[stackmanage_35.scala 57:49]
    .clock(Stack_21_clock),
    .reset(Stack_21_reset),
    .io_push(Stack_21_io_push),
    .io_pop(Stack_21_io_pop),
    .io_dataIn(Stack_21_io_dataIn),
    .io_clear(Stack_21_io_clear),
    .io_ray_id(Stack_21_io_ray_id),
    .io_dataOut(Stack_21_io_dataOut),
    .io_empty(Stack_21_io_empty),
    .io_hit_in(Stack_21_io_hit_in),
    .io_hit_out(Stack_21_io_hit_out),
    .io_ray_out(Stack_21_io_ray_out),
    .io_enable(Stack_21_io_enable)
  );
  Stack Stack_22 ( // @[stackmanage_35.scala 58:49]
    .clock(Stack_22_clock),
    .reset(Stack_22_reset),
    .io_push(Stack_22_io_push),
    .io_pop(Stack_22_io_pop),
    .io_dataIn(Stack_22_io_dataIn),
    .io_clear(Stack_22_io_clear),
    .io_ray_id(Stack_22_io_ray_id),
    .io_dataOut(Stack_22_io_dataOut),
    .io_empty(Stack_22_io_empty),
    .io_hit_in(Stack_22_io_hit_in),
    .io_hit_out(Stack_22_io_hit_out),
    .io_ray_out(Stack_22_io_ray_out),
    .io_enable(Stack_22_io_enable)
  );
  Stack Stack_23 ( // @[stackmanage_35.scala 59:48]
    .clock(Stack_23_clock),
    .reset(Stack_23_reset),
    .io_push(Stack_23_io_push),
    .io_pop(Stack_23_io_pop),
    .io_dataIn(Stack_23_io_dataIn),
    .io_clear(Stack_23_io_clear),
    .io_ray_id(Stack_23_io_ray_id),
    .io_dataOut(Stack_23_io_dataOut),
    .io_empty(Stack_23_io_empty),
    .io_hit_in(Stack_23_io_hit_in),
    .io_hit_out(Stack_23_io_hit_out),
    .io_ray_out(Stack_23_io_ray_out),
    .io_enable(Stack_23_io_enable)
  );
  Stack Stack_24 ( // @[stackmanage_35.scala 60:48]
    .clock(Stack_24_clock),
    .reset(Stack_24_reset),
    .io_push(Stack_24_io_push),
    .io_pop(Stack_24_io_pop),
    .io_dataIn(Stack_24_io_dataIn),
    .io_clear(Stack_24_io_clear),
    .io_ray_id(Stack_24_io_ray_id),
    .io_dataOut(Stack_24_io_dataOut),
    .io_empty(Stack_24_io_empty),
    .io_hit_in(Stack_24_io_hit_in),
    .io_hit_out(Stack_24_io_hit_out),
    .io_ray_out(Stack_24_io_ray_out),
    .io_enable(Stack_24_io_enable)
  );
  Stack Stack_25 ( // @[stackmanage_35.scala 61:49]
    .clock(Stack_25_clock),
    .reset(Stack_25_reset),
    .io_push(Stack_25_io_push),
    .io_pop(Stack_25_io_pop),
    .io_dataIn(Stack_25_io_dataIn),
    .io_clear(Stack_25_io_clear),
    .io_ray_id(Stack_25_io_ray_id),
    .io_dataOut(Stack_25_io_dataOut),
    .io_empty(Stack_25_io_empty),
    .io_hit_in(Stack_25_io_hit_in),
    .io_hit_out(Stack_25_io_hit_out),
    .io_ray_out(Stack_25_io_ray_out),
    .io_enable(Stack_25_io_enable)
  );
  Stack Stack_26 ( // @[stackmanage_35.scala 62:47]
    .clock(Stack_26_clock),
    .reset(Stack_26_reset),
    .io_push(Stack_26_io_push),
    .io_pop(Stack_26_io_pop),
    .io_dataIn(Stack_26_io_dataIn),
    .io_clear(Stack_26_io_clear),
    .io_ray_id(Stack_26_io_ray_id),
    .io_dataOut(Stack_26_io_dataOut),
    .io_empty(Stack_26_io_empty),
    .io_hit_in(Stack_26_io_hit_in),
    .io_hit_out(Stack_26_io_hit_out),
    .io_ray_out(Stack_26_io_ray_out),
    .io_enable(Stack_26_io_enable)
  );
  Stack Stack_27 ( // @[stackmanage_35.scala 63:47]
    .clock(Stack_27_clock),
    .reset(Stack_27_reset),
    .io_push(Stack_27_io_push),
    .io_pop(Stack_27_io_pop),
    .io_dataIn(Stack_27_io_dataIn),
    .io_clear(Stack_27_io_clear),
    .io_ray_id(Stack_27_io_ray_id),
    .io_dataOut(Stack_27_io_dataOut),
    .io_empty(Stack_27_io_empty),
    .io_hit_in(Stack_27_io_hit_in),
    .io_hit_out(Stack_27_io_hit_out),
    .io_ray_out(Stack_27_io_ray_out),
    .io_enable(Stack_27_io_enable)
  );
  Stack Stack_28 ( // @[stackmanage_35.scala 64:47]
    .clock(Stack_28_clock),
    .reset(Stack_28_reset),
    .io_push(Stack_28_io_push),
    .io_pop(Stack_28_io_pop),
    .io_dataIn(Stack_28_io_dataIn),
    .io_clear(Stack_28_io_clear),
    .io_ray_id(Stack_28_io_ray_id),
    .io_dataOut(Stack_28_io_dataOut),
    .io_empty(Stack_28_io_empty),
    .io_hit_in(Stack_28_io_hit_in),
    .io_hit_out(Stack_28_io_hit_out),
    .io_ray_out(Stack_28_io_ray_out),
    .io_enable(Stack_28_io_enable)
  );
  Stack Stack_29 ( // @[stackmanage_35.scala 65:47]
    .clock(Stack_29_clock),
    .reset(Stack_29_reset),
    .io_push(Stack_29_io_push),
    .io_pop(Stack_29_io_pop),
    .io_dataIn(Stack_29_io_dataIn),
    .io_clear(Stack_29_io_clear),
    .io_ray_id(Stack_29_io_ray_id),
    .io_dataOut(Stack_29_io_dataOut),
    .io_empty(Stack_29_io_empty),
    .io_hit_in(Stack_29_io_hit_in),
    .io_hit_out(Stack_29_io_hit_out),
    .io_ray_out(Stack_29_io_ray_out),
    .io_enable(Stack_29_io_enable)
  );
  Stack Stack_30 ( // @[stackmanage_35.scala 66:47]
    .clock(Stack_30_clock),
    .reset(Stack_30_reset),
    .io_push(Stack_30_io_push),
    .io_pop(Stack_30_io_pop),
    .io_dataIn(Stack_30_io_dataIn),
    .io_clear(Stack_30_io_clear),
    .io_ray_id(Stack_30_io_ray_id),
    .io_dataOut(Stack_30_io_dataOut),
    .io_empty(Stack_30_io_empty),
    .io_hit_in(Stack_30_io_hit_in),
    .io_hit_out(Stack_30_io_hit_out),
    .io_ray_out(Stack_30_io_ray_out),
    .io_enable(Stack_30_io_enable)
  );
  Stack Stack_31 ( // @[stackmanage_35.scala 67:47]
    .clock(Stack_31_clock),
    .reset(Stack_31_reset),
    .io_push(Stack_31_io_push),
    .io_pop(Stack_31_io_pop),
    .io_dataIn(Stack_31_io_dataIn),
    .io_clear(Stack_31_io_clear),
    .io_ray_id(Stack_31_io_ray_id),
    .io_dataOut(Stack_31_io_dataOut),
    .io_empty(Stack_31_io_empty),
    .io_hit_in(Stack_31_io_hit_in),
    .io_hit_out(Stack_31_io_hit_out),
    .io_ray_out(Stack_31_io_ray_out),
    .io_enable(Stack_31_io_enable)
  );
  Stack Stack_32 ( // @[stackmanage_35.scala 68:49]
    .clock(Stack_32_clock),
    .reset(Stack_32_reset),
    .io_push(Stack_32_io_push),
    .io_pop(Stack_32_io_pop),
    .io_dataIn(Stack_32_io_dataIn),
    .io_clear(Stack_32_io_clear),
    .io_ray_id(Stack_32_io_ray_id),
    .io_dataOut(Stack_32_io_dataOut),
    .io_empty(Stack_32_io_empty),
    .io_hit_in(Stack_32_io_hit_in),
    .io_hit_out(Stack_32_io_hit_out),
    .io_ray_out(Stack_32_io_ray_out),
    .io_enable(Stack_32_io_enable)
  );
  Stack Stack_33 ( // @[stackmanage_35.scala 69:48]
    .clock(Stack_33_clock),
    .reset(Stack_33_reset),
    .io_push(Stack_33_io_push),
    .io_pop(Stack_33_io_pop),
    .io_dataIn(Stack_33_io_dataIn),
    .io_clear(Stack_33_io_clear),
    .io_ray_id(Stack_33_io_ray_id),
    .io_dataOut(Stack_33_io_dataOut),
    .io_empty(Stack_33_io_empty),
    .io_hit_in(Stack_33_io_hit_in),
    .io_hit_out(Stack_33_io_hit_out),
    .io_ray_out(Stack_33_io_ray_out),
    .io_enable(Stack_33_io_enable)
  );
  Stack Stack_34 ( // @[stackmanage_35.scala 70:48]
    .clock(Stack_34_clock),
    .reset(Stack_34_reset),
    .io_push(Stack_34_io_push),
    .io_pop(Stack_34_io_pop),
    .io_dataIn(Stack_34_io_dataIn),
    .io_clear(Stack_34_io_clear),
    .io_ray_id(Stack_34_io_ray_id),
    .io_dataOut(Stack_34_io_dataOut),
    .io_empty(Stack_34_io_empty),
    .io_hit_in(Stack_34_io_hit_in),
    .io_hit_out(Stack_34_io_hit_out),
    .io_ray_out(Stack_34_io_ray_out),
    .io_enable(Stack_34_io_enable)
  );
  assign io_hitT_out = hitT_out_temp; // @[stackmanage_35.scala 4515:33]
  assign io_node_id_out = node_out_temp; // @[stackmanage_35.scala 4516:27]
  assign io_ray_id_out = ray_out_temp; // @[stackmanage_35.scala 4517:30]
  assign io_pop_valid = pop_valid_1; // @[stackmanage_35.scala 4518:31]
  assign io_Dis_en = _T_468 | dispatch_25 | dispatch_26 | dispatch_27 | dispatch_28 | dispatch_29 | dispatch_30 |
    dispatch_31 | dispatch_32 | dispatch_33 | dispatch_34 | dispatch_no_match; // @[stackmanage_35.scala 5989:275]
  assign io_Finish = _T_514 & Stack_25_io_empty & Stack_26_io_empty & Stack_27_io_empty & Stack_28_io_empty &
    Stack_29_io_empty & Stack_30_io_empty & Stack_31_io_empty & Stack_32_io_empty & Stack_33_io_empty &
    Stack_34_io_empty; // @[stackmanage_35.scala 5991:237]
  assign LUT_stack_clock = clock;
  assign LUT_stack_reset = reset;
  assign LUT_stack_io_push = io_push; // @[stackmanage_35.scala 234:38]
  assign LUT_stack_io_push_valid = io_push_en; // @[stackmanage_35.scala 235:38]
  assign LUT_stack_io_pop = io_pop; // @[stackmanage_35.scala 236:38]
  assign LUT_stack_io_pop_valid = io_pop_en; // @[stackmanage_35.scala 237:38]
  assign LUT_stack_io_clear = io_clear; // @[stackmanage_35.scala 243:38]
  assign LUT_stack_io_empty_0 = Stack_0_io_empty; // @[stackmanage_35.scala 72:29]
  assign LUT_stack_io_empty_1 = Stack_1_io_empty; // @[stackmanage_35.scala 73:29]
  assign LUT_stack_io_empty_2 = Stack_2_io_empty; // @[stackmanage_35.scala 74:29]
  assign LUT_stack_io_empty_3 = Stack_3_io_empty; // @[stackmanage_35.scala 75:29]
  assign LUT_stack_io_empty_4 = Stack_4_io_empty; // @[stackmanage_35.scala 76:29]
  assign LUT_stack_io_empty_5 = Stack_5_io_empty; // @[stackmanage_35.scala 77:29]
  assign LUT_stack_io_empty_6 = Stack_6_io_empty; // @[stackmanage_35.scala 78:29]
  assign LUT_stack_io_empty_7 = Stack_7_io_empty; // @[stackmanage_35.scala 79:29]
  assign LUT_stack_io_empty_8 = Stack_8_io_empty; // @[stackmanage_35.scala 80:29]
  assign LUT_stack_io_empty_9 = Stack_9_io_empty; // @[stackmanage_35.scala 81:29]
  assign LUT_stack_io_empty_10 = Stack_10_io_empty; // @[stackmanage_35.scala 83:30]
  assign LUT_stack_io_empty_11 = Stack_11_io_empty; // @[stackmanage_35.scala 84:30]
  assign LUT_stack_io_empty_12 = Stack_12_io_empty; // @[stackmanage_35.scala 85:30]
  assign LUT_stack_io_empty_13 = Stack_13_io_empty; // @[stackmanage_35.scala 86:30]
  assign LUT_stack_io_empty_14 = Stack_14_io_empty; // @[stackmanage_35.scala 87:30]
  assign LUT_stack_io_empty_15 = Stack_15_io_empty; // @[stackmanage_35.scala 88:30]
  assign LUT_stack_io_empty_16 = Stack_16_io_empty; // @[stackmanage_35.scala 89:30]
  assign LUT_stack_io_empty_17 = Stack_17_io_empty; // @[stackmanage_35.scala 90:30]
  assign LUT_stack_io_empty_18 = Stack_18_io_empty; // @[stackmanage_35.scala 91:30]
  assign LUT_stack_io_empty_19 = Stack_19_io_empty; // @[stackmanage_35.scala 92:30]
  assign LUT_stack_io_empty_20 = Stack_20_io_empty; // @[stackmanage_35.scala 94:30]
  assign LUT_stack_io_empty_21 = Stack_21_io_empty; // @[stackmanage_35.scala 95:30]
  assign LUT_stack_io_empty_22 = Stack_22_io_empty; // @[stackmanage_35.scala 96:30]
  assign LUT_stack_io_empty_23 = Stack_23_io_empty; // @[stackmanage_35.scala 97:30]
  assign LUT_stack_io_empty_24 = Stack_24_io_empty; // @[stackmanage_35.scala 98:30]
  assign LUT_stack_io_empty_25 = Stack_25_io_empty; // @[stackmanage_35.scala 99:30]
  assign LUT_stack_io_empty_26 = Stack_26_io_empty; // @[stackmanage_35.scala 100:30]
  assign LUT_stack_io_empty_27 = Stack_27_io_empty; // @[stackmanage_35.scala 101:30]
  assign LUT_stack_io_empty_28 = Stack_28_io_empty; // @[stackmanage_35.scala 102:30]
  assign LUT_stack_io_empty_29 = Stack_29_io_empty; // @[stackmanage_35.scala 103:30]
  assign LUT_stack_io_empty_30 = Stack_30_io_empty; // @[stackmanage_35.scala 105:30]
  assign LUT_stack_io_empty_31 = Stack_31_io_empty; // @[stackmanage_35.scala 106:30]
  assign LUT_stack_io_empty_32 = Stack_32_io_empty; // @[stackmanage_35.scala 107:30]
  assign LUT_stack_io_empty_33 = Stack_33_io_empty; // @[stackmanage_35.scala 108:30]
  assign LUT_stack_io_empty_34 = Stack_34_io_empty; // @[stackmanage_35.scala 109:30]
  assign LUT_stack_io_dispatch_0 = dispatch_0; // @[stackmanage_35.scala 5995:39]
  assign LUT_stack_io_dispatch_1 = dispatch_1; // @[stackmanage_35.scala 5996:39]
  assign LUT_stack_io_dispatch_2 = dispatch_2; // @[stackmanage_35.scala 5997:39]
  assign LUT_stack_io_dispatch_3 = dispatch_3; // @[stackmanage_35.scala 5998:39]
  assign LUT_stack_io_dispatch_4 = dispatch_4; // @[stackmanage_35.scala 5999:39]
  assign LUT_stack_io_dispatch_5 = dispatch_5; // @[stackmanage_35.scala 6000:39]
  assign LUT_stack_io_dispatch_6 = dispatch_6; // @[stackmanage_35.scala 6001:39]
  assign LUT_stack_io_dispatch_7 = dispatch_7; // @[stackmanage_35.scala 6002:39]
  assign LUT_stack_io_dispatch_8 = dispatch_8; // @[stackmanage_35.scala 6003:39]
  assign LUT_stack_io_dispatch_9 = dispatch_9; // @[stackmanage_35.scala 6004:39]
  assign LUT_stack_io_dispatch_10 = dispatch_10; // @[stackmanage_35.scala 6005:40]
  assign LUT_stack_io_dispatch_11 = dispatch_11; // @[stackmanage_35.scala 6006:40]
  assign LUT_stack_io_dispatch_12 = dispatch_12; // @[stackmanage_35.scala 6007:40]
  assign LUT_stack_io_dispatch_13 = dispatch_13; // @[stackmanage_35.scala 6008:40]
  assign LUT_stack_io_dispatch_14 = dispatch_14; // @[stackmanage_35.scala 6009:40]
  assign LUT_stack_io_dispatch_15 = dispatch_15; // @[stackmanage_35.scala 6010:40]
  assign LUT_stack_io_dispatch_16 = dispatch_16; // @[stackmanage_35.scala 6011:40]
  assign LUT_stack_io_dispatch_17 = dispatch_17; // @[stackmanage_35.scala 6012:40]
  assign LUT_stack_io_dispatch_18 = dispatch_18; // @[stackmanage_35.scala 6013:40]
  assign LUT_stack_io_dispatch_19 = dispatch_19; // @[stackmanage_35.scala 6014:40]
  assign LUT_stack_io_dispatch_20 = dispatch_20; // @[stackmanage_35.scala 6015:40]
  assign LUT_stack_io_dispatch_21 = dispatch_21; // @[stackmanage_35.scala 6016:40]
  assign LUT_stack_io_dispatch_22 = dispatch_22; // @[stackmanage_35.scala 6017:40]
  assign LUT_stack_io_dispatch_23 = dispatch_23; // @[stackmanage_35.scala 6018:40]
  assign LUT_stack_io_dispatch_24 = dispatch_24; // @[stackmanage_35.scala 6019:40]
  assign LUT_stack_io_dispatch_25 = dispatch_25; // @[stackmanage_35.scala 6020:40]
  assign LUT_stack_io_dispatch_26 = dispatch_26; // @[stackmanage_35.scala 6021:40]
  assign LUT_stack_io_dispatch_27 = dispatch_27; // @[stackmanage_35.scala 6022:40]
  assign LUT_stack_io_dispatch_28 = dispatch_28; // @[stackmanage_35.scala 6023:40]
  assign LUT_stack_io_dispatch_29 = dispatch_29; // @[stackmanage_35.scala 6024:40]
  assign LUT_stack_io_dispatch_30 = dispatch_30; // @[stackmanage_35.scala 6025:40]
  assign LUT_stack_io_dispatch_31 = dispatch_31; // @[stackmanage_35.scala 6026:40]
  assign LUT_stack_io_dispatch_32 = dispatch_32; // @[stackmanage_35.scala 6027:40]
  assign LUT_stack_io_dispatch_33 = dispatch_33; // @[stackmanage_35.scala 6028:40]
  assign LUT_stack_io_dispatch_34 = dispatch_34; // @[stackmanage_35.scala 6029:40]
  assign LUT_stack_io_ray_id_push = io_ray_id_push; // @[stackmanage_35.scala 238:38]
  assign LUT_stack_io_ray_id_pop = io_ray_id_pop; // @[stackmanage_35.scala 239:38]
  assign LUT_stack_io_node_id_push_in = io_node_id_push_in; // @[stackmanage_35.scala 240:38]
  assign LUT_stack_io_hitT_in = io_hitT_in; // @[stackmanage_35.scala 242:38]
  assign Stack_0_clock = clock;
  assign Stack_0_reset = reset;
  assign Stack_0_io_push = LUT_stack_io_push_0; // @[stackmanage_35.scala 151:37]
  assign Stack_0_io_pop = LUT_stack_io_pop_0; // @[stackmanage_35.scala 112:38]
  assign Stack_0_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 383:64 stackmanage_35.scala 384:28]
  assign Stack_0_io_clear = LUT_stack_io_clear_0; // @[stackmanage_35.scala 192:38]
  assign Stack_0_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1688:28]
  assign Stack_0_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1687:28]
  assign Stack_1_clock = clock;
  assign Stack_1_reset = reset;
  assign Stack_1_io_push = LUT_stack_io_push_1; // @[stackmanage_35.scala 152:37]
  assign Stack_1_io_pop = LUT_stack_io_pop_1; // @[stackmanage_35.scala 113:38]
  assign Stack_1_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_594); // @[stackmanage_35.scala 383:64 stackmanage_35.scala 385:30]
  assign Stack_1_io_clear = LUT_stack_io_clear_1; // @[stackmanage_35.scala 193:38]
  assign Stack_1_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1820; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1690:27]
  assign Stack_1_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1819; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1689:28]
  assign Stack_2_clock = clock;
  assign Stack_2_reset = reset;
  assign Stack_2_io_push = LUT_stack_io_push_2; // @[stackmanage_35.scala 153:37]
  assign Stack_2_io_pop = LUT_stack_io_pop_2; // @[stackmanage_35.scala 114:38]
  assign Stack_2_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_596); // @[stackmanage_35.scala 383:64 stackmanage_35.scala 386:30]
  assign Stack_2_io_clear = LUT_stack_io_clear_2; // @[stackmanage_35.scala 194:38]
  assign Stack_2_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1823; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1692:27]
  assign Stack_2_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1822; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1691:28]
  assign Stack_3_clock = clock;
  assign Stack_3_reset = reset;
  assign Stack_3_io_push = LUT_stack_io_push_3; // @[stackmanage_35.scala 154:37]
  assign Stack_3_io_pop = LUT_stack_io_pop_3; // @[stackmanage_35.scala 115:38]
  assign Stack_3_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_597); // @[stackmanage_35.scala 383:64 stackmanage_35.scala 387:30]
  assign Stack_3_io_clear = LUT_stack_io_clear_3; // @[stackmanage_35.scala 195:38]
  assign Stack_3_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1825; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1694:27]
  assign Stack_3_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1824; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1693:28]
  assign Stack_4_clock = clock;
  assign Stack_4_reset = reset;
  assign Stack_4_io_push = LUT_stack_io_push_4; // @[stackmanage_35.scala 155:37]
  assign Stack_4_io_pop = LUT_stack_io_pop_4; // @[stackmanage_35.scala 116:38]
  assign Stack_4_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_598); // @[stackmanage_35.scala 383:64 stackmanage_35.scala 388:30]
  assign Stack_4_io_clear = LUT_stack_io_clear_4; // @[stackmanage_35.scala 196:38]
  assign Stack_4_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1827; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1696:27]
  assign Stack_4_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1826; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1695:28]
  assign Stack_5_clock = clock;
  assign Stack_5_reset = reset;
  assign Stack_5_io_push = LUT_stack_io_push_5; // @[stackmanage_35.scala 156:37]
  assign Stack_5_io_pop = LUT_stack_io_pop_5; // @[stackmanage_35.scala 117:38]
  assign Stack_5_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_599); // @[stackmanage_35.scala 383:64 stackmanage_35.scala 389:30]
  assign Stack_5_io_clear = LUT_stack_io_clear_5; // @[stackmanage_35.scala 197:38]
  assign Stack_5_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1829; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1698:27]
  assign Stack_5_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1828; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1697:28]
  assign Stack_6_clock = clock;
  assign Stack_6_reset = reset;
  assign Stack_6_io_push = LUT_stack_io_push_6; // @[stackmanage_35.scala 157:37]
  assign Stack_6_io_pop = LUT_stack_io_pop_6; // @[stackmanage_35.scala 118:38]
  assign Stack_6_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_600); // @[stackmanage_35.scala 383:64 stackmanage_35.scala 390:30]
  assign Stack_6_io_clear = LUT_stack_io_clear_6; // @[stackmanage_35.scala 198:38]
  assign Stack_6_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1831; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1700:27]
  assign Stack_6_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1830; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1699:28]
  assign Stack_7_clock = clock;
  assign Stack_7_reset = reset;
  assign Stack_7_io_push = LUT_stack_io_push_7; // @[stackmanage_35.scala 158:37]
  assign Stack_7_io_pop = LUT_stack_io_pop_7; // @[stackmanage_35.scala 119:38]
  assign Stack_7_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_601); // @[stackmanage_35.scala 383:64 stackmanage_35.scala 391:30]
  assign Stack_7_io_clear = LUT_stack_io_clear_7; // @[stackmanage_35.scala 199:38]
  assign Stack_7_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1833; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1702:27]
  assign Stack_7_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1832; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1701:28]
  assign Stack_8_clock = clock;
  assign Stack_8_reset = reset;
  assign Stack_8_io_push = LUT_stack_io_push_8; // @[stackmanage_35.scala 159:37]
  assign Stack_8_io_pop = LUT_stack_io_pop_8; // @[stackmanage_35.scala 120:38]
  assign Stack_8_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_602); // @[stackmanage_35.scala 383:64 stackmanage_35.scala 392:30]
  assign Stack_8_io_clear = LUT_stack_io_clear_8; // @[stackmanage_35.scala 200:38]
  assign Stack_8_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1835; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1704:27]
  assign Stack_8_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1834; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1703:28]
  assign Stack_9_clock = clock;
  assign Stack_9_reset = reset;
  assign Stack_9_io_push = LUT_stack_io_push_9; // @[stackmanage_35.scala 160:37]
  assign Stack_9_io_pop = LUT_stack_io_pop_9; // @[stackmanage_35.scala 121:38]
  assign Stack_9_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_603); // @[stackmanage_35.scala 383:64 stackmanage_35.scala 393:30]
  assign Stack_9_io_clear = LUT_stack_io_clear_9; // @[stackmanage_35.scala 201:38]
  assign Stack_9_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1837; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1706:27]
  assign Stack_9_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1836; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1705:28]
  assign Stack_10_clock = clock;
  assign Stack_10_reset = reset;
  assign Stack_10_io_push = LUT_stack_io_push_10; // @[stackmanage_35.scala 162:38]
  assign Stack_10_io_pop = LUT_stack_io_pop_10; // @[stackmanage_35.scala 123:39]
  assign Stack_10_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_604); // @[stackmanage_35.scala 383:64 stackmanage_35.scala 394:31]
  assign Stack_10_io_clear = LUT_stack_io_clear_10; // @[stackmanage_35.scala 203:39]
  assign Stack_10_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1839; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1708:29]
  assign Stack_10_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1838; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1707:29]
  assign Stack_11_clock = clock;
  assign Stack_11_reset = reset;
  assign Stack_11_io_push = LUT_stack_io_push_11; // @[stackmanage_35.scala 163:38]
  assign Stack_11_io_pop = LUT_stack_io_pop_11; // @[stackmanage_35.scala 124:39]
  assign Stack_11_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_605); // @[stackmanage_35.scala 383:64 stackmanage_35.scala 395:31]
  assign Stack_11_io_clear = LUT_stack_io_clear_11; // @[stackmanage_35.scala 204:39]
  assign Stack_11_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1841; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1710:28]
  assign Stack_11_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1840; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1709:29]
  assign Stack_12_clock = clock;
  assign Stack_12_reset = reset;
  assign Stack_12_io_push = LUT_stack_io_push_12; // @[stackmanage_35.scala 164:38]
  assign Stack_12_io_pop = LUT_stack_io_pop_12; // @[stackmanage_35.scala 125:39]
  assign Stack_12_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_606); // @[stackmanage_35.scala 383:64 stackmanage_35.scala 396:31]
  assign Stack_12_io_clear = LUT_stack_io_clear_12; // @[stackmanage_35.scala 205:39]
  assign Stack_12_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1843; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1712:28]
  assign Stack_12_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1842; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1711:29]
  assign Stack_13_clock = clock;
  assign Stack_13_reset = reset;
  assign Stack_13_io_push = LUT_stack_io_push_13; // @[stackmanage_35.scala 165:38]
  assign Stack_13_io_pop = LUT_stack_io_pop_13; // @[stackmanage_35.scala 126:39]
  assign Stack_13_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_607); // @[stackmanage_35.scala 383:64 stackmanage_35.scala 397:31]
  assign Stack_13_io_clear = LUT_stack_io_clear_13; // @[stackmanage_35.scala 206:39]
  assign Stack_13_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1845; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1714:28]
  assign Stack_13_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1844; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1713:29]
  assign Stack_14_clock = clock;
  assign Stack_14_reset = reset;
  assign Stack_14_io_push = LUT_stack_io_push_14; // @[stackmanage_35.scala 166:38]
  assign Stack_14_io_pop = LUT_stack_io_pop_14; // @[stackmanage_35.scala 127:39]
  assign Stack_14_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_608); // @[stackmanage_35.scala 383:64 stackmanage_35.scala 398:31]
  assign Stack_14_io_clear = LUT_stack_io_clear_14; // @[stackmanage_35.scala 207:39]
  assign Stack_14_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1847; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1716:28]
  assign Stack_14_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1846; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1715:29]
  assign Stack_15_clock = clock;
  assign Stack_15_reset = reset;
  assign Stack_15_io_push = LUT_stack_io_push_15; // @[stackmanage_35.scala 167:38]
  assign Stack_15_io_pop = LUT_stack_io_pop_15; // @[stackmanage_35.scala 128:39]
  assign Stack_15_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_609); // @[stackmanage_35.scala 383:64 stackmanage_35.scala 399:31]
  assign Stack_15_io_clear = LUT_stack_io_clear_15; // @[stackmanage_35.scala 208:39]
  assign Stack_15_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1849; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1718:28]
  assign Stack_15_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1848; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1717:29]
  assign Stack_16_clock = clock;
  assign Stack_16_reset = reset;
  assign Stack_16_io_push = LUT_stack_io_push_16; // @[stackmanage_35.scala 168:38]
  assign Stack_16_io_pop = LUT_stack_io_pop_16; // @[stackmanage_35.scala 129:39]
  assign Stack_16_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_610); // @[stackmanage_35.scala 383:64 stackmanage_35.scala 400:31]
  assign Stack_16_io_clear = LUT_stack_io_clear_16; // @[stackmanage_35.scala 209:39]
  assign Stack_16_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1851; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1720:28]
  assign Stack_16_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1850; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1719:29]
  assign Stack_17_clock = clock;
  assign Stack_17_reset = reset;
  assign Stack_17_io_push = LUT_stack_io_push_17; // @[stackmanage_35.scala 169:38]
  assign Stack_17_io_pop = LUT_stack_io_pop_17; // @[stackmanage_35.scala 130:39]
  assign Stack_17_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_611); // @[stackmanage_35.scala 383:64 stackmanage_35.scala 401:31]
  assign Stack_17_io_clear = LUT_stack_io_clear_17; // @[stackmanage_35.scala 210:39]
  assign Stack_17_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1853; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1722:28]
  assign Stack_17_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1852; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1721:29]
  assign Stack_18_clock = clock;
  assign Stack_18_reset = reset;
  assign Stack_18_io_push = LUT_stack_io_push_18; // @[stackmanage_35.scala 170:38]
  assign Stack_18_io_pop = LUT_stack_io_pop_18; // @[stackmanage_35.scala 131:39]
  assign Stack_18_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_612); // @[stackmanage_35.scala 383:64 stackmanage_35.scala 402:31]
  assign Stack_18_io_clear = LUT_stack_io_clear_18; // @[stackmanage_35.scala 211:39]
  assign Stack_18_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1855; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1724:28]
  assign Stack_18_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1854; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1723:29]
  assign Stack_19_clock = clock;
  assign Stack_19_reset = reset;
  assign Stack_19_io_push = LUT_stack_io_push_19; // @[stackmanage_35.scala 171:38]
  assign Stack_19_io_pop = LUT_stack_io_pop_19; // @[stackmanage_35.scala 132:39]
  assign Stack_19_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_613); // @[stackmanage_35.scala 383:64 stackmanage_35.scala 403:31]
  assign Stack_19_io_clear = LUT_stack_io_clear_19; // @[stackmanage_35.scala 212:39]
  assign Stack_19_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1857; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1726:28]
  assign Stack_19_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1856; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1725:29]
  assign Stack_20_clock = clock;
  assign Stack_20_reset = reset;
  assign Stack_20_io_push = LUT_stack_io_push_20; // @[stackmanage_35.scala 173:38]
  assign Stack_20_io_pop = LUT_stack_io_pop_20; // @[stackmanage_35.scala 134:39]
  assign Stack_20_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_614); // @[stackmanage_35.scala 383:64 stackmanage_35.scala 404:31]
  assign Stack_20_io_clear = LUT_stack_io_clear_20; // @[stackmanage_35.scala 214:39]
  assign Stack_20_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1859; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1728:29]
  assign Stack_20_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1858; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1727:29]
  assign Stack_21_clock = clock;
  assign Stack_21_reset = reset;
  assign Stack_21_io_push = LUT_stack_io_push_21; // @[stackmanage_35.scala 174:38]
  assign Stack_21_io_pop = LUT_stack_io_pop_21; // @[stackmanage_35.scala 135:39]
  assign Stack_21_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_615); // @[stackmanage_35.scala 383:64 stackmanage_35.scala 405:31]
  assign Stack_21_io_clear = LUT_stack_io_clear_21; // @[stackmanage_35.scala 215:39]
  assign Stack_21_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1861; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1730:28]
  assign Stack_21_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1860; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1729:29]
  assign Stack_22_clock = clock;
  assign Stack_22_reset = reset;
  assign Stack_22_io_push = LUT_stack_io_push_22; // @[stackmanage_35.scala 175:38]
  assign Stack_22_io_pop = LUT_stack_io_pop_22; // @[stackmanage_35.scala 136:39]
  assign Stack_22_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_616); // @[stackmanage_35.scala 383:64 stackmanage_35.scala 406:31]
  assign Stack_22_io_clear = LUT_stack_io_clear_22; // @[stackmanage_35.scala 216:39]
  assign Stack_22_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1863; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1732:28]
  assign Stack_22_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1862; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1731:29]
  assign Stack_23_clock = clock;
  assign Stack_23_reset = reset;
  assign Stack_23_io_push = LUT_stack_io_push_23; // @[stackmanage_35.scala 176:38]
  assign Stack_23_io_pop = LUT_stack_io_pop_23; // @[stackmanage_35.scala 137:39]
  assign Stack_23_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_617); // @[stackmanage_35.scala 383:64 stackmanage_35.scala 407:31]
  assign Stack_23_io_clear = LUT_stack_io_clear_23; // @[stackmanage_35.scala 217:39]
  assign Stack_23_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1865; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1734:28]
  assign Stack_23_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1864; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1733:29]
  assign Stack_24_clock = clock;
  assign Stack_24_reset = reset;
  assign Stack_24_io_push = LUT_stack_io_push_24; // @[stackmanage_35.scala 177:38]
  assign Stack_24_io_pop = LUT_stack_io_pop_24; // @[stackmanage_35.scala 138:39]
  assign Stack_24_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_618); // @[stackmanage_35.scala 383:64 stackmanage_35.scala 408:31]
  assign Stack_24_io_clear = LUT_stack_io_clear_24; // @[stackmanage_35.scala 218:39]
  assign Stack_24_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1867; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1736:28]
  assign Stack_24_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1866; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1735:29]
  assign Stack_25_clock = clock;
  assign Stack_25_reset = reset;
  assign Stack_25_io_push = LUT_stack_io_push_25; // @[stackmanage_35.scala 178:38]
  assign Stack_25_io_pop = LUT_stack_io_pop_25; // @[stackmanage_35.scala 139:39]
  assign Stack_25_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_619); // @[stackmanage_35.scala 383:64 stackmanage_35.scala 409:31]
  assign Stack_25_io_clear = LUT_stack_io_clear_25; // @[stackmanage_35.scala 219:39]
  assign Stack_25_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1869; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1738:28]
  assign Stack_25_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1868; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1737:29]
  assign Stack_26_clock = clock;
  assign Stack_26_reset = reset;
  assign Stack_26_io_push = LUT_stack_io_push_26; // @[stackmanage_35.scala 179:38]
  assign Stack_26_io_pop = LUT_stack_io_pop_26; // @[stackmanage_35.scala 140:39]
  assign Stack_26_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_620); // @[stackmanage_35.scala 383:64 stackmanage_35.scala 410:31]
  assign Stack_26_io_clear = LUT_stack_io_clear_26; // @[stackmanage_35.scala 220:39]
  assign Stack_26_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1871; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1740:28]
  assign Stack_26_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1870; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1739:29]
  assign Stack_27_clock = clock;
  assign Stack_27_reset = reset;
  assign Stack_27_io_push = LUT_stack_io_push_27; // @[stackmanage_35.scala 180:38]
  assign Stack_27_io_pop = LUT_stack_io_pop_27; // @[stackmanage_35.scala 141:39]
  assign Stack_27_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_621); // @[stackmanage_35.scala 383:64 stackmanage_35.scala 411:31]
  assign Stack_27_io_clear = LUT_stack_io_clear_27; // @[stackmanage_35.scala 221:39]
  assign Stack_27_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1873; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1742:28]
  assign Stack_27_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1872; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1741:29]
  assign Stack_28_clock = clock;
  assign Stack_28_reset = reset;
  assign Stack_28_io_push = LUT_stack_io_push_28; // @[stackmanage_35.scala 181:38]
  assign Stack_28_io_pop = LUT_stack_io_pop_28; // @[stackmanage_35.scala 142:39]
  assign Stack_28_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_622); // @[stackmanage_35.scala 383:64 stackmanage_35.scala 412:31]
  assign Stack_28_io_clear = LUT_stack_io_clear_28; // @[stackmanage_35.scala 222:39]
  assign Stack_28_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1875; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1744:28]
  assign Stack_28_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1874; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1743:29]
  assign Stack_29_clock = clock;
  assign Stack_29_reset = reset;
  assign Stack_29_io_push = LUT_stack_io_push_29; // @[stackmanage_35.scala 182:38]
  assign Stack_29_io_pop = LUT_stack_io_pop_29; // @[stackmanage_35.scala 143:39]
  assign Stack_29_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_623); // @[stackmanage_35.scala 383:64 stackmanage_35.scala 413:31]
  assign Stack_29_io_clear = LUT_stack_io_clear_29; // @[stackmanage_35.scala 223:39]
  assign Stack_29_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1877; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1746:28]
  assign Stack_29_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1876; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1745:29]
  assign Stack_30_clock = clock;
  assign Stack_30_reset = reset;
  assign Stack_30_io_push = LUT_stack_io_push_30; // @[stackmanage_35.scala 184:38]
  assign Stack_30_io_pop = LUT_stack_io_pop_30; // @[stackmanage_35.scala 145:39]
  assign Stack_30_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_624); // @[stackmanage_35.scala 383:64 stackmanage_35.scala 414:31]
  assign Stack_30_io_clear = LUT_stack_io_clear_30; // @[stackmanage_35.scala 225:39]
  assign Stack_30_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1879; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1748:29]
  assign Stack_30_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1878; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1747:29]
  assign Stack_31_clock = clock;
  assign Stack_31_reset = reset;
  assign Stack_31_io_push = LUT_stack_io_push_31; // @[stackmanage_35.scala 185:38]
  assign Stack_31_io_pop = LUT_stack_io_pop_31; // @[stackmanage_35.scala 146:39]
  assign Stack_31_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_625); // @[stackmanage_35.scala 383:64 stackmanage_35.scala 415:31]
  assign Stack_31_io_clear = LUT_stack_io_clear_31; // @[stackmanage_35.scala 226:39]
  assign Stack_31_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1881; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1750:28]
  assign Stack_31_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1880; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1749:29]
  assign Stack_32_clock = clock;
  assign Stack_32_reset = reset;
  assign Stack_32_io_push = LUT_stack_io_push_32; // @[stackmanage_35.scala 186:38]
  assign Stack_32_io_pop = LUT_stack_io_pop_32; // @[stackmanage_35.scala 147:39]
  assign Stack_32_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_626); // @[stackmanage_35.scala 383:64 stackmanage_35.scala 416:31]
  assign Stack_32_io_clear = LUT_stack_io_clear_32; // @[stackmanage_35.scala 227:39]
  assign Stack_32_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1883; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1752:28]
  assign Stack_32_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1882; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1751:29]
  assign Stack_33_clock = clock;
  assign Stack_33_reset = reset;
  assign Stack_33_io_push = LUT_stack_io_push_33; // @[stackmanage_35.scala 187:38]
  assign Stack_33_io_pop = LUT_stack_io_pop_33; // @[stackmanage_35.scala 148:39]
  assign Stack_33_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_627); // @[stackmanage_35.scala 383:64 stackmanage_35.scala 417:31]
  assign Stack_33_io_clear = LUT_stack_io_clear_33; // @[stackmanage_35.scala 228:39]
  assign Stack_33_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1885; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1754:28]
  assign Stack_33_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1884; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1753:29]
  assign Stack_34_clock = clock;
  assign Stack_34_reset = reset;
  assign Stack_34_io_push = LUT_stack_io_push_34; // @[stackmanage_35.scala 188:38]
  assign Stack_34_io_pop = LUT_stack_io_pop_34; // @[stackmanage_35.scala 149:39]
  assign Stack_34_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_628); // @[stackmanage_35.scala 383:64 stackmanage_35.scala 418:31]
  assign Stack_34_io_clear = LUT_stack_io_clear_34; // @[stackmanage_35.scala 229:39]
  assign Stack_34_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1887; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1756:28]
  assign Stack_34_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1886; // @[stackmanage_35.scala 1686:63 stackmanage_35.scala 1755:29]
  always @(posedge clock) begin
    if (reset) begin // @[stackmanage_35.scala 375:34]
      node_push_in_1 <= 32'sh0; // @[stackmanage_35.scala 375:34]
    end else begin
      node_push_in_1 <= LUT_stack_io_node_id_push_in; // @[stackmanage_35.scala 379:29]
    end
    if (reset) begin // @[stackmanage_35.scala 376:34]
      node_push_in_2 <= 32'sh0; // @[stackmanage_35.scala 376:34]
    end else begin
      node_push_in_2 <= node_push_in_1; // @[stackmanage_35.scala 380:29]
    end
    if (reset) begin // @[stackmanage_35.scala 1682:34]
      hitT_out_temp <= 32'h0; // @[stackmanage_35.scala 1682:34]
    end else if (pop_0 & Stack_0_io_enable) begin // @[stackmanage_35.scala 4332:48]
      hitT_out_temp <= Stack_0_io_hit_out; // @[stackmanage_35.scala 4334:27]
    end else if (pop_1 & Stack_1_io_enable) begin // @[stackmanage_35.scala 4338:53]
      hitT_out_temp <= Stack_1_io_hit_out; // @[stackmanage_35.scala 4339:27]
    end else if (pop_2 & Stack_2_io_enable) begin // @[stackmanage_35.scala 4343:53]
      hitT_out_temp <= Stack_2_io_hit_out; // @[stackmanage_35.scala 4344:27]
    end else begin
      hitT_out_temp <= _GEN_2082;
    end
    if (reset) begin // @[stackmanage_35.scala 1683:35]
      ray_out_temp <= 32'h0; // @[stackmanage_35.scala 1683:35]
    end else if (pop_0 & Stack_0_io_enable) begin // @[stackmanage_35.scala 4332:48]
      ray_out_temp <= Stack_0_io_ray_out; // @[stackmanage_35.scala 4335:28]
    end else if (pop_1 & Stack_1_io_enable) begin // @[stackmanage_35.scala 4338:53]
      ray_out_temp <= Stack_1_io_ray_out; // @[stackmanage_35.scala 4340:28]
    end else if (pop_2 & Stack_2_io_enable) begin // @[stackmanage_35.scala 4343:53]
      ray_out_temp <= Stack_2_io_ray_out; // @[stackmanage_35.scala 4345:28]
    end else begin
      ray_out_temp <= _GEN_2083;
    end
    if (reset) begin // @[stackmanage_35.scala 1684:32]
      node_out_temp <= 32'sh0; // @[stackmanage_35.scala 1684:32]
    end else if (pop_0 & Stack_0_io_enable) begin // @[stackmanage_35.scala 4332:48]
      node_out_temp <= Stack_0_io_dataOut; // @[stackmanage_35.scala 4336:25]
    end else if (pop_1 & Stack_1_io_enable) begin // @[stackmanage_35.scala 4338:53]
      node_out_temp <= Stack_1_io_dataOut; // @[stackmanage_35.scala 4341:25]
    end else if (pop_2 & Stack_2_io_enable) begin // @[stackmanage_35.scala 4343:53]
      node_out_temp <= Stack_2_io_dataOut; // @[stackmanage_35.scala 4346:25]
    end else begin
      node_out_temp <= _GEN_2084;
    end
    if (reset) begin // @[stackmanage_35.scala 1685:38]
      pop_valid_1 <= 1'h0; // @[stackmanage_35.scala 1685:38]
    end else begin
      pop_valid_1 <= _GEN_2097;
    end
    if (reset) begin // @[stackmanage_35.scala 4245:46]
      pop_0 <= 1'h0; // @[stackmanage_35.scala 4245:46]
    end else begin
      pop_0 <= LUT_stack_io_pop_0; // @[stackmanage_35.scala 4295:40]
    end
    if (reset) begin // @[stackmanage_35.scala 4246:46]
      pop_1 <= 1'h0; // @[stackmanage_35.scala 4246:46]
    end else begin
      pop_1 <= LUT_stack_io_pop_1; // @[stackmanage_35.scala 4296:40]
    end
    if (reset) begin // @[stackmanage_35.scala 4247:46]
      pop_2 <= 1'h0; // @[stackmanage_35.scala 4247:46]
    end else begin
      pop_2 <= LUT_stack_io_pop_2; // @[stackmanage_35.scala 4297:40]
    end
    if (reset) begin // @[stackmanage_35.scala 4248:46]
      pop_3 <= 1'h0; // @[stackmanage_35.scala 4248:46]
    end else begin
      pop_3 <= LUT_stack_io_pop_3; // @[stackmanage_35.scala 4298:40]
    end
    if (reset) begin // @[stackmanage_35.scala 4249:46]
      pop_4 <= 1'h0; // @[stackmanage_35.scala 4249:46]
    end else begin
      pop_4 <= LUT_stack_io_pop_4; // @[stackmanage_35.scala 4299:40]
    end
    if (reset) begin // @[stackmanage_35.scala 4250:46]
      pop_5 <= 1'h0; // @[stackmanage_35.scala 4250:46]
    end else begin
      pop_5 <= LUT_stack_io_pop_5; // @[stackmanage_35.scala 4300:40]
    end
    if (reset) begin // @[stackmanage_35.scala 4251:46]
      pop_6 <= 1'h0; // @[stackmanage_35.scala 4251:46]
    end else begin
      pop_6 <= LUT_stack_io_pop_6; // @[stackmanage_35.scala 4301:40]
    end
    if (reset) begin // @[stackmanage_35.scala 4252:46]
      pop_7 <= 1'h0; // @[stackmanage_35.scala 4252:46]
    end else begin
      pop_7 <= LUT_stack_io_pop_7; // @[stackmanage_35.scala 4302:40]
    end
    if (reset) begin // @[stackmanage_35.scala 4253:46]
      pop_8 <= 1'h0; // @[stackmanage_35.scala 4253:46]
    end else begin
      pop_8 <= LUT_stack_io_pop_8; // @[stackmanage_35.scala 4303:40]
    end
    if (reset) begin // @[stackmanage_35.scala 4254:46]
      pop_9 <= 1'h0; // @[stackmanage_35.scala 4254:46]
    end else begin
      pop_9 <= LUT_stack_io_pop_9; // @[stackmanage_35.scala 4304:40]
    end
    if (reset) begin // @[stackmanage_35.scala 4256:47]
      pop_10 <= 1'h0; // @[stackmanage_35.scala 4256:47]
    end else begin
      pop_10 <= LUT_stack_io_pop_10; // @[stackmanage_35.scala 4305:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4257:47]
      pop_11 <= 1'h0; // @[stackmanage_35.scala 4257:47]
    end else begin
      pop_11 <= LUT_stack_io_pop_11; // @[stackmanage_35.scala 4306:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4258:47]
      pop_12 <= 1'h0; // @[stackmanage_35.scala 4258:47]
    end else begin
      pop_12 <= LUT_stack_io_pop_12; // @[stackmanage_35.scala 4307:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4259:47]
      pop_13 <= 1'h0; // @[stackmanage_35.scala 4259:47]
    end else begin
      pop_13 <= LUT_stack_io_pop_13; // @[stackmanage_35.scala 4308:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4260:47]
      pop_14 <= 1'h0; // @[stackmanage_35.scala 4260:47]
    end else begin
      pop_14 <= LUT_stack_io_pop_14; // @[stackmanage_35.scala 4309:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4261:47]
      pop_15 <= 1'h0; // @[stackmanage_35.scala 4261:47]
    end else begin
      pop_15 <= LUT_stack_io_pop_15; // @[stackmanage_35.scala 4310:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4262:47]
      pop_16 <= 1'h0; // @[stackmanage_35.scala 4262:47]
    end else begin
      pop_16 <= LUT_stack_io_pop_16; // @[stackmanage_35.scala 4311:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4263:47]
      pop_17 <= 1'h0; // @[stackmanage_35.scala 4263:47]
    end else begin
      pop_17 <= LUT_stack_io_pop_17; // @[stackmanage_35.scala 4312:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4264:47]
      pop_18 <= 1'h0; // @[stackmanage_35.scala 4264:47]
    end else begin
      pop_18 <= LUT_stack_io_pop_18; // @[stackmanage_35.scala 4313:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4265:47]
      pop_19 <= 1'h0; // @[stackmanage_35.scala 4265:47]
    end else begin
      pop_19 <= LUT_stack_io_pop_19; // @[stackmanage_35.scala 4314:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4267:47]
      pop_20 <= 1'h0; // @[stackmanage_35.scala 4267:47]
    end else begin
      pop_20 <= LUT_stack_io_pop_20; // @[stackmanage_35.scala 4315:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4268:47]
      pop_21 <= 1'h0; // @[stackmanage_35.scala 4268:47]
    end else begin
      pop_21 <= LUT_stack_io_pop_21; // @[stackmanage_35.scala 4316:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4269:47]
      pop_22 <= 1'h0; // @[stackmanage_35.scala 4269:47]
    end else begin
      pop_22 <= LUT_stack_io_pop_22; // @[stackmanage_35.scala 4317:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4270:47]
      pop_23 <= 1'h0; // @[stackmanage_35.scala 4270:47]
    end else begin
      pop_23 <= LUT_stack_io_pop_23; // @[stackmanage_35.scala 4318:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4271:47]
      pop_24 <= 1'h0; // @[stackmanage_35.scala 4271:47]
    end else begin
      pop_24 <= LUT_stack_io_pop_24; // @[stackmanage_35.scala 4319:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4272:47]
      pop_25 <= 1'h0; // @[stackmanage_35.scala 4272:47]
    end else begin
      pop_25 <= LUT_stack_io_pop_25; // @[stackmanage_35.scala 4320:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4273:47]
      pop_26 <= 1'h0; // @[stackmanage_35.scala 4273:47]
    end else begin
      pop_26 <= LUT_stack_io_pop_26; // @[stackmanage_35.scala 4321:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4274:47]
      pop_27 <= 1'h0; // @[stackmanage_35.scala 4274:47]
    end else begin
      pop_27 <= LUT_stack_io_pop_27; // @[stackmanage_35.scala 4322:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4275:47]
      pop_28 <= 1'h0; // @[stackmanage_35.scala 4275:47]
    end else begin
      pop_28 <= LUT_stack_io_pop_28; // @[stackmanage_35.scala 4323:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4276:47]
      pop_29 <= 1'h0; // @[stackmanage_35.scala 4276:47]
    end else begin
      pop_29 <= LUT_stack_io_pop_29; // @[stackmanage_35.scala 4324:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4278:47]
      pop_30 <= 1'h0; // @[stackmanage_35.scala 4278:47]
    end else begin
      pop_30 <= LUT_stack_io_pop_30; // @[stackmanage_35.scala 4325:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4279:47]
      pop_31 <= 1'h0; // @[stackmanage_35.scala 4279:47]
    end else begin
      pop_31 <= LUT_stack_io_pop_31; // @[stackmanage_35.scala 4326:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4280:47]
      pop_32 <= 1'h0; // @[stackmanage_35.scala 4280:47]
    end else begin
      pop_32 <= LUT_stack_io_pop_32; // @[stackmanage_35.scala 4327:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4281:47]
      pop_33 <= 1'h0; // @[stackmanage_35.scala 4281:47]
    end else begin
      pop_33 <= LUT_stack_io_pop_33; // @[stackmanage_35.scala 4328:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4282:47]
      pop_34 <= 1'h0; // @[stackmanage_35.scala 4282:47]
    end else begin
      pop_34 <= LUT_stack_io_pop_34; // @[stackmanage_35.scala 4329:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4520:41]
      dispatch_0 <= 1'h0; // @[stackmanage_35.scala 4520:41]
    end else begin
      dispatch_0 <= _T_317;
    end
    if (reset) begin // @[stackmanage_35.scala 4521:41]
      dispatch_1 <= 1'h0; // @[stackmanage_35.scala 4521:41]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4643:38]
      dispatch_1 <= 1'h0; // @[stackmanage_35.scala 4645:33]
    end else begin
      dispatch_1 <= _T_320;
    end
    if (reset) begin // @[stackmanage_35.scala 4522:41]
      dispatch_2 <= 1'h0; // @[stackmanage_35.scala 4522:41]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4643:38]
      dispatch_2 <= 1'h0; // @[stackmanage_35.scala 4646:33]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4679:43]
      dispatch_2 <= 1'h0; // @[stackmanage_35.scala 4682:33]
    end else begin
      dispatch_2 <= _T_323;
    end
    if (reset) begin // @[stackmanage_35.scala 4523:41]
      dispatch_3 <= 1'h0; // @[stackmanage_35.scala 4523:41]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4643:38]
      dispatch_3 <= 1'h0; // @[stackmanage_35.scala 4647:33]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4679:43]
      dispatch_3 <= 1'h0; // @[stackmanage_35.scala 4683:33]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4716:43]
      dispatch_3 <= 1'h0; // @[stackmanage_35.scala 4720:33]
    end else begin
      dispatch_3 <= _T_326;
    end
    if (reset) begin // @[stackmanage_35.scala 4524:41]
      dispatch_4 <= 1'h0; // @[stackmanage_35.scala 4524:41]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4643:38]
      dispatch_4 <= 1'h0; // @[stackmanage_35.scala 4648:33]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4679:43]
      dispatch_4 <= 1'h0; // @[stackmanage_35.scala 4684:33]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4716:43]
      dispatch_4 <= 1'h0; // @[stackmanage_35.scala 4722:33]
    end else begin
      dispatch_4 <= _GEN_2627;
    end
    if (reset) begin // @[stackmanage_35.scala 4525:41]
      dispatch_5 <= 1'h0; // @[stackmanage_35.scala 4525:41]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4643:38]
      dispatch_5 <= 1'h0; // @[stackmanage_35.scala 4649:33]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4679:43]
      dispatch_5 <= 1'h0; // @[stackmanage_35.scala 4685:33]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4716:43]
      dispatch_5 <= 1'h0; // @[stackmanage_35.scala 4723:33]
    end else begin
      dispatch_5 <= _GEN_2628;
    end
    if (reset) begin // @[stackmanage_35.scala 4526:41]
      dispatch_6 <= 1'h0; // @[stackmanage_35.scala 4526:41]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4643:38]
      dispatch_6 <= 1'h0; // @[stackmanage_35.scala 4650:33]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4679:43]
      dispatch_6 <= 1'h0; // @[stackmanage_35.scala 4686:33]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4716:43]
      dispatch_6 <= 1'h0; // @[stackmanage_35.scala 4724:33]
    end else begin
      dispatch_6 <= _GEN_2629;
    end
    if (reset) begin // @[stackmanage_35.scala 4527:41]
      dispatch_7 <= 1'h0; // @[stackmanage_35.scala 4527:41]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4643:38]
      dispatch_7 <= 1'h0; // @[stackmanage_35.scala 4651:33]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4679:43]
      dispatch_7 <= 1'h0; // @[stackmanage_35.scala 4687:33]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4716:43]
      dispatch_7 <= 1'h0; // @[stackmanage_35.scala 4725:33]
    end else begin
      dispatch_7 <= _GEN_2630;
    end
    if (reset) begin // @[stackmanage_35.scala 4528:41]
      dispatch_8 <= 1'h0; // @[stackmanage_35.scala 4528:41]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4643:38]
      dispatch_8 <= 1'h0; // @[stackmanage_35.scala 4652:33]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4679:43]
      dispatch_8 <= 1'h0; // @[stackmanage_35.scala 4688:33]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4716:43]
      dispatch_8 <= 1'h0; // @[stackmanage_35.scala 4726:33]
    end else begin
      dispatch_8 <= _GEN_2631;
    end
    if (reset) begin // @[stackmanage_35.scala 4529:41]
      dispatch_9 <= 1'h0; // @[stackmanage_35.scala 4529:41]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4643:38]
      dispatch_9 <= 1'h0; // @[stackmanage_35.scala 4653:33]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4679:43]
      dispatch_9 <= 1'h0; // @[stackmanage_35.scala 4689:33]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4716:43]
      dispatch_9 <= 1'h0; // @[stackmanage_35.scala 4727:33]
    end else begin
      dispatch_9 <= _GEN_2632;
    end
    if (reset) begin // @[stackmanage_35.scala 4531:42]
      dispatch_10 <= 1'h0; // @[stackmanage_35.scala 4531:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4643:38]
      dispatch_10 <= 1'h0; // @[stackmanage_35.scala 4654:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4679:43]
      dispatch_10 <= 1'h0; // @[stackmanage_35.scala 4690:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4716:43]
      dispatch_10 <= 1'h0; // @[stackmanage_35.scala 4728:34]
    end else begin
      dispatch_10 <= _GEN_2633;
    end
    if (reset) begin // @[stackmanage_35.scala 4532:42]
      dispatch_11 <= 1'h0; // @[stackmanage_35.scala 4532:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4643:38]
      dispatch_11 <= 1'h0; // @[stackmanage_35.scala 4655:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4679:43]
      dispatch_11 <= 1'h0; // @[stackmanage_35.scala 4691:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4716:43]
      dispatch_11 <= 1'h0; // @[stackmanage_35.scala 4729:34]
    end else begin
      dispatch_11 <= _GEN_2634;
    end
    if (reset) begin // @[stackmanage_35.scala 4533:42]
      dispatch_12 <= 1'h0; // @[stackmanage_35.scala 4533:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4643:38]
      dispatch_12 <= 1'h0; // @[stackmanage_35.scala 4656:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4679:43]
      dispatch_12 <= 1'h0; // @[stackmanage_35.scala 4692:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4716:43]
      dispatch_12 <= 1'h0; // @[stackmanage_35.scala 4730:34]
    end else begin
      dispatch_12 <= _GEN_2635;
    end
    if (reset) begin // @[stackmanage_35.scala 4534:42]
      dispatch_13 <= 1'h0; // @[stackmanage_35.scala 4534:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4643:38]
      dispatch_13 <= 1'h0; // @[stackmanage_35.scala 4657:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4679:43]
      dispatch_13 <= 1'h0; // @[stackmanage_35.scala 4693:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4716:43]
      dispatch_13 <= 1'h0; // @[stackmanage_35.scala 4731:34]
    end else begin
      dispatch_13 <= _GEN_2636;
    end
    if (reset) begin // @[stackmanage_35.scala 4535:42]
      dispatch_14 <= 1'h0; // @[stackmanage_35.scala 4535:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4643:38]
      dispatch_14 <= 1'h0; // @[stackmanage_35.scala 4658:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4679:43]
      dispatch_14 <= 1'h0; // @[stackmanage_35.scala 4694:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4716:43]
      dispatch_14 <= 1'h0; // @[stackmanage_35.scala 4732:34]
    end else begin
      dispatch_14 <= _GEN_2637;
    end
    if (reset) begin // @[stackmanage_35.scala 4536:42]
      dispatch_15 <= 1'h0; // @[stackmanage_35.scala 4536:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4643:38]
      dispatch_15 <= 1'h0; // @[stackmanage_35.scala 4659:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4679:43]
      dispatch_15 <= 1'h0; // @[stackmanage_35.scala 4695:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4716:43]
      dispatch_15 <= 1'h0; // @[stackmanage_35.scala 4733:34]
    end else begin
      dispatch_15 <= _GEN_2638;
    end
    if (reset) begin // @[stackmanage_35.scala 4537:42]
      dispatch_16 <= 1'h0; // @[stackmanage_35.scala 4537:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4643:38]
      dispatch_16 <= 1'h0; // @[stackmanage_35.scala 4660:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4679:43]
      dispatch_16 <= 1'h0; // @[stackmanage_35.scala 4696:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4716:43]
      dispatch_16 <= 1'h0; // @[stackmanage_35.scala 4734:34]
    end else begin
      dispatch_16 <= _GEN_2639;
    end
    if (reset) begin // @[stackmanage_35.scala 4538:42]
      dispatch_17 <= 1'h0; // @[stackmanage_35.scala 4538:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4643:38]
      dispatch_17 <= 1'h0; // @[stackmanage_35.scala 4661:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4679:43]
      dispatch_17 <= 1'h0; // @[stackmanage_35.scala 4697:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4716:43]
      dispatch_17 <= 1'h0; // @[stackmanage_35.scala 4735:34]
    end else begin
      dispatch_17 <= _GEN_2640;
    end
    if (reset) begin // @[stackmanage_35.scala 4539:42]
      dispatch_18 <= 1'h0; // @[stackmanage_35.scala 4539:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4643:38]
      dispatch_18 <= 1'h0; // @[stackmanage_35.scala 4662:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4679:43]
      dispatch_18 <= 1'h0; // @[stackmanage_35.scala 4698:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4716:43]
      dispatch_18 <= 1'h0; // @[stackmanage_35.scala 4736:34]
    end else begin
      dispatch_18 <= _GEN_2641;
    end
    if (reset) begin // @[stackmanage_35.scala 4540:42]
      dispatch_19 <= 1'h0; // @[stackmanage_35.scala 4540:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4643:38]
      dispatch_19 <= 1'h0; // @[stackmanage_35.scala 4663:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4679:43]
      dispatch_19 <= 1'h0; // @[stackmanage_35.scala 4699:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4716:43]
      dispatch_19 <= 1'h0; // @[stackmanage_35.scala 4737:34]
    end else begin
      dispatch_19 <= _GEN_2642;
    end
    if (reset) begin // @[stackmanage_35.scala 4542:42]
      dispatch_20 <= 1'h0; // @[stackmanage_35.scala 4542:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4643:38]
      dispatch_20 <= 1'h0; // @[stackmanage_35.scala 4664:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4679:43]
      dispatch_20 <= 1'h0; // @[stackmanage_35.scala 4700:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4716:43]
      dispatch_20 <= 1'h0; // @[stackmanage_35.scala 4738:34]
    end else begin
      dispatch_20 <= _GEN_2643;
    end
    if (reset) begin // @[stackmanage_35.scala 4543:42]
      dispatch_21 <= 1'h0; // @[stackmanage_35.scala 4543:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4643:38]
      dispatch_21 <= 1'h0; // @[stackmanage_35.scala 4665:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4679:43]
      dispatch_21 <= 1'h0; // @[stackmanage_35.scala 4701:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4716:43]
      dispatch_21 <= 1'h0; // @[stackmanage_35.scala 4739:34]
    end else begin
      dispatch_21 <= _GEN_2644;
    end
    if (reset) begin // @[stackmanage_35.scala 4544:42]
      dispatch_22 <= 1'h0; // @[stackmanage_35.scala 4544:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4643:38]
      dispatch_22 <= 1'h0; // @[stackmanage_35.scala 4666:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4679:43]
      dispatch_22 <= 1'h0; // @[stackmanage_35.scala 4702:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4716:43]
      dispatch_22 <= 1'h0; // @[stackmanage_35.scala 4740:34]
    end else begin
      dispatch_22 <= _GEN_2645;
    end
    if (reset) begin // @[stackmanage_35.scala 4545:42]
      dispatch_23 <= 1'h0; // @[stackmanage_35.scala 4545:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4643:38]
      dispatch_23 <= 1'h0; // @[stackmanage_35.scala 4667:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4679:43]
      dispatch_23 <= 1'h0; // @[stackmanage_35.scala 4703:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4716:43]
      dispatch_23 <= 1'h0; // @[stackmanage_35.scala 4741:34]
    end else begin
      dispatch_23 <= _GEN_2646;
    end
    if (reset) begin // @[stackmanage_35.scala 4546:42]
      dispatch_24 <= 1'h0; // @[stackmanage_35.scala 4546:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4643:38]
      dispatch_24 <= 1'h0; // @[stackmanage_35.scala 4668:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4679:43]
      dispatch_24 <= 1'h0; // @[stackmanage_35.scala 4704:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4716:43]
      dispatch_24 <= 1'h0; // @[stackmanage_35.scala 4742:34]
    end else begin
      dispatch_24 <= _GEN_2647;
    end
    if (reset) begin // @[stackmanage_35.scala 4547:42]
      dispatch_25 <= 1'h0; // @[stackmanage_35.scala 4547:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4643:38]
      dispatch_25 <= 1'h0; // @[stackmanage_35.scala 4669:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4679:43]
      dispatch_25 <= 1'h0; // @[stackmanage_35.scala 4705:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4716:43]
      dispatch_25 <= 1'h0; // @[stackmanage_35.scala 4743:34]
    end else begin
      dispatch_25 <= _GEN_2648;
    end
    if (reset) begin // @[stackmanage_35.scala 4548:42]
      dispatch_26 <= 1'h0; // @[stackmanage_35.scala 4548:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4643:38]
      dispatch_26 <= 1'h0; // @[stackmanage_35.scala 4670:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4679:43]
      dispatch_26 <= 1'h0; // @[stackmanage_35.scala 4706:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4716:43]
      dispatch_26 <= 1'h0; // @[stackmanage_35.scala 4744:34]
    end else begin
      dispatch_26 <= _GEN_2649;
    end
    if (reset) begin // @[stackmanage_35.scala 4549:42]
      dispatch_27 <= 1'h0; // @[stackmanage_35.scala 4549:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4643:38]
      dispatch_27 <= 1'h0; // @[stackmanage_35.scala 4671:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4679:43]
      dispatch_27 <= 1'h0; // @[stackmanage_35.scala 4707:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4716:43]
      dispatch_27 <= 1'h0; // @[stackmanage_35.scala 4745:34]
    end else begin
      dispatch_27 <= _GEN_2650;
    end
    if (reset) begin // @[stackmanage_35.scala 4550:42]
      dispatch_28 <= 1'h0; // @[stackmanage_35.scala 4550:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4643:38]
      dispatch_28 <= 1'h0; // @[stackmanage_35.scala 4672:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4679:43]
      dispatch_28 <= 1'h0; // @[stackmanage_35.scala 4708:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4716:43]
      dispatch_28 <= 1'h0; // @[stackmanage_35.scala 4746:34]
    end else begin
      dispatch_28 <= _GEN_2651;
    end
    if (reset) begin // @[stackmanage_35.scala 4551:42]
      dispatch_29 <= 1'h0; // @[stackmanage_35.scala 4551:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4643:38]
      dispatch_29 <= 1'h0; // @[stackmanage_35.scala 4673:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4679:43]
      dispatch_29 <= 1'h0; // @[stackmanage_35.scala 4709:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4716:43]
      dispatch_29 <= 1'h0; // @[stackmanage_35.scala 4747:34]
    end else begin
      dispatch_29 <= _GEN_2652;
    end
    if (reset) begin // @[stackmanage_35.scala 4553:42]
      dispatch_30 <= 1'h0; // @[stackmanage_35.scala 4553:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4643:38]
      dispatch_30 <= 1'h0; // @[stackmanage_35.scala 4674:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4679:43]
      dispatch_30 <= 1'h0; // @[stackmanage_35.scala 4710:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4716:43]
      dispatch_30 <= 1'h0; // @[stackmanage_35.scala 4748:34]
    end else begin
      dispatch_30 <= _GEN_2653;
    end
    if (reset) begin // @[stackmanage_35.scala 4554:42]
      dispatch_31 <= 1'h0; // @[stackmanage_35.scala 4554:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4643:38]
      dispatch_31 <= 1'h0; // @[stackmanage_35.scala 4675:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4679:43]
      dispatch_31 <= 1'h0; // @[stackmanage_35.scala 4711:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4716:43]
      dispatch_31 <= 1'h0; // @[stackmanage_35.scala 4749:34]
    end else begin
      dispatch_31 <= _GEN_2654;
    end
    if (reset) begin // @[stackmanage_35.scala 4555:42]
      dispatch_32 <= 1'h0; // @[stackmanage_35.scala 4555:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4643:38]
      dispatch_32 <= 1'h0; // @[stackmanage_35.scala 4676:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4679:43]
      dispatch_32 <= 1'h0; // @[stackmanage_35.scala 4712:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4716:43]
      dispatch_32 <= 1'h0; // @[stackmanage_35.scala 4750:34]
    end else begin
      dispatch_32 <= _GEN_2655;
    end
    if (reset) begin // @[stackmanage_35.scala 4556:42]
      dispatch_33 <= 1'h0; // @[stackmanage_35.scala 4556:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4643:38]
      dispatch_33 <= 1'h0; // @[stackmanage_35.scala 4677:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4679:43]
      dispatch_33 <= 1'h0; // @[stackmanage_35.scala 4713:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4716:43]
      dispatch_33 <= 1'h0; // @[stackmanage_35.scala 4751:34]
    end else begin
      dispatch_33 <= _GEN_2656;
    end
    if (reset) begin // @[stackmanage_35.scala 4557:42]
      dispatch_34 <= 1'h0; // @[stackmanage_35.scala 4557:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4643:38]
      dispatch_34 <= 1'h0; // @[stackmanage_35.scala 4678:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4679:43]
      dispatch_34 <= 1'h0; // @[stackmanage_35.scala 4714:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4716:43]
      dispatch_34 <= 1'h0; // @[stackmanage_35.scala 4752:34]
    end else begin
      dispatch_34 <= _GEN_2657;
    end
    if (reset) begin // @[stackmanage_35.scala 4558:42]
      dispatch_no_match <= 1'h0; // @[stackmanage_35.scala 4558:42]
    end else begin
      dispatch_no_match <= LUT_stack_io_no_match; // @[stackmanage_35.scala 5984:25]
    end
    if (reset) begin // @[stackmanage_35.scala 4562:42]
      empty_0 <= 1'h0; // @[stackmanage_35.scala 4562:42]
    end else begin
      empty_0 <= Stack_0_io_empty; // @[stackmanage_35.scala 4601:35]
    end
    if (reset) begin // @[stackmanage_35.scala 4563:42]
      empty_1 <= 1'h0; // @[stackmanage_35.scala 4563:42]
    end else begin
      empty_1 <= Stack_1_io_empty; // @[stackmanage_35.scala 4602:35]
    end
    if (reset) begin // @[stackmanage_35.scala 4564:42]
      empty_2 <= 1'h0; // @[stackmanage_35.scala 4564:42]
    end else begin
      empty_2 <= Stack_2_io_empty; // @[stackmanage_35.scala 4603:35]
    end
    if (reset) begin // @[stackmanage_35.scala 4565:42]
      empty_3 <= 1'h0; // @[stackmanage_35.scala 4565:42]
    end else begin
      empty_3 <= Stack_3_io_empty; // @[stackmanage_35.scala 4604:35]
    end
    if (reset) begin // @[stackmanage_35.scala 4566:42]
      empty_4 <= 1'h0; // @[stackmanage_35.scala 4566:42]
    end else begin
      empty_4 <= Stack_4_io_empty; // @[stackmanage_35.scala 4605:35]
    end
    if (reset) begin // @[stackmanage_35.scala 4567:42]
      empty_5 <= 1'h0; // @[stackmanage_35.scala 4567:42]
    end else begin
      empty_5 <= Stack_5_io_empty; // @[stackmanage_35.scala 4606:35]
    end
    if (reset) begin // @[stackmanage_35.scala 4568:42]
      empty_6 <= 1'h0; // @[stackmanage_35.scala 4568:42]
    end else begin
      empty_6 <= Stack_6_io_empty; // @[stackmanage_35.scala 4607:35]
    end
    if (reset) begin // @[stackmanage_35.scala 4569:42]
      empty_7 <= 1'h0; // @[stackmanage_35.scala 4569:42]
    end else begin
      empty_7 <= Stack_7_io_empty; // @[stackmanage_35.scala 4608:35]
    end
    if (reset) begin // @[stackmanage_35.scala 4570:42]
      empty_8 <= 1'h0; // @[stackmanage_35.scala 4570:42]
    end else begin
      empty_8 <= Stack_8_io_empty; // @[stackmanage_35.scala 4609:35]
    end
    if (reset) begin // @[stackmanage_35.scala 4571:42]
      empty_9 <= 1'h0; // @[stackmanage_35.scala 4571:42]
    end else begin
      empty_9 <= Stack_9_io_empty; // @[stackmanage_35.scala 4610:35]
    end
    if (reset) begin // @[stackmanage_35.scala 4573:43]
      empty_10 <= 1'h0; // @[stackmanage_35.scala 4573:43]
    end else begin
      empty_10 <= Stack_10_io_empty; // @[stackmanage_35.scala 4612:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4574:43]
      empty_11 <= 1'h0; // @[stackmanage_35.scala 4574:43]
    end else begin
      empty_11 <= Stack_11_io_empty; // @[stackmanage_35.scala 4613:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4575:43]
      empty_12 <= 1'h0; // @[stackmanage_35.scala 4575:43]
    end else begin
      empty_12 <= Stack_12_io_empty; // @[stackmanage_35.scala 4614:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4576:43]
      empty_13 <= 1'h0; // @[stackmanage_35.scala 4576:43]
    end else begin
      empty_13 <= Stack_13_io_empty; // @[stackmanage_35.scala 4615:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4577:43]
      empty_14 <= 1'h0; // @[stackmanage_35.scala 4577:43]
    end else begin
      empty_14 <= Stack_14_io_empty; // @[stackmanage_35.scala 4616:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4578:43]
      empty_15 <= 1'h0; // @[stackmanage_35.scala 4578:43]
    end else begin
      empty_15 <= Stack_15_io_empty; // @[stackmanage_35.scala 4617:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4579:43]
      empty_16 <= 1'h0; // @[stackmanage_35.scala 4579:43]
    end else begin
      empty_16 <= Stack_16_io_empty; // @[stackmanage_35.scala 4618:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4580:43]
      empty_17 <= 1'h0; // @[stackmanage_35.scala 4580:43]
    end else begin
      empty_17 <= Stack_17_io_empty; // @[stackmanage_35.scala 4619:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4581:43]
      empty_18 <= 1'h0; // @[stackmanage_35.scala 4581:43]
    end else begin
      empty_18 <= Stack_18_io_empty; // @[stackmanage_35.scala 4620:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4582:43]
      empty_19 <= 1'h0; // @[stackmanage_35.scala 4582:43]
    end else begin
      empty_19 <= Stack_19_io_empty; // @[stackmanage_35.scala 4621:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4584:43]
      empty_20 <= 1'h0; // @[stackmanage_35.scala 4584:43]
    end else begin
      empty_20 <= Stack_20_io_empty; // @[stackmanage_35.scala 4623:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4585:43]
      empty_21 <= 1'h0; // @[stackmanage_35.scala 4585:43]
    end else begin
      empty_21 <= Stack_21_io_empty; // @[stackmanage_35.scala 4624:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4586:43]
      empty_22 <= 1'h0; // @[stackmanage_35.scala 4586:43]
    end else begin
      empty_22 <= Stack_22_io_empty; // @[stackmanage_35.scala 4625:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4587:43]
      empty_23 <= 1'h0; // @[stackmanage_35.scala 4587:43]
    end else begin
      empty_23 <= Stack_23_io_empty; // @[stackmanage_35.scala 4626:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4588:43]
      empty_24 <= 1'h0; // @[stackmanage_35.scala 4588:43]
    end else begin
      empty_24 <= Stack_24_io_empty; // @[stackmanage_35.scala 4627:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4589:43]
      empty_25 <= 1'h0; // @[stackmanage_35.scala 4589:43]
    end else begin
      empty_25 <= Stack_25_io_empty; // @[stackmanage_35.scala 4628:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4590:43]
      empty_26 <= 1'h0; // @[stackmanage_35.scala 4590:43]
    end else begin
      empty_26 <= Stack_26_io_empty; // @[stackmanage_35.scala 4629:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4591:43]
      empty_27 <= 1'h0; // @[stackmanage_35.scala 4591:43]
    end else begin
      empty_27 <= Stack_27_io_empty; // @[stackmanage_35.scala 4630:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4592:43]
      empty_28 <= 1'h0; // @[stackmanage_35.scala 4592:43]
    end else begin
      empty_28 <= Stack_28_io_empty; // @[stackmanage_35.scala 4631:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4593:43]
      empty_29 <= 1'h0; // @[stackmanage_35.scala 4593:43]
    end else begin
      empty_29 <= Stack_29_io_empty; // @[stackmanage_35.scala 4632:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4595:43]
      empty_30 <= 1'h0; // @[stackmanage_35.scala 4595:43]
    end else begin
      empty_30 <= Stack_30_io_empty; // @[stackmanage_35.scala 4634:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4596:43]
      empty_31 <= 1'h0; // @[stackmanage_35.scala 4596:43]
    end else begin
      empty_31 <= Stack_31_io_empty; // @[stackmanage_35.scala 4635:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4597:43]
      empty_32 <= 1'h0; // @[stackmanage_35.scala 4597:43]
    end else begin
      empty_32 <= Stack_32_io_empty; // @[stackmanage_35.scala 4636:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4598:43]
      empty_33 <= 1'h0; // @[stackmanage_35.scala 4598:43]
    end else begin
      empty_33 <= Stack_33_io_empty; // @[stackmanage_35.scala 4637:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4599:43]
      empty_34 <= 1'h0; // @[stackmanage_35.scala 4599:43]
    end else begin
      empty_34 <= Stack_34_io_empty; // @[stackmanage_35.scala 4638:36]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  node_push_in_1 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  node_push_in_2 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  hitT_out_temp = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  ray_out_temp = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  node_out_temp = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  pop_valid_1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  pop_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  pop_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  pop_2 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  pop_3 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  pop_4 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  pop_5 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  pop_6 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  pop_7 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  pop_8 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  pop_9 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  pop_10 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  pop_11 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  pop_12 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  pop_13 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  pop_14 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  pop_15 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  pop_16 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  pop_17 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  pop_18 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  pop_19 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  pop_20 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  pop_21 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  pop_22 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  pop_23 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  pop_24 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  pop_25 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  pop_26 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  pop_27 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  pop_28 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  pop_29 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  pop_30 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  pop_31 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  pop_32 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  pop_33 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  pop_34 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  dispatch_0 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  dispatch_1 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  dispatch_2 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  dispatch_3 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  dispatch_4 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  dispatch_5 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  dispatch_6 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  dispatch_7 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  dispatch_8 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  dispatch_9 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  dispatch_10 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  dispatch_11 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  dispatch_12 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  dispatch_13 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  dispatch_14 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  dispatch_15 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  dispatch_16 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  dispatch_17 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  dispatch_18 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  dispatch_19 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  dispatch_20 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  dispatch_21 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  dispatch_22 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  dispatch_23 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  dispatch_24 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  dispatch_25 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  dispatch_26 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  dispatch_27 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  dispatch_28 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  dispatch_29 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  dispatch_30 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  dispatch_31 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  dispatch_32 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  dispatch_33 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  dispatch_34 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  dispatch_no_match = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  empty_0 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  empty_1 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  empty_2 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  empty_3 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  empty_4 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  empty_5 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  empty_6 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  empty_7 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  empty_8 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  empty_9 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  empty_10 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  empty_11 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  empty_12 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  empty_13 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  empty_14 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  empty_15 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  empty_16 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  empty_17 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  empty_18 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  empty_19 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  empty_20 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  empty_21 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  empty_22 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  empty_23 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  empty_24 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  empty_25 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  empty_26 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  empty_27 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  empty_28 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  empty_29 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  empty_30 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  empty_31 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  empty_32 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  empty_33 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  empty_34 = _RAND_111[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MY_MUL(
  input         clock,
  input         reset,
  input  [31:0] io_a,
  input  [31:0] io_b,
  output [31:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_REG_INIT
  wire [32:0] mulAddRecFNToRaw_preMul_io_a; // @[FMUL_1.scala 36:15]
  wire [32:0] mulAddRecFNToRaw_preMul_io_b; // @[FMUL_1.scala 36:15]
  wire [32:0] mulAddRecFNToRaw_preMul_io_c; // @[FMUL_1.scala 36:15]
  wire [23:0] mulAddRecFNToRaw_preMul_io_mulAddA; // @[FMUL_1.scala 36:15]
  wire [23:0] mulAddRecFNToRaw_preMul_io_mulAddB; // @[FMUL_1.scala 36:15]
  wire [47:0] mulAddRecFNToRaw_preMul_io_mulAddC; // @[FMUL_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny; // @[FMUL_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB; // @[FMUL_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfA; // @[FMUL_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA; // @[FMUL_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfB; // @[FMUL_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB; // @[FMUL_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_signProd; // @[FMUL_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC; // @[FMUL_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfC; // @[FMUL_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC; // @[FMUL_1.scala 36:15]
  wire [9:0] mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum; // @[FMUL_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags; // @[FMUL_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant; // @[FMUL_1.scala 36:15]
  wire [4:0] mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist; // @[FMUL_1.scala 36:15]
  wire [25:0] mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC; // @[FMUL_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC; // @[FMUL_1.scala 36:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny; // @[FMUL_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB; // @[FMUL_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA; // @[FMUL_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA; // @[FMUL_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB; // @[FMUL_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB; // @[FMUL_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_signProd; // @[FMUL_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC; // @[FMUL_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC; // @[FMUL_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC; // @[FMUL_1.scala 116:15]
  wire [9:0] mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum; // @[FMUL_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags; // @[FMUL_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant; // @[FMUL_1.scala 116:15]
  wire [4:0] mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist; // @[FMUL_1.scala 116:15]
  wire [25:0] mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC; // @[FMUL_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC; // @[FMUL_1.scala 116:15]
  wire [48:0] mulAddRecFNToRaw_postMul_io_mulAddResult; // @[FMUL_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_invalidExc; // @[FMUL_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isNaN; // @[FMUL_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isInf; // @[FMUL_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isZero; // @[FMUL_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_sign; // @[FMUL_1.scala 116:15]
  wire [9:0] mulAddRecFNToRaw_postMul_io_rawOut_sExp; // @[FMUL_1.scala 116:15]
  wire [26:0] mulAddRecFNToRaw_postMul_io_rawOut_sig; // @[FMUL_1.scala 116:15]
  wire  roundRawFNToRecFN_io_invalidExc; // @[FMUL_1.scala 137:15]
  wire  roundRawFNToRecFN_io_in_isNaN; // @[FMUL_1.scala 137:15]
  wire  roundRawFNToRecFN_io_in_isInf; // @[FMUL_1.scala 137:15]
  wire  roundRawFNToRecFN_io_in_isZero; // @[FMUL_1.scala 137:15]
  wire  roundRawFNToRecFN_io_in_sign; // @[FMUL_1.scala 137:15]
  wire [9:0] roundRawFNToRecFN_io_in_sExp; // @[FMUL_1.scala 137:15]
  wire [26:0] roundRawFNToRecFN_io_in_sig; // @[FMUL_1.scala 137:15]
  wire [32:0] roundRawFNToRecFN_io_out; // @[FMUL_1.scala 137:15]
  reg [23:0] premul_a; // @[FMUL_1.scala 15:37]
  reg [23:0] premul_b; // @[FMUL_1.scala 16:37]
  reg [47:0] premul_c; // @[FMUL_1.scala 17:37]
  reg  isSigNaNAny; // @[FMUL_1.scala 18:33]
  reg  isNaNAOrB; // @[FMUL_1.scala 19:34]
  reg  isInfA; // @[FMUL_1.scala 20:43]
  reg  isZeroA; // @[FMUL_1.scala 21:40]
  reg  isInfB; // @[FMUL_1.scala 22:43]
  reg  isZeroB; // @[FMUL_1.scala 23:40]
  reg  signProd; // @[FMUL_1.scala 24:38]
  reg  isNaNC; // @[FMUL_1.scala 25:39]
  reg  isInfC; // @[FMUL_1.scala 26:42]
  reg  isZeroC; // @[FMUL_1.scala 27:39]
  reg [9:0] sExpSum; // @[FMUL_1.scala 28:36]
  reg  doSubMags; // @[FMUL_1.scala 29:33]
  reg  CIsDominant; // @[FMUL_1.scala 30:33]
  reg [4:0] CDom_CAlignDist; // @[FMUL_1.scala 31:34]
  reg [25:0] highAlignedSigC; // @[FMUL_1.scala 32:37]
  reg  bit0AlignedSigC; // @[FMUL_1.scala 33:38]
  wire  _T_3 = io_a[30:23] == 8'h0; // @[rawFloatFromFN.scala 50:34]
  wire  _T_4 = io_a[22:0] == 23'h0; // @[rawFloatFromFN.scala 51:38]
  wire [4:0] _T_28 = io_a[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:69]
  wire [4:0] _T_29 = io_a[2] ? 5'h14 : _T_28; // @[Mux.scala 47:69]
  wire [4:0] _T_30 = io_a[3] ? 5'h13 : _T_29; // @[Mux.scala 47:69]
  wire [4:0] _T_31 = io_a[4] ? 5'h12 : _T_30; // @[Mux.scala 47:69]
  wire [4:0] _T_32 = io_a[5] ? 5'h11 : _T_31; // @[Mux.scala 47:69]
  wire [4:0] _T_33 = io_a[6] ? 5'h10 : _T_32; // @[Mux.scala 47:69]
  wire [4:0] _T_34 = io_a[7] ? 5'hf : _T_33; // @[Mux.scala 47:69]
  wire [4:0] _T_35 = io_a[8] ? 5'he : _T_34; // @[Mux.scala 47:69]
  wire [4:0] _T_36 = io_a[9] ? 5'hd : _T_35; // @[Mux.scala 47:69]
  wire [4:0] _T_37 = io_a[10] ? 5'hc : _T_36; // @[Mux.scala 47:69]
  wire [4:0] _T_38 = io_a[11] ? 5'hb : _T_37; // @[Mux.scala 47:69]
  wire [4:0] _T_39 = io_a[12] ? 5'ha : _T_38; // @[Mux.scala 47:69]
  wire [4:0] _T_40 = io_a[13] ? 5'h9 : _T_39; // @[Mux.scala 47:69]
  wire [4:0] _T_41 = io_a[14] ? 5'h8 : _T_40; // @[Mux.scala 47:69]
  wire [4:0] _T_42 = io_a[15] ? 5'h7 : _T_41; // @[Mux.scala 47:69]
  wire [4:0] _T_43 = io_a[16] ? 5'h6 : _T_42; // @[Mux.scala 47:69]
  wire [4:0] _T_44 = io_a[17] ? 5'h5 : _T_43; // @[Mux.scala 47:69]
  wire [4:0] _T_45 = io_a[18] ? 5'h4 : _T_44; // @[Mux.scala 47:69]
  wire [4:0] _T_46 = io_a[19] ? 5'h3 : _T_45; // @[Mux.scala 47:69]
  wire [4:0] _T_47 = io_a[20] ? 5'h2 : _T_46; // @[Mux.scala 47:69]
  wire [4:0] _T_48 = io_a[21] ? 5'h1 : _T_47; // @[Mux.scala 47:69]
  wire [4:0] _T_49 = io_a[22] ? 5'h0 : _T_48; // @[Mux.scala 47:69]
  wire [53:0] _GEN_0 = {{31'd0}, io_a[22:0]}; // @[rawFloatFromFN.scala 54:36]
  wire [53:0] _T_50 = _GEN_0 << _T_49; // @[rawFloatFromFN.scala 54:36]
  wire [22:0] _T_52 = {_T_50[21:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  wire [8:0] _GEN_1 = {{4'd0}, _T_49}; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_53 = _GEN_1 ^ 9'h1ff; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_54 = _T_3 ? _T_53 : {{1'd0}, io_a[30:23]}; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_55 = _T_3 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  wire [7:0] _GEN_2 = {{6'd0}, _T_55}; // @[rawFloatFromFN.scala 60:22]
  wire [7:0] _T_56 = 8'h80 | _GEN_2; // @[rawFloatFromFN.scala 60:22]
  wire [8:0] _GEN_3 = {{1'd0}, _T_56}; // @[rawFloatFromFN.scala 59:15]
  wire [8:0] _T_58 = _T_54 + _GEN_3; // @[rawFloatFromFN.scala 59:15]
  wire  _T_59 = _T_3 & _T_4; // @[rawFloatFromFN.scala 62:34]
  wire  _T_61 = _T_58[8:7] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  wire  _T_63 = _T_61 & ~_T_4; // @[rawFloatFromFN.scala 66:33]
  wire [9:0] _T_66 = {1'b0,$signed(_T_58)}; // @[rawFloatFromFN.scala 70:48]
  wire  hi_lo = ~_T_59; // @[rawFloatFromFN.scala 72:29]
  wire [22:0] lo = _T_3 ? _T_52 : io_a[22:0]; // @[rawFloatFromFN.scala 72:42]
  wire [24:0] _T_67 = {1'h0,hi_lo,lo}; // @[Cat.scala 30:58]
  wire [2:0] _T_69 = _T_59 ? 3'h0 : _T_66[8:6]; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_4 = {{2'd0}, _T_63}; // @[recFNFromFN.scala 48:79]
  wire [2:0] hi_lo_1 = _T_69 | _GEN_4; // @[recFNFromFN.scala 48:79]
  wire [5:0] lo_hi = _T_66[5:0]; // @[recFNFromFN.scala 50:23]
  wire [22:0] lo_lo = _T_67[22:0]; // @[recFNFromFN.scala 51:22]
  wire [28:0] lo_1 = {lo_hi,lo_lo}; // @[Cat.scala 30:58]
  wire [3:0] hi_1 = {io_a[31],hi_lo_1}; // @[Cat.scala 30:58]
  wire  _T_75 = io_b[30:23] == 8'h0; // @[rawFloatFromFN.scala 50:34]
  wire  _T_76 = io_b[22:0] == 23'h0; // @[rawFloatFromFN.scala 51:38]
  wire [4:0] _T_100 = io_b[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:69]
  wire [4:0] _T_101 = io_b[2] ? 5'h14 : _T_100; // @[Mux.scala 47:69]
  wire [4:0] _T_102 = io_b[3] ? 5'h13 : _T_101; // @[Mux.scala 47:69]
  wire [4:0] _T_103 = io_b[4] ? 5'h12 : _T_102; // @[Mux.scala 47:69]
  wire [4:0] _T_104 = io_b[5] ? 5'h11 : _T_103; // @[Mux.scala 47:69]
  wire [4:0] _T_105 = io_b[6] ? 5'h10 : _T_104; // @[Mux.scala 47:69]
  wire [4:0] _T_106 = io_b[7] ? 5'hf : _T_105; // @[Mux.scala 47:69]
  wire [4:0] _T_107 = io_b[8] ? 5'he : _T_106; // @[Mux.scala 47:69]
  wire [4:0] _T_108 = io_b[9] ? 5'hd : _T_107; // @[Mux.scala 47:69]
  wire [4:0] _T_109 = io_b[10] ? 5'hc : _T_108; // @[Mux.scala 47:69]
  wire [4:0] _T_110 = io_b[11] ? 5'hb : _T_109; // @[Mux.scala 47:69]
  wire [4:0] _T_111 = io_b[12] ? 5'ha : _T_110; // @[Mux.scala 47:69]
  wire [4:0] _T_112 = io_b[13] ? 5'h9 : _T_111; // @[Mux.scala 47:69]
  wire [4:0] _T_113 = io_b[14] ? 5'h8 : _T_112; // @[Mux.scala 47:69]
  wire [4:0] _T_114 = io_b[15] ? 5'h7 : _T_113; // @[Mux.scala 47:69]
  wire [4:0] _T_115 = io_b[16] ? 5'h6 : _T_114; // @[Mux.scala 47:69]
  wire [4:0] _T_116 = io_b[17] ? 5'h5 : _T_115; // @[Mux.scala 47:69]
  wire [4:0] _T_117 = io_b[18] ? 5'h4 : _T_116; // @[Mux.scala 47:69]
  wire [4:0] _T_118 = io_b[19] ? 5'h3 : _T_117; // @[Mux.scala 47:69]
  wire [4:0] _T_119 = io_b[20] ? 5'h2 : _T_118; // @[Mux.scala 47:69]
  wire [4:0] _T_120 = io_b[21] ? 5'h1 : _T_119; // @[Mux.scala 47:69]
  wire [4:0] _T_121 = io_b[22] ? 5'h0 : _T_120; // @[Mux.scala 47:69]
  wire [53:0] _GEN_5 = {{31'd0}, io_b[22:0]}; // @[rawFloatFromFN.scala 54:36]
  wire [53:0] _T_122 = _GEN_5 << _T_121; // @[rawFloatFromFN.scala 54:36]
  wire [22:0] _T_124 = {_T_122[21:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  wire [8:0] _GEN_6 = {{4'd0}, _T_121}; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_125 = _GEN_6 ^ 9'h1ff; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_126 = _T_75 ? _T_125 : {{1'd0}, io_b[30:23]}; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_127 = _T_75 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  wire [7:0] _GEN_7 = {{6'd0}, _T_127}; // @[rawFloatFromFN.scala 60:22]
  wire [7:0] _T_128 = 8'h80 | _GEN_7; // @[rawFloatFromFN.scala 60:22]
  wire [8:0] _GEN_8 = {{1'd0}, _T_128}; // @[rawFloatFromFN.scala 59:15]
  wire [8:0] _T_130 = _T_126 + _GEN_8; // @[rawFloatFromFN.scala 59:15]
  wire  _T_131 = _T_75 & _T_76; // @[rawFloatFromFN.scala 62:34]
  wire  _T_133 = _T_130[8:7] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  wire  _T_135 = _T_133 & ~_T_76; // @[rawFloatFromFN.scala 66:33]
  wire [9:0] _T_138 = {1'b0,$signed(_T_130)}; // @[rawFloatFromFN.scala 70:48]
  wire  hi_lo_2 = ~_T_131; // @[rawFloatFromFN.scala 72:29]
  wire [22:0] lo_2 = _T_75 ? _T_124 : io_b[22:0]; // @[rawFloatFromFN.scala 72:42]
  wire [24:0] _T_139 = {1'h0,hi_lo_2,lo_2}; // @[Cat.scala 30:58]
  wire [2:0] _T_141 = _T_131 ? 3'h0 : _T_138[8:6]; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_9 = {{2'd0}, _T_135}; // @[recFNFromFN.scala 48:79]
  wire [2:0] hi_lo_3 = _T_141 | _GEN_9; // @[recFNFromFN.scala 48:79]
  wire [5:0] lo_hi_1 = _T_138[5:0]; // @[recFNFromFN.scala 50:23]
  wire [22:0] lo_lo_1 = _T_139[22:0]; // @[recFNFromFN.scala 51:22]
  wire [28:0] lo_3 = {lo_hi_1,lo_lo_1}; // @[Cat.scala 30:58]
  wire [3:0] hi_3 = {io_b[31],hi_lo_3}; // @[Cat.scala 30:58]
  wire [31:0] _T_144 = io_a ^ io_b; // @[FMUL_1.scala 41:45]
  wire [31:0] _T_145 = _T_144 & 32'h80000000; // @[FMUL_1.scala 41:53]
  wire [47:0] _T_147 = premul_a * premul_b; // @[FMUL_1.scala 113:19]
  wire  _T_150 = roundRawFNToRecFN_io_out[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_152 = roundRawFNToRecFN_io_out[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  wire  _T_154 = _T_152 & roundRawFNToRecFN_io_out[29]; // @[rawFloatFromRecFN.scala 55:33]
  wire  _T_157 = _T_152 & ~roundRawFNToRecFN_io_out[29]; // @[rawFloatFromRecFN.scala 56:33]
  wire [9:0] _T_159 = {1'b0,$signed(roundRawFNToRecFN_io_out[31:23])}; // @[rawFloatFromRecFN.scala 59:27]
  wire  hi_lo_4 = ~_T_150; // @[rawFloatFromRecFN.scala 60:39]
  wire [22:0] lo_4 = roundRawFNToRecFN_io_out[22:0]; // @[rawFloatFromRecFN.scala 60:51]
  wire [24:0] _T_160 = {1'h0,hi_lo_4,lo_4}; // @[Cat.scala 30:58]
  wire  _T_161 = $signed(_T_159) < 10'sh82; // @[fNFromRecFN.scala 50:39]
  wire [4:0] _T_164 = 5'h1 - _T_159[4:0]; // @[fNFromRecFN.scala 51:39]
  wire [23:0] _T_166 = _T_160[24:1] >> _T_164; // @[fNFromRecFN.scala 52:42]
  wire [7:0] _T_170 = _T_159[7:0] - 8'h81; // @[fNFromRecFN.scala 57:45]
  wire [7:0] _T_171 = _T_161 ? 8'h0 : _T_170; // @[fNFromRecFN.scala 55:16]
  wire  _T_172 = _T_154 | _T_157; // @[fNFromRecFN.scala 59:44]
  wire [7:0] _T_174 = _T_172 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] hi_lo_5 = _T_171 | _T_174; // @[fNFromRecFN.scala 59:15]
  wire [22:0] _T_176 = _T_157 ? 23'h0 : _T_160[22:0]; // @[fNFromRecFN.scala 63:20]
  wire [22:0] lo_5 = _T_161 ? _T_166[22:0] : _T_176; // @[fNFromRecFN.scala 61:16]
  wire [8:0] hi_5 = {roundRawFNToRecFN_io_out[32],hi_lo_5}; // @[Cat.scala 30:58]
  MulAddRecFNToRaw_preMul mulAddRecFNToRaw_preMul ( // @[FMUL_1.scala 36:15]
    .io_a(mulAddRecFNToRaw_preMul_io_a),
    .io_b(mulAddRecFNToRaw_preMul_io_b),
    .io_c(mulAddRecFNToRaw_preMul_io_c),
    .io_mulAddA(mulAddRecFNToRaw_preMul_io_mulAddA),
    .io_mulAddB(mulAddRecFNToRaw_preMul_io_mulAddB),
    .io_mulAddC(mulAddRecFNToRaw_preMul_io_mulAddC),
    .io_toPostMul_isSigNaNAny(mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny),
    .io_toPostMul_isNaNAOrB(mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB),
    .io_toPostMul_isInfA(mulAddRecFNToRaw_preMul_io_toPostMul_isInfA),
    .io_toPostMul_isZeroA(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA),
    .io_toPostMul_isInfB(mulAddRecFNToRaw_preMul_io_toPostMul_isInfB),
    .io_toPostMul_isZeroB(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB),
    .io_toPostMul_signProd(mulAddRecFNToRaw_preMul_io_toPostMul_signProd),
    .io_toPostMul_isNaNC(mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC),
    .io_toPostMul_isInfC(mulAddRecFNToRaw_preMul_io_toPostMul_isInfC),
    .io_toPostMul_isZeroC(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC),
    .io_toPostMul_sExpSum(mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum),
    .io_toPostMul_doSubMags(mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags),
    .io_toPostMul_CIsDominant(mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant),
    .io_toPostMul_CDom_CAlignDist(mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist),
    .io_toPostMul_highAlignedSigC(mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC),
    .io_toPostMul_bit0AlignedSigC(mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC)
  );
  MulAddRecFNToRaw_postMul mulAddRecFNToRaw_postMul ( // @[FMUL_1.scala 116:15]
    .io_fromPreMul_isSigNaNAny(mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny),
    .io_fromPreMul_isNaNAOrB(mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB),
    .io_fromPreMul_isInfA(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA),
    .io_fromPreMul_isZeroA(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA),
    .io_fromPreMul_isInfB(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB),
    .io_fromPreMul_isZeroB(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB),
    .io_fromPreMul_signProd(mulAddRecFNToRaw_postMul_io_fromPreMul_signProd),
    .io_fromPreMul_isNaNC(mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC),
    .io_fromPreMul_isInfC(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC),
    .io_fromPreMul_isZeroC(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC),
    .io_fromPreMul_sExpSum(mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum),
    .io_fromPreMul_doSubMags(mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags),
    .io_fromPreMul_CIsDominant(mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant),
    .io_fromPreMul_CDom_CAlignDist(mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist),
    .io_fromPreMul_highAlignedSigC(mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC),
    .io_fromPreMul_bit0AlignedSigC(mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC),
    .io_mulAddResult(mulAddRecFNToRaw_postMul_io_mulAddResult),
    .io_invalidExc(mulAddRecFNToRaw_postMul_io_invalidExc),
    .io_rawOut_isNaN(mulAddRecFNToRaw_postMul_io_rawOut_isNaN),
    .io_rawOut_isInf(mulAddRecFNToRaw_postMul_io_rawOut_isInf),
    .io_rawOut_isZero(mulAddRecFNToRaw_postMul_io_rawOut_isZero),
    .io_rawOut_sign(mulAddRecFNToRaw_postMul_io_rawOut_sign),
    .io_rawOut_sExp(mulAddRecFNToRaw_postMul_io_rawOut_sExp),
    .io_rawOut_sig(mulAddRecFNToRaw_postMul_io_rawOut_sig)
  );
  RoundRawFNToRecFN roundRawFNToRecFN ( // @[FMUL_1.scala 137:15]
    .io_invalidExc(roundRawFNToRecFN_io_invalidExc),
    .io_in_isNaN(roundRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundRawFNToRecFN_io_in_sig),
    .io_out(roundRawFNToRecFN_io_out)
  );
  assign io_out = {hi_5,lo_5}; // @[Cat.scala 30:58]
  assign mulAddRecFNToRaw_preMul_io_a = {hi_1,lo_1}; // @[Cat.scala 30:58]
  assign mulAddRecFNToRaw_preMul_io_b = {hi_3,lo_3}; // @[Cat.scala 30:58]
  assign mulAddRecFNToRaw_preMul_io_c = {_T_145, 1'h0}; // @[FMUL_1.scala 41:75]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny = isSigNaNAny; // @[FMUL_1.scala 119:84]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB = isNaNAOrB; // @[FMUL_1.scala 120:86]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA = isInfA; // @[FMUL_1.scala 121:94]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA = isZeroA; // @[FMUL_1.scala 122:91]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB = isInfB; // @[FMUL_1.scala 123:94]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB = isZeroB; // @[FMUL_1.scala 124:91]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_signProd = signProd; // @[FMUL_1.scala 125:89]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC = isNaNC; // @[FMUL_1.scala 126:90]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC = isInfC; // @[FMUL_1.scala 127:94]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC = isZeroC; // @[FMUL_1.scala 128:91]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum = sExpSum; // @[FMUL_1.scala 129:88]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags = doSubMags; // @[FMUL_1.scala 130:85]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant = CIsDominant; // @[FMUL_1.scala 131:84]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist = CDom_CAlignDist; // @[FMUL_1.scala 132:78]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC = highAlignedSigC; // @[FMUL_1.scala 133:80]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC = bit0AlignedSigC; // @[FMUL_1.scala 134:82]
  assign mulAddRecFNToRaw_postMul_io_mulAddResult = _T_147 + premul_c; // @[FMUL_1.scala 113:31]
  assign roundRawFNToRecFN_io_invalidExc = mulAddRecFNToRaw_postMul_io_invalidExc; // @[FMUL_1.scala 138:39]
  assign roundRawFNToRecFN_io_in_isNaN = mulAddRecFNToRaw_postMul_io_rawOut_isNaN; // @[FMUL_1.scala 140:39]
  assign roundRawFNToRecFN_io_in_isInf = mulAddRecFNToRaw_postMul_io_rawOut_isInf; // @[FMUL_1.scala 140:39]
  assign roundRawFNToRecFN_io_in_isZero = mulAddRecFNToRaw_postMul_io_rawOut_isZero; // @[FMUL_1.scala 140:39]
  assign roundRawFNToRecFN_io_in_sign = mulAddRecFNToRaw_postMul_io_rawOut_sign; // @[FMUL_1.scala 140:39]
  assign roundRawFNToRecFN_io_in_sExp = mulAddRecFNToRaw_postMul_io_rawOut_sExp; // @[FMUL_1.scala 140:39]
  assign roundRawFNToRecFN_io_in_sig = mulAddRecFNToRaw_postMul_io_rawOut_sig; // @[FMUL_1.scala 140:39]
  always @(posedge clock) begin
    if (reset) begin // @[FMUL_1.scala 15:37]
      premul_a <= 24'h0; // @[FMUL_1.scala 15:37]
    end else begin
      premul_a <= mulAddRecFNToRaw_preMul_io_mulAddA; // @[FMUL_1.scala 103:63]
    end
    if (reset) begin // @[FMUL_1.scala 16:37]
      premul_b <= 24'h0; // @[FMUL_1.scala 16:37]
    end else begin
      premul_b <= mulAddRecFNToRaw_preMul_io_mulAddB; // @[FMUL_1.scala 104:63]
    end
    if (reset) begin // @[FMUL_1.scala 17:37]
      premul_c <= 48'h0; // @[FMUL_1.scala 17:37]
    end else begin
      premul_c <= mulAddRecFNToRaw_preMul_io_mulAddC; // @[FMUL_1.scala 105:63]
    end
    if (reset) begin // @[FMUL_1.scala 18:33]
      isSigNaNAny <= 1'h0; // @[FMUL_1.scala 18:33]
    end else begin
      isSigNaNAny <= mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny; // @[FMUL_1.scala 43:61]
    end
    if (reset) begin // @[FMUL_1.scala 19:34]
      isNaNAOrB <= 1'h0; // @[FMUL_1.scala 19:34]
    end else begin
      isNaNAOrB <= mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB; // @[FMUL_1.scala 44:62]
    end
    if (reset) begin // @[FMUL_1.scala 20:43]
      isInfA <= 1'h0; // @[FMUL_1.scala 20:43]
    end else begin
      isInfA <= mulAddRecFNToRaw_preMul_io_toPostMul_isInfA; // @[FMUL_1.scala 45:70]
    end
    if (reset) begin // @[FMUL_1.scala 21:40]
      isZeroA <= 1'h0; // @[FMUL_1.scala 21:40]
    end else begin
      isZeroA <= mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA; // @[FMUL_1.scala 46:67]
    end
    if (reset) begin // @[FMUL_1.scala 22:43]
      isInfB <= 1'h0; // @[FMUL_1.scala 22:43]
    end else begin
      isInfB <= mulAddRecFNToRaw_preMul_io_toPostMul_isInfB; // @[FMUL_1.scala 47:70]
    end
    if (reset) begin // @[FMUL_1.scala 23:40]
      isZeroB <= 1'h0; // @[FMUL_1.scala 23:40]
    end else begin
      isZeroB <= mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB; // @[FMUL_1.scala 48:67]
    end
    if (reset) begin // @[FMUL_1.scala 24:38]
      signProd <= 1'h0; // @[FMUL_1.scala 24:38]
    end else begin
      signProd <= mulAddRecFNToRaw_preMul_io_toPostMul_signProd; // @[FMUL_1.scala 49:65]
    end
    if (reset) begin // @[FMUL_1.scala 25:39]
      isNaNC <= 1'h0; // @[FMUL_1.scala 25:39]
    end else begin
      isNaNC <= mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC; // @[FMUL_1.scala 50:66]
    end
    if (reset) begin // @[FMUL_1.scala 26:42]
      isInfC <= 1'h0; // @[FMUL_1.scala 26:42]
    end else begin
      isInfC <= mulAddRecFNToRaw_preMul_io_toPostMul_isInfC; // @[FMUL_1.scala 51:69]
    end
    if (reset) begin // @[FMUL_1.scala 27:39]
      isZeroC <= 1'h0; // @[FMUL_1.scala 27:39]
    end else begin
      isZeroC <= mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC; // @[FMUL_1.scala 52:66]
    end
    if (reset) begin // @[FMUL_1.scala 28:36]
      sExpSum <= 10'sh0; // @[FMUL_1.scala 28:36]
    end else begin
      sExpSum <= mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum; // @[FMUL_1.scala 53:63]
    end
    if (reset) begin // @[FMUL_1.scala 29:33]
      doSubMags <= 1'h0; // @[FMUL_1.scala 29:33]
    end else begin
      doSubMags <= mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags; // @[FMUL_1.scala 54:60]
    end
    if (reset) begin // @[FMUL_1.scala 30:33]
      CIsDominant <= 1'h0; // @[FMUL_1.scala 30:33]
    end else begin
      CIsDominant <= mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant; // @[FMUL_1.scala 55:59]
    end
    if (reset) begin // @[FMUL_1.scala 31:34]
      CDom_CAlignDist <= 5'h0; // @[FMUL_1.scala 31:34]
    end else begin
      CDom_CAlignDist <= mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist; // @[FMUL_1.scala 56:54]
    end
    if (reset) begin // @[FMUL_1.scala 32:37]
      highAlignedSigC <= 26'h0; // @[FMUL_1.scala 32:37]
    end else begin
      highAlignedSigC <= mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC; // @[FMUL_1.scala 57:56]
    end
    if (reset) begin // @[FMUL_1.scala 33:38]
      bit0AlignedSigC <= 1'h0; // @[FMUL_1.scala 33:38]
    end else begin
      bit0AlignedSigC <= mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC; // @[FMUL_1.scala 58:57]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  premul_a = _RAND_0[23:0];
  _RAND_1 = {1{`RANDOM}};
  premul_b = _RAND_1[23:0];
  _RAND_2 = {2{`RANDOM}};
  premul_c = _RAND_2[47:0];
  _RAND_3 = {1{`RANDOM}};
  isSigNaNAny = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  isNaNAOrB = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  isInfA = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  isZeroA = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  isInfB = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  isZeroB = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  signProd = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  isNaNC = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  isInfC = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  isZeroC = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  sExpSum = _RAND_13[9:0];
  _RAND_14 = {1{`RANDOM}};
  doSubMags = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  CIsDominant = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  CDom_CAlignDist = _RAND_16[4:0];
  _RAND_17 = {1{`RANDOM}};
  highAlignedSigC = _RAND_17[25:0];
  _RAND_18 = {1{`RANDOM}};
  bit0AlignedSigC = _RAND_18[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MY_ADD(
  input         clock,
  input         reset,
  input  [31:0] io_a,
  input  [31:0] io_b,
  output [31:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_REG_INIT
  wire [32:0] mulAddRecFNToRaw_preMul_io_a; // @[FADD_1.scala 36:15]
  wire [32:0] mulAddRecFNToRaw_preMul_io_b; // @[FADD_1.scala 36:15]
  wire [32:0] mulAddRecFNToRaw_preMul_io_c; // @[FADD_1.scala 36:15]
  wire [23:0] mulAddRecFNToRaw_preMul_io_mulAddA; // @[FADD_1.scala 36:15]
  wire [23:0] mulAddRecFNToRaw_preMul_io_mulAddB; // @[FADD_1.scala 36:15]
  wire [47:0] mulAddRecFNToRaw_preMul_io_mulAddC; // @[FADD_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny; // @[FADD_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB; // @[FADD_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfA; // @[FADD_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA; // @[FADD_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfB; // @[FADD_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB; // @[FADD_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_signProd; // @[FADD_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC; // @[FADD_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfC; // @[FADD_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC; // @[FADD_1.scala 36:15]
  wire [9:0] mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum; // @[FADD_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags; // @[FADD_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant; // @[FADD_1.scala 36:15]
  wire [4:0] mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist; // @[FADD_1.scala 36:15]
  wire [25:0] mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC; // @[FADD_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC; // @[FADD_1.scala 36:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny; // @[FADD_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB; // @[FADD_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA; // @[FADD_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA; // @[FADD_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB; // @[FADD_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB; // @[FADD_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_signProd; // @[FADD_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC; // @[FADD_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC; // @[FADD_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC; // @[FADD_1.scala 116:15]
  wire [9:0] mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum; // @[FADD_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags; // @[FADD_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant; // @[FADD_1.scala 116:15]
  wire [4:0] mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist; // @[FADD_1.scala 116:15]
  wire [25:0] mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC; // @[FADD_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC; // @[FADD_1.scala 116:15]
  wire [48:0] mulAddRecFNToRaw_postMul_io_mulAddResult; // @[FADD_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_invalidExc; // @[FADD_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isNaN; // @[FADD_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isInf; // @[FADD_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isZero; // @[FADD_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_sign; // @[FADD_1.scala 116:15]
  wire [9:0] mulAddRecFNToRaw_postMul_io_rawOut_sExp; // @[FADD_1.scala 116:15]
  wire [26:0] mulAddRecFNToRaw_postMul_io_rawOut_sig; // @[FADD_1.scala 116:15]
  wire  roundRawFNToRecFN_io_invalidExc; // @[FADD_1.scala 137:15]
  wire  roundRawFNToRecFN_io_in_isNaN; // @[FADD_1.scala 137:15]
  wire  roundRawFNToRecFN_io_in_isInf; // @[FADD_1.scala 137:15]
  wire  roundRawFNToRecFN_io_in_isZero; // @[FADD_1.scala 137:15]
  wire  roundRawFNToRecFN_io_in_sign; // @[FADD_1.scala 137:15]
  wire [9:0] roundRawFNToRecFN_io_in_sExp; // @[FADD_1.scala 137:15]
  wire [26:0] roundRawFNToRecFN_io_in_sig; // @[FADD_1.scala 137:15]
  wire [32:0] roundRawFNToRecFN_io_out; // @[FADD_1.scala 137:15]
  reg [23:0] premul_a; // @[FADD_1.scala 15:37]
  reg [23:0] premul_b; // @[FADD_1.scala 16:37]
  reg [47:0] premul_c; // @[FADD_1.scala 17:37]
  reg  isSigNaNAny; // @[FADD_1.scala 18:33]
  reg  isNaNAOrB; // @[FADD_1.scala 19:34]
  reg  isInfA; // @[FADD_1.scala 20:43]
  reg  isZeroA; // @[FADD_1.scala 21:40]
  reg  isInfB; // @[FADD_1.scala 22:43]
  reg  isZeroB; // @[FADD_1.scala 23:40]
  reg  signProd; // @[FADD_1.scala 24:38]
  reg  isNaNC; // @[FADD_1.scala 25:39]
  reg  isInfC; // @[FADD_1.scala 26:42]
  reg  isZeroC; // @[FADD_1.scala 27:39]
  reg [9:0] sExpSum; // @[FADD_1.scala 28:36]
  reg  doSubMags; // @[FADD_1.scala 29:33]
  reg  CIsDominant; // @[FADD_1.scala 30:33]
  reg [4:0] CDom_CAlignDist; // @[FADD_1.scala 31:34]
  reg [25:0] highAlignedSigC; // @[FADD_1.scala 32:37]
  reg  bit0AlignedSigC; // @[FADD_1.scala 33:38]
  wire  _T_3 = io_a[30:23] == 8'h0; // @[rawFloatFromFN.scala 50:34]
  wire  _T_4 = io_a[22:0] == 23'h0; // @[rawFloatFromFN.scala 51:38]
  wire [4:0] _T_28 = io_a[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:69]
  wire [4:0] _T_29 = io_a[2] ? 5'h14 : _T_28; // @[Mux.scala 47:69]
  wire [4:0] _T_30 = io_a[3] ? 5'h13 : _T_29; // @[Mux.scala 47:69]
  wire [4:0] _T_31 = io_a[4] ? 5'h12 : _T_30; // @[Mux.scala 47:69]
  wire [4:0] _T_32 = io_a[5] ? 5'h11 : _T_31; // @[Mux.scala 47:69]
  wire [4:0] _T_33 = io_a[6] ? 5'h10 : _T_32; // @[Mux.scala 47:69]
  wire [4:0] _T_34 = io_a[7] ? 5'hf : _T_33; // @[Mux.scala 47:69]
  wire [4:0] _T_35 = io_a[8] ? 5'he : _T_34; // @[Mux.scala 47:69]
  wire [4:0] _T_36 = io_a[9] ? 5'hd : _T_35; // @[Mux.scala 47:69]
  wire [4:0] _T_37 = io_a[10] ? 5'hc : _T_36; // @[Mux.scala 47:69]
  wire [4:0] _T_38 = io_a[11] ? 5'hb : _T_37; // @[Mux.scala 47:69]
  wire [4:0] _T_39 = io_a[12] ? 5'ha : _T_38; // @[Mux.scala 47:69]
  wire [4:0] _T_40 = io_a[13] ? 5'h9 : _T_39; // @[Mux.scala 47:69]
  wire [4:0] _T_41 = io_a[14] ? 5'h8 : _T_40; // @[Mux.scala 47:69]
  wire [4:0] _T_42 = io_a[15] ? 5'h7 : _T_41; // @[Mux.scala 47:69]
  wire [4:0] _T_43 = io_a[16] ? 5'h6 : _T_42; // @[Mux.scala 47:69]
  wire [4:0] _T_44 = io_a[17] ? 5'h5 : _T_43; // @[Mux.scala 47:69]
  wire [4:0] _T_45 = io_a[18] ? 5'h4 : _T_44; // @[Mux.scala 47:69]
  wire [4:0] _T_46 = io_a[19] ? 5'h3 : _T_45; // @[Mux.scala 47:69]
  wire [4:0] _T_47 = io_a[20] ? 5'h2 : _T_46; // @[Mux.scala 47:69]
  wire [4:0] _T_48 = io_a[21] ? 5'h1 : _T_47; // @[Mux.scala 47:69]
  wire [4:0] _T_49 = io_a[22] ? 5'h0 : _T_48; // @[Mux.scala 47:69]
  wire [53:0] _GEN_0 = {{31'd0}, io_a[22:0]}; // @[rawFloatFromFN.scala 54:36]
  wire [53:0] _T_50 = _GEN_0 << _T_49; // @[rawFloatFromFN.scala 54:36]
  wire [22:0] _T_52 = {_T_50[21:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  wire [8:0] _GEN_1 = {{4'd0}, _T_49}; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_53 = _GEN_1 ^ 9'h1ff; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_54 = _T_3 ? _T_53 : {{1'd0}, io_a[30:23]}; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_55 = _T_3 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  wire [7:0] _GEN_2 = {{6'd0}, _T_55}; // @[rawFloatFromFN.scala 60:22]
  wire [7:0] _T_56 = 8'h80 | _GEN_2; // @[rawFloatFromFN.scala 60:22]
  wire [8:0] _GEN_3 = {{1'd0}, _T_56}; // @[rawFloatFromFN.scala 59:15]
  wire [8:0] _T_58 = _T_54 + _GEN_3; // @[rawFloatFromFN.scala 59:15]
  wire  _T_59 = _T_3 & _T_4; // @[rawFloatFromFN.scala 62:34]
  wire  _T_61 = _T_58[8:7] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  wire  _T_63 = _T_61 & ~_T_4; // @[rawFloatFromFN.scala 66:33]
  wire [9:0] _T_66 = {1'b0,$signed(_T_58)}; // @[rawFloatFromFN.scala 70:48]
  wire  hi_lo = ~_T_59; // @[rawFloatFromFN.scala 72:29]
  wire [22:0] lo = _T_3 ? _T_52 : io_a[22:0]; // @[rawFloatFromFN.scala 72:42]
  wire [24:0] _T_67 = {1'h0,hi_lo,lo}; // @[Cat.scala 30:58]
  wire [2:0] _T_69 = _T_59 ? 3'h0 : _T_66[8:6]; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_4 = {{2'd0}, _T_63}; // @[recFNFromFN.scala 48:79]
  wire [2:0] hi_lo_1 = _T_69 | _GEN_4; // @[recFNFromFN.scala 48:79]
  wire [5:0] lo_hi = _T_66[5:0]; // @[recFNFromFN.scala 50:23]
  wire [22:0] lo_lo = _T_67[22:0]; // @[recFNFromFN.scala 51:22]
  wire [28:0] lo_1 = {lo_hi,lo_lo}; // @[Cat.scala 30:58]
  wire [3:0] hi_1 = {io_a[31],hi_lo_1}; // @[Cat.scala 30:58]
  wire  _T_75 = io_b[30:23] == 8'h0; // @[rawFloatFromFN.scala 50:34]
  wire  _T_76 = io_b[22:0] == 23'h0; // @[rawFloatFromFN.scala 51:38]
  wire [4:0] _T_100 = io_b[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:69]
  wire [4:0] _T_101 = io_b[2] ? 5'h14 : _T_100; // @[Mux.scala 47:69]
  wire [4:0] _T_102 = io_b[3] ? 5'h13 : _T_101; // @[Mux.scala 47:69]
  wire [4:0] _T_103 = io_b[4] ? 5'h12 : _T_102; // @[Mux.scala 47:69]
  wire [4:0] _T_104 = io_b[5] ? 5'h11 : _T_103; // @[Mux.scala 47:69]
  wire [4:0] _T_105 = io_b[6] ? 5'h10 : _T_104; // @[Mux.scala 47:69]
  wire [4:0] _T_106 = io_b[7] ? 5'hf : _T_105; // @[Mux.scala 47:69]
  wire [4:0] _T_107 = io_b[8] ? 5'he : _T_106; // @[Mux.scala 47:69]
  wire [4:0] _T_108 = io_b[9] ? 5'hd : _T_107; // @[Mux.scala 47:69]
  wire [4:0] _T_109 = io_b[10] ? 5'hc : _T_108; // @[Mux.scala 47:69]
  wire [4:0] _T_110 = io_b[11] ? 5'hb : _T_109; // @[Mux.scala 47:69]
  wire [4:0] _T_111 = io_b[12] ? 5'ha : _T_110; // @[Mux.scala 47:69]
  wire [4:0] _T_112 = io_b[13] ? 5'h9 : _T_111; // @[Mux.scala 47:69]
  wire [4:0] _T_113 = io_b[14] ? 5'h8 : _T_112; // @[Mux.scala 47:69]
  wire [4:0] _T_114 = io_b[15] ? 5'h7 : _T_113; // @[Mux.scala 47:69]
  wire [4:0] _T_115 = io_b[16] ? 5'h6 : _T_114; // @[Mux.scala 47:69]
  wire [4:0] _T_116 = io_b[17] ? 5'h5 : _T_115; // @[Mux.scala 47:69]
  wire [4:0] _T_117 = io_b[18] ? 5'h4 : _T_116; // @[Mux.scala 47:69]
  wire [4:0] _T_118 = io_b[19] ? 5'h3 : _T_117; // @[Mux.scala 47:69]
  wire [4:0] _T_119 = io_b[20] ? 5'h2 : _T_118; // @[Mux.scala 47:69]
  wire [4:0] _T_120 = io_b[21] ? 5'h1 : _T_119; // @[Mux.scala 47:69]
  wire [4:0] _T_121 = io_b[22] ? 5'h0 : _T_120; // @[Mux.scala 47:69]
  wire [53:0] _GEN_5 = {{31'd0}, io_b[22:0]}; // @[rawFloatFromFN.scala 54:36]
  wire [53:0] _T_122 = _GEN_5 << _T_121; // @[rawFloatFromFN.scala 54:36]
  wire [22:0] _T_124 = {_T_122[21:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  wire [8:0] _GEN_6 = {{4'd0}, _T_121}; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_125 = _GEN_6 ^ 9'h1ff; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_126 = _T_75 ? _T_125 : {{1'd0}, io_b[30:23]}; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_127 = _T_75 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  wire [7:0] _GEN_7 = {{6'd0}, _T_127}; // @[rawFloatFromFN.scala 60:22]
  wire [7:0] _T_128 = 8'h80 | _GEN_7; // @[rawFloatFromFN.scala 60:22]
  wire [8:0] _GEN_8 = {{1'd0}, _T_128}; // @[rawFloatFromFN.scala 59:15]
  wire [8:0] _T_130 = _T_126 + _GEN_8; // @[rawFloatFromFN.scala 59:15]
  wire  _T_131 = _T_75 & _T_76; // @[rawFloatFromFN.scala 62:34]
  wire  _T_133 = _T_130[8:7] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  wire  _T_135 = _T_133 & ~_T_76; // @[rawFloatFromFN.scala 66:33]
  wire [9:0] _T_138 = {1'b0,$signed(_T_130)}; // @[rawFloatFromFN.scala 70:48]
  wire  hi_lo_2 = ~_T_131; // @[rawFloatFromFN.scala 72:29]
  wire [22:0] lo_2 = _T_75 ? _T_124 : io_b[22:0]; // @[rawFloatFromFN.scala 72:42]
  wire [24:0] _T_139 = {1'h0,hi_lo_2,lo_2}; // @[Cat.scala 30:58]
  wire [2:0] _T_141 = _T_131 ? 3'h0 : _T_138[8:6]; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_9 = {{2'd0}, _T_135}; // @[recFNFromFN.scala 48:79]
  wire [2:0] hi_lo_3 = _T_141 | _GEN_9; // @[recFNFromFN.scala 48:79]
  wire [5:0] lo_hi_1 = _T_138[5:0]; // @[recFNFromFN.scala 50:23]
  wire [22:0] lo_lo_1 = _T_139[22:0]; // @[recFNFromFN.scala 51:22]
  wire [28:0] lo_3 = {lo_hi_1,lo_lo_1}; // @[Cat.scala 30:58]
  wire [3:0] hi_3 = {io_b[31],hi_lo_3}; // @[Cat.scala 30:58]
  wire [47:0] _T_144 = premul_a * premul_b; // @[FADD_1.scala 113:19]
  wire  _T_147 = roundRawFNToRecFN_io_out[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_149 = roundRawFNToRecFN_io_out[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  wire  _T_151 = _T_149 & roundRawFNToRecFN_io_out[29]; // @[rawFloatFromRecFN.scala 55:33]
  wire  _T_154 = _T_149 & ~roundRawFNToRecFN_io_out[29]; // @[rawFloatFromRecFN.scala 56:33]
  wire [9:0] _T_156 = {1'b0,$signed(roundRawFNToRecFN_io_out[31:23])}; // @[rawFloatFromRecFN.scala 59:27]
  wire  hi_lo_4 = ~_T_147; // @[rawFloatFromRecFN.scala 60:39]
  wire [22:0] lo_4 = roundRawFNToRecFN_io_out[22:0]; // @[rawFloatFromRecFN.scala 60:51]
  wire [24:0] _T_157 = {1'h0,hi_lo_4,lo_4}; // @[Cat.scala 30:58]
  wire  _T_158 = $signed(_T_156) < 10'sh82; // @[fNFromRecFN.scala 50:39]
  wire [4:0] _T_161 = 5'h1 - _T_156[4:0]; // @[fNFromRecFN.scala 51:39]
  wire [23:0] _T_163 = _T_157[24:1] >> _T_161; // @[fNFromRecFN.scala 52:42]
  wire [7:0] _T_167 = _T_156[7:0] - 8'h81; // @[fNFromRecFN.scala 57:45]
  wire [7:0] _T_168 = _T_158 ? 8'h0 : _T_167; // @[fNFromRecFN.scala 55:16]
  wire  _T_169 = _T_151 | _T_154; // @[fNFromRecFN.scala 59:44]
  wire [7:0] _T_171 = _T_169 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] hi_lo_5 = _T_168 | _T_171; // @[fNFromRecFN.scala 59:15]
  wire [22:0] _T_173 = _T_154 ? 23'h0 : _T_157[22:0]; // @[fNFromRecFN.scala 63:20]
  wire [22:0] lo_5 = _T_158 ? _T_163[22:0] : _T_173; // @[fNFromRecFN.scala 61:16]
  wire [8:0] hi_5 = {roundRawFNToRecFN_io_out[32],hi_lo_5}; // @[Cat.scala 30:58]
  MulAddRecFNToRaw_preMul mulAddRecFNToRaw_preMul ( // @[FADD_1.scala 36:15]
    .io_a(mulAddRecFNToRaw_preMul_io_a),
    .io_b(mulAddRecFNToRaw_preMul_io_b),
    .io_c(mulAddRecFNToRaw_preMul_io_c),
    .io_mulAddA(mulAddRecFNToRaw_preMul_io_mulAddA),
    .io_mulAddB(mulAddRecFNToRaw_preMul_io_mulAddB),
    .io_mulAddC(mulAddRecFNToRaw_preMul_io_mulAddC),
    .io_toPostMul_isSigNaNAny(mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny),
    .io_toPostMul_isNaNAOrB(mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB),
    .io_toPostMul_isInfA(mulAddRecFNToRaw_preMul_io_toPostMul_isInfA),
    .io_toPostMul_isZeroA(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA),
    .io_toPostMul_isInfB(mulAddRecFNToRaw_preMul_io_toPostMul_isInfB),
    .io_toPostMul_isZeroB(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB),
    .io_toPostMul_signProd(mulAddRecFNToRaw_preMul_io_toPostMul_signProd),
    .io_toPostMul_isNaNC(mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC),
    .io_toPostMul_isInfC(mulAddRecFNToRaw_preMul_io_toPostMul_isInfC),
    .io_toPostMul_isZeroC(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC),
    .io_toPostMul_sExpSum(mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum),
    .io_toPostMul_doSubMags(mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags),
    .io_toPostMul_CIsDominant(mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant),
    .io_toPostMul_CDom_CAlignDist(mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist),
    .io_toPostMul_highAlignedSigC(mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC),
    .io_toPostMul_bit0AlignedSigC(mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC)
  );
  MulAddRecFNToRaw_postMul mulAddRecFNToRaw_postMul ( // @[FADD_1.scala 116:15]
    .io_fromPreMul_isSigNaNAny(mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny),
    .io_fromPreMul_isNaNAOrB(mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB),
    .io_fromPreMul_isInfA(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA),
    .io_fromPreMul_isZeroA(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA),
    .io_fromPreMul_isInfB(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB),
    .io_fromPreMul_isZeroB(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB),
    .io_fromPreMul_signProd(mulAddRecFNToRaw_postMul_io_fromPreMul_signProd),
    .io_fromPreMul_isNaNC(mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC),
    .io_fromPreMul_isInfC(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC),
    .io_fromPreMul_isZeroC(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC),
    .io_fromPreMul_sExpSum(mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum),
    .io_fromPreMul_doSubMags(mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags),
    .io_fromPreMul_CIsDominant(mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant),
    .io_fromPreMul_CDom_CAlignDist(mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist),
    .io_fromPreMul_highAlignedSigC(mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC),
    .io_fromPreMul_bit0AlignedSigC(mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC),
    .io_mulAddResult(mulAddRecFNToRaw_postMul_io_mulAddResult),
    .io_invalidExc(mulAddRecFNToRaw_postMul_io_invalidExc),
    .io_rawOut_isNaN(mulAddRecFNToRaw_postMul_io_rawOut_isNaN),
    .io_rawOut_isInf(mulAddRecFNToRaw_postMul_io_rawOut_isInf),
    .io_rawOut_isZero(mulAddRecFNToRaw_postMul_io_rawOut_isZero),
    .io_rawOut_sign(mulAddRecFNToRaw_postMul_io_rawOut_sign),
    .io_rawOut_sExp(mulAddRecFNToRaw_postMul_io_rawOut_sExp),
    .io_rawOut_sig(mulAddRecFNToRaw_postMul_io_rawOut_sig)
  );
  RoundRawFNToRecFN roundRawFNToRecFN ( // @[FADD_1.scala 137:15]
    .io_invalidExc(roundRawFNToRecFN_io_invalidExc),
    .io_in_isNaN(roundRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundRawFNToRecFN_io_in_sig),
    .io_out(roundRawFNToRecFN_io_out)
  );
  assign io_out = {hi_5,lo_5}; // @[Cat.scala 30:58]
  assign mulAddRecFNToRaw_preMul_io_a = {hi_1,lo_1}; // @[Cat.scala 30:58]
  assign mulAddRecFNToRaw_preMul_io_b = 33'h80000000; // @[FADD_1.scala 40:35]
  assign mulAddRecFNToRaw_preMul_io_c = {hi_3,lo_3}; // @[Cat.scala 30:58]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny = isSigNaNAny; // @[FADD_1.scala 119:84]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB = isNaNAOrB; // @[FADD_1.scala 120:86]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA = isInfA; // @[FADD_1.scala 121:94]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA = isZeroA; // @[FADD_1.scala 122:91]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB = isInfB; // @[FADD_1.scala 123:94]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB = isZeroB; // @[FADD_1.scala 124:91]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_signProd = signProd; // @[FADD_1.scala 125:89]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC = isNaNC; // @[FADD_1.scala 126:90]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC = isInfC; // @[FADD_1.scala 127:94]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC = isZeroC; // @[FADD_1.scala 128:91]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum = sExpSum; // @[FADD_1.scala 129:88]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags = doSubMags; // @[FADD_1.scala 130:85]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant = CIsDominant; // @[FADD_1.scala 131:84]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist = CDom_CAlignDist; // @[FADD_1.scala 132:78]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC = highAlignedSigC; // @[FADD_1.scala 133:80]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC = bit0AlignedSigC; // @[FADD_1.scala 134:82]
  assign mulAddRecFNToRaw_postMul_io_mulAddResult = _T_144 + premul_c; // @[FADD_1.scala 113:31]
  assign roundRawFNToRecFN_io_invalidExc = mulAddRecFNToRaw_postMul_io_invalidExc; // @[FADD_1.scala 138:39]
  assign roundRawFNToRecFN_io_in_isNaN = mulAddRecFNToRaw_postMul_io_rawOut_isNaN; // @[FADD_1.scala 140:39]
  assign roundRawFNToRecFN_io_in_isInf = mulAddRecFNToRaw_postMul_io_rawOut_isInf; // @[FADD_1.scala 140:39]
  assign roundRawFNToRecFN_io_in_isZero = mulAddRecFNToRaw_postMul_io_rawOut_isZero; // @[FADD_1.scala 140:39]
  assign roundRawFNToRecFN_io_in_sign = mulAddRecFNToRaw_postMul_io_rawOut_sign; // @[FADD_1.scala 140:39]
  assign roundRawFNToRecFN_io_in_sExp = mulAddRecFNToRaw_postMul_io_rawOut_sExp; // @[FADD_1.scala 140:39]
  assign roundRawFNToRecFN_io_in_sig = mulAddRecFNToRaw_postMul_io_rawOut_sig; // @[FADD_1.scala 140:39]
  always @(posedge clock) begin
    if (reset) begin // @[FADD_1.scala 15:37]
      premul_a <= 24'h0; // @[FADD_1.scala 15:37]
    end else begin
      premul_a <= mulAddRecFNToRaw_preMul_io_mulAddA; // @[FADD_1.scala 103:63]
    end
    if (reset) begin // @[FADD_1.scala 16:37]
      premul_b <= 24'h0; // @[FADD_1.scala 16:37]
    end else begin
      premul_b <= mulAddRecFNToRaw_preMul_io_mulAddB; // @[FADD_1.scala 104:63]
    end
    if (reset) begin // @[FADD_1.scala 17:37]
      premul_c <= 48'h0; // @[FADD_1.scala 17:37]
    end else begin
      premul_c <= mulAddRecFNToRaw_preMul_io_mulAddC; // @[FADD_1.scala 105:63]
    end
    if (reset) begin // @[FADD_1.scala 18:33]
      isSigNaNAny <= 1'h0; // @[FADD_1.scala 18:33]
    end else begin
      isSigNaNAny <= mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny; // @[FADD_1.scala 43:61]
    end
    if (reset) begin // @[FADD_1.scala 19:34]
      isNaNAOrB <= 1'h0; // @[FADD_1.scala 19:34]
    end else begin
      isNaNAOrB <= mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB; // @[FADD_1.scala 44:62]
    end
    if (reset) begin // @[FADD_1.scala 20:43]
      isInfA <= 1'h0; // @[FADD_1.scala 20:43]
    end else begin
      isInfA <= mulAddRecFNToRaw_preMul_io_toPostMul_isInfA; // @[FADD_1.scala 45:70]
    end
    if (reset) begin // @[FADD_1.scala 21:40]
      isZeroA <= 1'h0; // @[FADD_1.scala 21:40]
    end else begin
      isZeroA <= mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA; // @[FADD_1.scala 46:67]
    end
    if (reset) begin // @[FADD_1.scala 22:43]
      isInfB <= 1'h0; // @[FADD_1.scala 22:43]
    end else begin
      isInfB <= mulAddRecFNToRaw_preMul_io_toPostMul_isInfB; // @[FADD_1.scala 47:70]
    end
    if (reset) begin // @[FADD_1.scala 23:40]
      isZeroB <= 1'h0; // @[FADD_1.scala 23:40]
    end else begin
      isZeroB <= mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB; // @[FADD_1.scala 48:67]
    end
    if (reset) begin // @[FADD_1.scala 24:38]
      signProd <= 1'h0; // @[FADD_1.scala 24:38]
    end else begin
      signProd <= mulAddRecFNToRaw_preMul_io_toPostMul_signProd; // @[FADD_1.scala 49:65]
    end
    if (reset) begin // @[FADD_1.scala 25:39]
      isNaNC <= 1'h0; // @[FADD_1.scala 25:39]
    end else begin
      isNaNC <= mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC; // @[FADD_1.scala 50:66]
    end
    if (reset) begin // @[FADD_1.scala 26:42]
      isInfC <= 1'h0; // @[FADD_1.scala 26:42]
    end else begin
      isInfC <= mulAddRecFNToRaw_preMul_io_toPostMul_isInfC; // @[FADD_1.scala 51:69]
    end
    if (reset) begin // @[FADD_1.scala 27:39]
      isZeroC <= 1'h0; // @[FADD_1.scala 27:39]
    end else begin
      isZeroC <= mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC; // @[FADD_1.scala 52:66]
    end
    if (reset) begin // @[FADD_1.scala 28:36]
      sExpSum <= 10'sh0; // @[FADD_1.scala 28:36]
    end else begin
      sExpSum <= mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum; // @[FADD_1.scala 53:63]
    end
    if (reset) begin // @[FADD_1.scala 29:33]
      doSubMags <= 1'h0; // @[FADD_1.scala 29:33]
    end else begin
      doSubMags <= mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags; // @[FADD_1.scala 54:60]
    end
    if (reset) begin // @[FADD_1.scala 30:33]
      CIsDominant <= 1'h0; // @[FADD_1.scala 30:33]
    end else begin
      CIsDominant <= mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant; // @[FADD_1.scala 55:59]
    end
    if (reset) begin // @[FADD_1.scala 31:34]
      CDom_CAlignDist <= 5'h0; // @[FADD_1.scala 31:34]
    end else begin
      CDom_CAlignDist <= mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist; // @[FADD_1.scala 56:54]
    end
    if (reset) begin // @[FADD_1.scala 32:37]
      highAlignedSigC <= 26'h0; // @[FADD_1.scala 32:37]
    end else begin
      highAlignedSigC <= mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC; // @[FADD_1.scala 57:56]
    end
    if (reset) begin // @[FADD_1.scala 33:38]
      bit0AlignedSigC <= 1'h0; // @[FADD_1.scala 33:38]
    end else begin
      bit0AlignedSigC <= mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC; // @[FADD_1.scala 58:57]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  premul_a = _RAND_0[23:0];
  _RAND_1 = {1{`RANDOM}};
  premul_b = _RAND_1[23:0];
  _RAND_2 = {2{`RANDOM}};
  premul_c = _RAND_2[47:0];
  _RAND_3 = {1{`RANDOM}};
  isSigNaNAny = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  isNaNAOrB = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  isInfA = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  isZeroA = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  isInfB = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  isZeroB = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  signProd = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  isNaNC = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  isInfC = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  isZeroC = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  sExpSum = _RAND_13[9:0];
  _RAND_14 = {1{`RANDOM}};
  doSubMags = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  CIsDominant = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  CDom_CAlignDist = _RAND_16[4:0];
  _RAND_17 = {1{`RANDOM}};
  highAlignedSigC = _RAND_17[25:0];
  _RAND_18 = {1{`RANDOM}};
  bit0AlignedSigC = _RAND_18[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IST0(
  input         clock,
  input         reset,
  input         io_enable_IST0,
  input  [31:0] io_nodeid_leaf,
  input  [31:0] io_rayid_leaf,
  input  [31:0] io_hiT_in,
  input  [31:0] io_v00_x,
  input  [31:0] io_v00_y,
  input  [31:0] io_v00_z,
  input  [31:0] io_v00_w,
  input  [31:0] io_v11_in_x,
  input  [31:0] io_v11_in_y,
  input  [31:0] io_v11_in_z,
  input  [31:0] io_v11_in_w,
  input  [31:0] io_v22_in_x,
  input  [31:0] io_v22_in_y,
  input  [31:0] io_v22_in_z,
  input  [31:0] io_v22_in_w,
  input  [31:0] io_ray_o_in_x,
  input  [31:0] io_ray_o_in_y,
  input  [31:0] io_ray_o_in_z,
  input  [31:0] io_ray_d_in_x,
  input  [31:0] io_ray_d_in_y,
  input  [31:0] io_ray_d_in_z,
  input         io_RAY_AABB_1,
  input         io_RAY_AABB_2,
  input         io_break_in,
  output [31:0] io_Oz,
  output [31:0] io_invDz_div,
  output [31:0] io_nodeid_ist0_out,
  output [31:0] io_rayid_ist0_out,
  output [31:0] io_hiT_out,
  output [31:0] io_v11_out_x,
  output [31:0] io_v11_out_y,
  output [31:0] io_v11_out_z,
  output [31:0] io_v11_out_w,
  output [31:0] io_v22_out_x,
  output [31:0] io_v22_out_y,
  output [31:0] io_v22_out_z,
  output [31:0] io_v22_out_w,
  output [31:0] io_ray_o_out_x,
  output [31:0] io_ray_o_out_y,
  output [31:0] io_ray_o_out_z,
  output [31:0] io_ray_d_out_x,
  output [31:0] io_ray_d_out_y,
  output [31:0] io_ray_d_out_z,
  output        io_enable_SU_out,
  output        io_break_out,
  output        io_RAY_AABB_1_out,
  output        io_RAY_AABB_2_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [127:0] _RAND_10;
  reg [127:0] _RAND_11;
  reg [95:0] _RAND_12;
  reg [95:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [127:0] _RAND_20;
  reg [127:0] _RAND_21;
  reg [95:0] _RAND_22;
  reg [95:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [127:0] _RAND_31;
  reg [127:0] _RAND_32;
  reg [95:0] _RAND_33;
  reg [95:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [127:0] _RAND_46;
  reg [127:0] _RAND_47;
  reg [95:0] _RAND_48;
  reg [95:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [127:0] _RAND_59;
  reg [127:0] _RAND_60;
  reg [95:0] _RAND_61;
  reg [95:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
`endif // RANDOMIZE_REG_INIT
  wire  FADD_MUL_13_clock; // @[IST0.scala 73:33]
  wire  FADD_MUL_13_reset; // @[IST0.scala 73:33]
  wire [31:0] FADD_MUL_13_io_a; // @[IST0.scala 73:33]
  wire [31:0] FADD_MUL_13_io_b; // @[IST0.scala 73:33]
  wire [31:0] FADD_MUL_13_io_c; // @[IST0.scala 73:33]
  wire [31:0] FADD_MUL_13_io_out; // @[IST0.scala 73:33]
  wire  FMUL_1_clock; // @[IST0.scala 79:24]
  wire  FMUL_1_reset; // @[IST0.scala 79:24]
  wire [31:0] FMUL_1_io_a; // @[IST0.scala 79:24]
  wire [31:0] FMUL_1_io_b; // @[IST0.scala 79:24]
  wire [31:0] FMUL_1_io_out; // @[IST0.scala 79:24]
  wire  FMUL_2_clock; // @[IST0.scala 84:24]
  wire  FMUL_2_reset; // @[IST0.scala 84:24]
  wire [31:0] FMUL_2_io_a; // @[IST0.scala 84:24]
  wire [31:0] FMUL_2_io_b; // @[IST0.scala 84:24]
  wire [31:0] FMUL_2_io_out; // @[IST0.scala 84:24]
  wire  FMUL_3_clock; // @[IST0.scala 89:24]
  wire  FMUL_3_reset; // @[IST0.scala 89:24]
  wire [31:0] FMUL_3_io_a; // @[IST0.scala 89:24]
  wire [31:0] FMUL_3_io_b; // @[IST0.scala 89:24]
  wire [31:0] FMUL_3_io_out; // @[IST0.scala 89:24]
  wire  FMUL_4_clock; // @[IST0.scala 94:24]
  wire  FMUL_4_reset; // @[IST0.scala 94:24]
  wire [31:0] FMUL_4_io_a; // @[IST0.scala 94:24]
  wire [31:0] FMUL_4_io_b; // @[IST0.scala 94:24]
  wire [31:0] FMUL_4_io_out; // @[IST0.scala 94:24]
  wire  FMUL_5_clock; // @[IST0.scala 99:24]
  wire  FMUL_5_reset; // @[IST0.scala 99:24]
  wire [31:0] FMUL_5_io_a; // @[IST0.scala 99:24]
  wire [31:0] FMUL_5_io_b; // @[IST0.scala 99:24]
  wire [31:0] FMUL_5_io_out; // @[IST0.scala 99:24]
  wire  FADD_1_clock; // @[IST0.scala 164:24]
  wire  FADD_1_reset; // @[IST0.scala 164:24]
  wire [31:0] FADD_1_io_a; // @[IST0.scala 164:24]
  wire [31:0] FADD_1_io_b; // @[IST0.scala 164:24]
  wire [31:0] FADD_1_io_out; // @[IST0.scala 164:24]
  wire  FADD_2_clock; // @[IST0.scala 173:24]
  wire  FADD_2_reset; // @[IST0.scala 173:24]
  wire [31:0] FADD_2_io_a; // @[IST0.scala 173:24]
  wire [31:0] FADD_2_io_b; // @[IST0.scala 173:24]
  wire [31:0] FADD_2_io_out; // @[IST0.scala 173:24]
  wire  FADD_3_clock; // @[IST0.scala 262:24]
  wire  FADD_3_reset; // @[IST0.scala 262:24]
  wire [31:0] FADD_3_io_a; // @[IST0.scala 262:24]
  wire [31:0] FADD_3_io_b; // @[IST0.scala 262:24]
  wire [31:0] FADD_3_io_out; // @[IST0.scala 262:24]
  wire  FADD_4_clock; // @[IST0.scala 271:24]
  wire  FADD_4_reset; // @[IST0.scala 271:24]
  wire [31:0] FADD_4_io_a; // @[IST0.scala 271:24]
  wire [31:0] FADD_4_io_b; // @[IST0.scala 271:24]
  wire [31:0] FADD_4_io_out; // @[IST0.scala 271:24]
  reg [31:0] temp_0; // @[IST0.scala 42:33]
  reg [31:0] temp_1; // @[IST0.scala 43:33]
  reg [31:0] temp_2; // @[IST0.scala 44:33]
  reg [31:0] temp_3; // @[IST0.scala 45:33]
  reg [31:0] temp_4; // @[IST0.scala 46:33]
  reg [31:0] temp_5; // @[IST0.scala 47:33]
  reg  enable_1; // @[IST0.scala 49:51]
  reg [31:0] nodeid_ist0_temp_1; // @[IST0.scala 50:38]
  reg [31:0] rayid_ist0_temp_1; // @[IST0.scala 51:41]
  reg [31:0] hitT_temp_1; // @[IST0.scala 52:47]
  reg [127:0] v11_1; // @[IST0.scala 53:56]
  reg [127:0] v22_1; // @[IST0.scala 54:56]
  reg [95:0] ray_o_in_1; // @[IST0.scala 55:50]
  reg [95:0] ray_d_in_1; // @[IST0.scala 56:50]
  reg  break_1; // @[IST0.scala 57:51]
  reg  ray_aabb_1; // @[IST0.scala 58:46]
  reg  ray_aabb_2; // @[IST0.scala 59:46]
  wire [127:0] _T = {io_v11_in_w,io_v11_in_z,io_v11_in_y,io_v11_in_x}; // @[Cat.scala 30:58]
  wire [127:0] _T_1 = {io_v22_in_w,io_v22_in_z,io_v22_in_y,io_v22_in_x}; // @[Cat.scala 30:58]
  wire [95:0] _T_2 = {io_ray_o_in_z,io_ray_o_in_y,io_ray_o_in_x}; // @[Cat.scala 30:58]
  wire [95:0] _T_3 = {io_ray_d_in_z,io_ray_d_in_y,io_ray_d_in_x}; // @[Cat.scala 30:58]
  wire  hi_4 = ~io_ray_o_in_x[31]; // @[common.scala 90:20]
  wire [30:0] lo_2 = io_ray_o_in_x[30:0]; // @[common.scala 90:30]
  reg [31:0] nodeid_ist0_temp_temp; // @[IST0.scala 104:41]
  reg [31:0] rayid_ist0_temp_temp; // @[IST0.scala 105:44]
  reg [31:0] hitT_temp_temp; // @[IST0.scala 106:50]
  reg [127:0] v11_temp; // @[IST0.scala 107:59]
  reg [127:0] v22_temp; // @[IST0.scala 108:59]
  reg [95:0] ray_o_in_temp; // @[IST0.scala 109:53]
  reg [95:0] ray_d_in_temp; // @[IST0.scala 110:53]
  reg  enable_temp; // @[IST0.scala 111:54]
  reg  break_temp; // @[IST0.scala 112:54]
  reg  ray_aabb_1_temp; // @[IST0.scala 113:46]
  reg  ray_aabb_2_temp; // @[IST0.scala 114:46]
  reg [31:0] nodeid_ist0_temp_2; // @[IST0.scala 131:38]
  reg [31:0] rayid_ist0_temp_2; // @[IST0.scala 132:41]
  reg [31:0] hitT_temp_2; // @[IST0.scala 133:47]
  reg [127:0] v11_2; // @[IST0.scala 134:56]
  reg [127:0] v22_2; // @[IST0.scala 135:56]
  reg [95:0] ray_o_in_2; // @[IST0.scala 136:50]
  reg [95:0] ray_d_in_2; // @[IST0.scala 137:50]
  reg  enable_2; // @[IST0.scala 138:51]
  reg  break_2; // @[IST0.scala 139:51]
  reg  ray_aabb_1_2; // @[IST0.scala 140:43]
  reg  ray_aabb_2_2; // @[IST0.scala 141:44]
  reg [31:0] temp_6; // @[IST0.scala 156:50]
  reg [31:0] temp_7; // @[IST0.scala 157:50]
  reg [31:0] temp_0_2; // @[IST0.scala 158:47]
  reg [31:0] temp_5_2; // @[IST0.scala 159:46]
  reg [31:0] add_nodeid_ist0_temp_2; // @[IST0.scala 182:42]
  reg [31:0] add_rayid_ist0_temp_2; // @[IST0.scala 183:45]
  reg [31:0] add_hitT_temp_2; // @[IST0.scala 184:51]
  reg [127:0] add_v11_2; // @[IST0.scala 185:60]
  reg [127:0] add_v22_2; // @[IST0.scala 186:60]
  reg [95:0] add_ray_o_in_2; // @[IST0.scala 187:54]
  reg [95:0] add_ray_d_in_2; // @[IST0.scala 188:54]
  reg  add_enable_2; // @[IST0.scala 189:55]
  reg  add_break_2; // @[IST0.scala 190:55]
  reg  add_ray_aabb_1_2; // @[IST0.scala 191:47]
  reg  add_ray_aabb_2_2; // @[IST0.scala 192:48]
  reg [31:0] add_temp_0_2; // @[IST0.scala 206:51]
  reg [31:0] add_temp_5_2; // @[IST0.scala 207:50]
  reg [31:0] add2_nodeid_ist0_temp_2; // @[IST0.scala 214:43]
  reg [31:0] add2_rayid_ist0_temp_2; // @[IST0.scala 215:46]
  reg [31:0] add2_hitT_temp_2; // @[IST0.scala 216:52]
  reg [127:0] add2_v11_2; // @[IST0.scala 217:61]
  reg [127:0] add2_v22_2; // @[IST0.scala 218:61]
  reg [95:0] add2_ray_o_in_2; // @[IST0.scala 219:55]
  reg [95:0] add2_ray_d_in_2; // @[IST0.scala 220:55]
  reg  add2_enable_2; // @[IST0.scala 221:56]
  reg  add2_break_2; // @[IST0.scala 222:56]
  reg  add2_ray_aabb_1_2; // @[IST0.scala 223:48]
  reg  add2_ray_aabb_2_2; // @[IST0.scala 224:49]
  wire  hi_5 = ~temp_6[31]; // @[common.scala 90:20]
  wire [30:0] lo_3 = temp_6[30:0]; // @[common.scala 90:30]
  MY_MULADD FADD_MUL_13 ( // @[IST0.scala 73:33]
    .clock(FADD_MUL_13_clock),
    .reset(FADD_MUL_13_reset),
    .io_a(FADD_MUL_13_io_a),
    .io_b(FADD_MUL_13_io_b),
    .io_c(FADD_MUL_13_io_c),
    .io_out(FADD_MUL_13_io_out)
  );
  MY_MUL FMUL_1 ( // @[IST0.scala 79:24]
    .clock(FMUL_1_clock),
    .reset(FMUL_1_reset),
    .io_a(FMUL_1_io_a),
    .io_b(FMUL_1_io_b),
    .io_out(FMUL_1_io_out)
  );
  MY_MUL FMUL_2 ( // @[IST0.scala 84:24]
    .clock(FMUL_2_clock),
    .reset(FMUL_2_reset),
    .io_a(FMUL_2_io_a),
    .io_b(FMUL_2_io_b),
    .io_out(FMUL_2_io_out)
  );
  MY_MUL FMUL_3 ( // @[IST0.scala 89:24]
    .clock(FMUL_3_clock),
    .reset(FMUL_3_reset),
    .io_a(FMUL_3_io_a),
    .io_b(FMUL_3_io_b),
    .io_out(FMUL_3_io_out)
  );
  MY_MUL FMUL_4 ( // @[IST0.scala 94:24]
    .clock(FMUL_4_clock),
    .reset(FMUL_4_reset),
    .io_a(FMUL_4_io_a),
    .io_b(FMUL_4_io_b),
    .io_out(FMUL_4_io_out)
  );
  MY_MUL FMUL_5 ( // @[IST0.scala 99:24]
    .clock(FMUL_5_clock),
    .reset(FMUL_5_reset),
    .io_a(FMUL_5_io_a),
    .io_b(FMUL_5_io_b),
    .io_out(FMUL_5_io_out)
  );
  MY_ADD FADD_1 ( // @[IST0.scala 164:24]
    .clock(FADD_1_clock),
    .reset(FADD_1_reset),
    .io_a(FADD_1_io_a),
    .io_b(FADD_1_io_b),
    .io_out(FADD_1_io_out)
  );
  MY_ADD FADD_2 ( // @[IST0.scala 173:24]
    .clock(FADD_2_clock),
    .reset(FADD_2_reset),
    .io_a(FADD_2_io_a),
    .io_b(FADD_2_io_b),
    .io_out(FADD_2_io_out)
  );
  MY_ADD FADD_3 ( // @[IST0.scala 262:24]
    .clock(FADD_3_clock),
    .reset(FADD_3_reset),
    .io_a(FADD_3_io_a),
    .io_b(FADD_3_io_b),
    .io_out(FADD_3_io_out)
  );
  MY_ADD FADD_4 ( // @[IST0.scala 271:24]
    .clock(FADD_4_clock),
    .reset(FADD_4_reset),
    .io_a(FADD_4_io_a),
    .io_b(FADD_4_io_b),
    .io_out(FADD_4_io_out)
  );
  assign io_Oz = FADD_3_io_out; // @[IST0.scala 269:29]
  assign io_invDz_div = FADD_4_io_out; // @[IST0.scala 278:22]
  assign io_nodeid_ist0_out = add2_nodeid_ist0_temp_2; // @[IST0.scala 238:32]
  assign io_rayid_ist0_out = add2_rayid_ist0_temp_2; // @[IST0.scala 239:35]
  assign io_hiT_out = add2_hitT_temp_2; // @[IST0.scala 240:42]
  assign io_v11_out_x = add2_v11_2[31:0]; // @[IST0.scala 241:53]
  assign io_v11_out_y = add2_v11_2[63:32]; // @[IST0.scala 242:53]
  assign io_v11_out_z = add2_v11_2[95:64]; // @[IST0.scala 243:53]
  assign io_v11_out_w = add2_v11_2[127:96]; // @[IST0.scala 244:52]
  assign io_v22_out_x = add2_v22_2[31:0]; // @[IST0.scala 246:57]
  assign io_v22_out_y = add2_v22_2[63:32]; // @[IST0.scala 247:57]
  assign io_v22_out_z = add2_v22_2[95:64]; // @[IST0.scala 248:57]
  assign io_v22_out_w = add2_v22_2[127:96]; // @[IST0.scala 249:55]
  assign io_ray_o_out_x = add2_ray_o_in_2[31:0]; // @[IST0.scala 252:59]
  assign io_ray_o_out_y = add2_ray_o_in_2[63:32]; // @[IST0.scala 253:59]
  assign io_ray_o_out_z = add2_ray_o_in_2[95:64]; // @[IST0.scala 254:59]
  assign io_ray_d_out_x = add2_ray_d_in_2[31:0]; // @[IST0.scala 255:59]
  assign io_ray_d_out_y = add2_ray_d_in_2[63:32]; // @[IST0.scala 256:59]
  assign io_ray_d_out_z = add2_ray_d_in_2[95:64]; // @[IST0.scala 257:59]
  assign io_enable_SU_out = add2_enable_2; // @[IST0.scala 258:36]
  assign io_break_out = add2_break_2; // @[IST0.scala 259:42]
  assign io_RAY_AABB_1_out = add2_ray_aabb_1_2; // @[IST0.scala 260:33]
  assign io_RAY_AABB_2_out = add2_ray_aabb_2_2; // @[IST0.scala 261:33]
  assign FADD_MUL_13_clock = clock;
  assign FADD_MUL_13_reset = reset;
  assign FADD_MUL_13_io_a = {hi_4,lo_2}; // @[Cat.scala 30:58]
  assign FADD_MUL_13_io_b = io_v00_x; // @[IST0.scala 75:26]
  assign FADD_MUL_13_io_c = io_v00_w; // @[IST0.scala 76:26]
  assign FMUL_1_clock = clock;
  assign FMUL_1_reset = reset;
  assign FMUL_1_io_a = io_ray_o_in_y; // @[IST0.scala 80:21]
  assign FMUL_1_io_b = io_v00_y; // @[IST0.scala 81:21]
  assign FMUL_2_clock = clock;
  assign FMUL_2_reset = reset;
  assign FMUL_2_io_a = io_ray_o_in_z; // @[IST0.scala 85:21]
  assign FMUL_2_io_b = io_v00_z; // @[IST0.scala 86:21]
  assign FMUL_3_clock = clock;
  assign FMUL_3_reset = reset;
  assign FMUL_3_io_a = io_ray_d_in_x; // @[IST0.scala 90:21]
  assign FMUL_3_io_b = io_v00_x; // @[IST0.scala 91:21]
  assign FMUL_4_clock = clock;
  assign FMUL_4_reset = reset;
  assign FMUL_4_io_a = io_ray_d_in_y; // @[IST0.scala 95:21]
  assign FMUL_4_io_b = io_v00_y; // @[IST0.scala 96:21]
  assign FMUL_5_clock = clock;
  assign FMUL_5_reset = reset;
  assign FMUL_5_io_a = io_ray_d_in_z; // @[IST0.scala 100:21]
  assign FMUL_5_io_b = io_v00_z; // @[IST0.scala 101:21]
  assign FADD_1_clock = clock;
  assign FADD_1_reset = reset;
  assign FADD_1_io_a = temp_1; // @[IST0.scala 165:21]
  assign FADD_1_io_b = temp_2; // @[IST0.scala 166:21]
  assign FADD_2_clock = clock;
  assign FADD_2_reset = reset;
  assign FADD_2_io_a = temp_3; // @[IST0.scala 174:21]
  assign FADD_2_io_b = temp_4; // @[IST0.scala 175:21]
  assign FADD_3_clock = clock;
  assign FADD_3_reset = reset;
  assign FADD_3_io_a = add_temp_0_2; // @[IST0.scala 263:21]
  assign FADD_3_io_b = {hi_5,lo_3}; // @[Cat.scala 30:58]
  assign FADD_4_clock = clock;
  assign FADD_4_reset = reset;
  assign FADD_4_io_a = add_temp_5_2; // @[IST0.scala 272:21]
  assign FADD_4_io_b = temp_7; // @[IST0.scala 273:21]
  always @(posedge clock) begin
    if (reset) begin // @[IST0.scala 42:33]
      temp_0 <= 32'h0; // @[IST0.scala 42:33]
    end else begin
      temp_0 <= FADD_MUL_13_io_out; // @[IST0.scala 77:42]
    end
    if (reset) begin // @[IST0.scala 43:33]
      temp_1 <= 32'h0; // @[IST0.scala 43:33]
    end else begin
      temp_1 <= FMUL_1_io_out; // @[IST0.scala 82:42]
    end
    if (reset) begin // @[IST0.scala 44:33]
      temp_2 <= 32'h0; // @[IST0.scala 44:33]
    end else begin
      temp_2 <= FMUL_2_io_out; // @[IST0.scala 87:42]
    end
    if (reset) begin // @[IST0.scala 45:33]
      temp_3 <= 32'h0; // @[IST0.scala 45:33]
    end else begin
      temp_3 <= FMUL_3_io_out; // @[IST0.scala 92:42]
    end
    if (reset) begin // @[IST0.scala 46:33]
      temp_4 <= 32'h0; // @[IST0.scala 46:33]
    end else begin
      temp_4 <= FMUL_4_io_out; // @[IST0.scala 97:42]
    end
    if (reset) begin // @[IST0.scala 47:33]
      temp_5 <= 32'h0; // @[IST0.scala 47:33]
    end else begin
      temp_5 <= FMUL_5_io_out; // @[IST0.scala 102:42]
    end
    if (reset) begin // @[IST0.scala 49:51]
      enable_1 <= 1'h0; // @[IST0.scala 49:51]
    end else begin
      enable_1 <= io_enable_IST0; // @[IST0.scala 68:42]
    end
    if (reset) begin // @[IST0.scala 50:38]
      nodeid_ist0_temp_1 <= 32'sh0; // @[IST0.scala 50:38]
    end else begin
      nodeid_ist0_temp_1 <= io_nodeid_leaf; // @[IST0.scala 61:29]
    end
    if (reset) begin // @[IST0.scala 51:41]
      rayid_ist0_temp_1 <= 32'h0; // @[IST0.scala 51:41]
    end else begin
      rayid_ist0_temp_1 <= io_rayid_leaf; // @[IST0.scala 62:32]
    end
    if (reset) begin // @[IST0.scala 52:47]
      hitT_temp_1 <= 32'h0; // @[IST0.scala 52:47]
    end else begin
      hitT_temp_1 <= io_hiT_in; // @[IST0.scala 63:38]
    end
    if (reset) begin // @[IST0.scala 53:56]
      v11_1 <= 128'h0; // @[IST0.scala 53:56]
    end else begin
      v11_1 <= _T; // @[IST0.scala 64:46]
    end
    if (reset) begin // @[IST0.scala 54:56]
      v22_1 <= 128'h0; // @[IST0.scala 54:56]
    end else begin
      v22_1 <= _T_1; // @[IST0.scala 65:46]
    end
    if (reset) begin // @[IST0.scala 55:50]
      ray_o_in_1 <= 96'h0; // @[IST0.scala 55:50]
    end else begin
      ray_o_in_1 <= _T_2; // @[IST0.scala 66:40]
    end
    if (reset) begin // @[IST0.scala 56:50]
      ray_d_in_1 <= 96'h0; // @[IST0.scala 56:50]
    end else begin
      ray_d_in_1 <= _T_3; // @[IST0.scala 67:40]
    end
    if (reset) begin // @[IST0.scala 57:51]
      break_1 <= 1'h0; // @[IST0.scala 57:51]
    end else begin
      break_1 <= io_break_in; // @[IST0.scala 69:44]
    end
    if (reset) begin // @[IST0.scala 58:46]
      ray_aabb_1 <= 1'h0; // @[IST0.scala 58:46]
    end else begin
      ray_aabb_1 <= io_RAY_AABB_1; // @[IST0.scala 70:40]
    end
    if (reset) begin // @[IST0.scala 59:46]
      ray_aabb_2 <= 1'h0; // @[IST0.scala 59:46]
    end else begin
      ray_aabb_2 <= io_RAY_AABB_2; // @[IST0.scala 71:40]
    end
    if (reset) begin // @[IST0.scala 104:41]
      nodeid_ist0_temp_temp <= 32'sh0; // @[IST0.scala 104:41]
    end else begin
      nodeid_ist0_temp_temp <= nodeid_ist0_temp_1; // @[IST0.scala 116:32]
    end
    if (reset) begin // @[IST0.scala 105:44]
      rayid_ist0_temp_temp <= 32'h0; // @[IST0.scala 105:44]
    end else begin
      rayid_ist0_temp_temp <= rayid_ist0_temp_1; // @[IST0.scala 117:35]
    end
    if (reset) begin // @[IST0.scala 106:50]
      hitT_temp_temp <= 32'h0; // @[IST0.scala 106:50]
    end else begin
      hitT_temp_temp <= hitT_temp_1; // @[IST0.scala 118:41]
    end
    if (reset) begin // @[IST0.scala 107:59]
      v11_temp <= 128'h0; // @[IST0.scala 107:59]
    end else begin
      v11_temp <= v11_1; // @[IST0.scala 119:49]
    end
    if (reset) begin // @[IST0.scala 108:59]
      v22_temp <= 128'h0; // @[IST0.scala 108:59]
    end else begin
      v22_temp <= v22_1; // @[IST0.scala 120:49]
    end
    if (reset) begin // @[IST0.scala 109:53]
      ray_o_in_temp <= 96'h0; // @[IST0.scala 109:53]
    end else begin
      ray_o_in_temp <= ray_o_in_1; // @[IST0.scala 121:43]
    end
    if (reset) begin // @[IST0.scala 110:53]
      ray_d_in_temp <= 96'h0; // @[IST0.scala 110:53]
    end else begin
      ray_d_in_temp <= ray_d_in_1; // @[IST0.scala 122:43]
    end
    if (reset) begin // @[IST0.scala 111:54]
      enable_temp <= 1'h0; // @[IST0.scala 111:54]
    end else begin
      enable_temp <= enable_1; // @[IST0.scala 123:45]
    end
    if (reset) begin // @[IST0.scala 112:54]
      break_temp <= 1'h0; // @[IST0.scala 112:54]
    end else begin
      break_temp <= break_1; // @[IST0.scala 124:47]
    end
    if (reset) begin // @[IST0.scala 113:46]
      ray_aabb_1_temp <= 1'h0; // @[IST0.scala 113:46]
    end else begin
      ray_aabb_1_temp <= ray_aabb_1; // @[IST0.scala 125:39]
    end
    if (reset) begin // @[IST0.scala 114:46]
      ray_aabb_2_temp <= 1'h0; // @[IST0.scala 114:46]
    end else begin
      ray_aabb_2_temp <= ray_aabb_2; // @[IST0.scala 126:39]
    end
    if (reset) begin // @[IST0.scala 131:38]
      nodeid_ist0_temp_2 <= 32'sh0; // @[IST0.scala 131:38]
    end else begin
      nodeid_ist0_temp_2 <= nodeid_ist0_temp_temp; // @[IST0.scala 143:29]
    end
    if (reset) begin // @[IST0.scala 132:41]
      rayid_ist0_temp_2 <= 32'h0; // @[IST0.scala 132:41]
    end else begin
      rayid_ist0_temp_2 <= rayid_ist0_temp_temp; // @[IST0.scala 144:32]
    end
    if (reset) begin // @[IST0.scala 133:47]
      hitT_temp_2 <= 32'h0; // @[IST0.scala 133:47]
    end else begin
      hitT_temp_2 <= hitT_temp_temp; // @[IST0.scala 145:38]
    end
    if (reset) begin // @[IST0.scala 134:56]
      v11_2 <= 128'h0; // @[IST0.scala 134:56]
    end else begin
      v11_2 <= v11_temp; // @[IST0.scala 146:46]
    end
    if (reset) begin // @[IST0.scala 135:56]
      v22_2 <= 128'h0; // @[IST0.scala 135:56]
    end else begin
      v22_2 <= v22_temp; // @[IST0.scala 147:46]
    end
    if (reset) begin // @[IST0.scala 136:50]
      ray_o_in_2 <= 96'h0; // @[IST0.scala 136:50]
    end else begin
      ray_o_in_2 <= ray_o_in_temp; // @[IST0.scala 148:40]
    end
    if (reset) begin // @[IST0.scala 137:50]
      ray_d_in_2 <= 96'h0; // @[IST0.scala 137:50]
    end else begin
      ray_d_in_2 <= ray_d_in_temp; // @[IST0.scala 149:40]
    end
    if (reset) begin // @[IST0.scala 138:51]
      enable_2 <= 1'h0; // @[IST0.scala 138:51]
    end else begin
      enable_2 <= enable_temp; // @[IST0.scala 152:42]
    end
    if (reset) begin // @[IST0.scala 139:51]
      break_2 <= 1'h0; // @[IST0.scala 139:51]
    end else begin
      break_2 <= break_temp; // @[IST0.scala 153:44]
    end
    if (reset) begin // @[IST0.scala 140:43]
      ray_aabb_1_2 <= 1'h0; // @[IST0.scala 140:43]
    end else begin
      ray_aabb_1_2 <= ray_aabb_1_temp; // @[IST0.scala 154:37]
    end
    if (reset) begin // @[IST0.scala 141:44]
      ray_aabb_2_2 <= 1'h0; // @[IST0.scala 141:44]
    end else begin
      ray_aabb_2_2 <= ray_aabb_2_temp; // @[IST0.scala 155:37]
    end
    if (reset) begin // @[IST0.scala 156:50]
      temp_6 <= 32'h0; // @[IST0.scala 156:50]
    end else begin
      temp_6 <= FADD_1_io_out; // @[IST0.scala 171:26]
    end
    if (reset) begin // @[IST0.scala 157:50]
      temp_7 <= 32'h0; // @[IST0.scala 157:50]
    end else begin
      temp_7 <= FADD_2_io_out; // @[IST0.scala 180:26]
    end
    if (reset) begin // @[IST0.scala 158:47]
      temp_0_2 <= 32'h0; // @[IST0.scala 158:47]
    end else begin
      temp_0_2 <= temp_0; // @[IST0.scala 161:41]
    end
    if (reset) begin // @[IST0.scala 159:46]
      temp_5_2 <= 32'h0; // @[IST0.scala 159:46]
    end else begin
      temp_5_2 <= temp_5; // @[IST0.scala 162:41]
    end
    if (reset) begin // @[IST0.scala 182:42]
      add_nodeid_ist0_temp_2 <= 32'sh0; // @[IST0.scala 182:42]
    end else begin
      add_nodeid_ist0_temp_2 <= nodeid_ist0_temp_2; // @[IST0.scala 194:33]
    end
    if (reset) begin // @[IST0.scala 183:45]
      add_rayid_ist0_temp_2 <= 32'h0; // @[IST0.scala 183:45]
    end else begin
      add_rayid_ist0_temp_2 <= rayid_ist0_temp_2; // @[IST0.scala 195:36]
    end
    if (reset) begin // @[IST0.scala 184:51]
      add_hitT_temp_2 <= 32'h0; // @[IST0.scala 184:51]
    end else begin
      add_hitT_temp_2 <= hitT_temp_2; // @[IST0.scala 196:42]
    end
    if (reset) begin // @[IST0.scala 185:60]
      add_v11_2 <= 128'h0; // @[IST0.scala 185:60]
    end else begin
      add_v11_2 <= v11_2; // @[IST0.scala 197:50]
    end
    if (reset) begin // @[IST0.scala 186:60]
      add_v22_2 <= 128'h0; // @[IST0.scala 186:60]
    end else begin
      add_v22_2 <= v22_2; // @[IST0.scala 198:50]
    end
    if (reset) begin // @[IST0.scala 187:54]
      add_ray_o_in_2 <= 96'h0; // @[IST0.scala 187:54]
    end else begin
      add_ray_o_in_2 <= ray_o_in_2; // @[IST0.scala 199:44]
    end
    if (reset) begin // @[IST0.scala 188:54]
      add_ray_d_in_2 <= 96'h0; // @[IST0.scala 188:54]
    end else begin
      add_ray_d_in_2 <= ray_d_in_2; // @[IST0.scala 200:44]
    end
    if (reset) begin // @[IST0.scala 189:55]
      add_enable_2 <= 1'h0; // @[IST0.scala 189:55]
    end else begin
      add_enable_2 <= enable_2; // @[IST0.scala 201:46]
    end
    if (reset) begin // @[IST0.scala 190:55]
      add_break_2 <= 1'h0; // @[IST0.scala 190:55]
    end else begin
      add_break_2 <= break_2; // @[IST0.scala 202:48]
    end
    if (reset) begin // @[IST0.scala 191:47]
      add_ray_aabb_1_2 <= 1'h0; // @[IST0.scala 191:47]
    end else begin
      add_ray_aabb_1_2 <= ray_aabb_1_2; // @[IST0.scala 203:41]
    end
    if (reset) begin // @[IST0.scala 192:48]
      add_ray_aabb_2_2 <= 1'h0; // @[IST0.scala 192:48]
    end else begin
      add_ray_aabb_2_2 <= ray_aabb_2_2; // @[IST0.scala 204:41]
    end
    if (reset) begin // @[IST0.scala 206:51]
      add_temp_0_2 <= 32'h0; // @[IST0.scala 206:51]
    end else begin
      add_temp_0_2 <= temp_0_2; // @[IST0.scala 209:45]
    end
    if (reset) begin // @[IST0.scala 207:50]
      add_temp_5_2 <= 32'h0; // @[IST0.scala 207:50]
    end else begin
      add_temp_5_2 <= temp_5_2; // @[IST0.scala 210:45]
    end
    if (reset) begin // @[IST0.scala 214:43]
      add2_nodeid_ist0_temp_2 <= 32'sh0; // @[IST0.scala 214:43]
    end else begin
      add2_nodeid_ist0_temp_2 <= add_nodeid_ist0_temp_2; // @[IST0.scala 226:34]
    end
    if (reset) begin // @[IST0.scala 215:46]
      add2_rayid_ist0_temp_2 <= 32'h0; // @[IST0.scala 215:46]
    end else begin
      add2_rayid_ist0_temp_2 <= add_rayid_ist0_temp_2; // @[IST0.scala 227:37]
    end
    if (reset) begin // @[IST0.scala 216:52]
      add2_hitT_temp_2 <= 32'h0; // @[IST0.scala 216:52]
    end else begin
      add2_hitT_temp_2 <= add_hitT_temp_2; // @[IST0.scala 228:43]
    end
    if (reset) begin // @[IST0.scala 217:61]
      add2_v11_2 <= 128'h0; // @[IST0.scala 217:61]
    end else begin
      add2_v11_2 <= add_v11_2; // @[IST0.scala 229:51]
    end
    if (reset) begin // @[IST0.scala 218:61]
      add2_v22_2 <= 128'h0; // @[IST0.scala 218:61]
    end else begin
      add2_v22_2 <= add_v22_2; // @[IST0.scala 230:51]
    end
    if (reset) begin // @[IST0.scala 219:55]
      add2_ray_o_in_2 <= 96'h0; // @[IST0.scala 219:55]
    end else begin
      add2_ray_o_in_2 <= add_ray_o_in_2; // @[IST0.scala 231:45]
    end
    if (reset) begin // @[IST0.scala 220:55]
      add2_ray_d_in_2 <= 96'h0; // @[IST0.scala 220:55]
    end else begin
      add2_ray_d_in_2 <= add_ray_d_in_2; // @[IST0.scala 232:45]
    end
    if (reset) begin // @[IST0.scala 221:56]
      add2_enable_2 <= 1'h0; // @[IST0.scala 221:56]
    end else begin
      add2_enable_2 <= add_enable_2; // @[IST0.scala 233:47]
    end
    if (reset) begin // @[IST0.scala 222:56]
      add2_break_2 <= 1'h0; // @[IST0.scala 222:56]
    end else begin
      add2_break_2 <= add_break_2; // @[IST0.scala 234:49]
    end
    if (reset) begin // @[IST0.scala 223:48]
      add2_ray_aabb_1_2 <= 1'h0; // @[IST0.scala 223:48]
    end else begin
      add2_ray_aabb_1_2 <= add_ray_aabb_1_2; // @[IST0.scala 235:42]
    end
    if (reset) begin // @[IST0.scala 224:49]
      add2_ray_aabb_2_2 <= 1'h0; // @[IST0.scala 224:49]
    end else begin
      add2_ray_aabb_2_2 <= add_ray_aabb_2_2; // @[IST0.scala 236:42]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  temp_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  temp_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  temp_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  temp_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  temp_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  temp_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  enable_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  nodeid_ist0_temp_1 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  rayid_ist0_temp_1 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  hitT_temp_1 = _RAND_9[31:0];
  _RAND_10 = {4{`RANDOM}};
  v11_1 = _RAND_10[127:0];
  _RAND_11 = {4{`RANDOM}};
  v22_1 = _RAND_11[127:0];
  _RAND_12 = {3{`RANDOM}};
  ray_o_in_1 = _RAND_12[95:0];
  _RAND_13 = {3{`RANDOM}};
  ray_d_in_1 = _RAND_13[95:0];
  _RAND_14 = {1{`RANDOM}};
  break_1 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  ray_aabb_1 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  ray_aabb_2 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  nodeid_ist0_temp_temp = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  rayid_ist0_temp_temp = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  hitT_temp_temp = _RAND_19[31:0];
  _RAND_20 = {4{`RANDOM}};
  v11_temp = _RAND_20[127:0];
  _RAND_21 = {4{`RANDOM}};
  v22_temp = _RAND_21[127:0];
  _RAND_22 = {3{`RANDOM}};
  ray_o_in_temp = _RAND_22[95:0];
  _RAND_23 = {3{`RANDOM}};
  ray_d_in_temp = _RAND_23[95:0];
  _RAND_24 = {1{`RANDOM}};
  enable_temp = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  break_temp = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  ray_aabb_1_temp = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  ray_aabb_2_temp = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  nodeid_ist0_temp_2 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  rayid_ist0_temp_2 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  hitT_temp_2 = _RAND_30[31:0];
  _RAND_31 = {4{`RANDOM}};
  v11_2 = _RAND_31[127:0];
  _RAND_32 = {4{`RANDOM}};
  v22_2 = _RAND_32[127:0];
  _RAND_33 = {3{`RANDOM}};
  ray_o_in_2 = _RAND_33[95:0];
  _RAND_34 = {3{`RANDOM}};
  ray_d_in_2 = _RAND_34[95:0];
  _RAND_35 = {1{`RANDOM}};
  enable_2 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  break_2 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  ray_aabb_1_2 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  ray_aabb_2_2 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  temp_6 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  temp_7 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  temp_0_2 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  temp_5_2 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  add_nodeid_ist0_temp_2 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  add_rayid_ist0_temp_2 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  add_hitT_temp_2 = _RAND_45[31:0];
  _RAND_46 = {4{`RANDOM}};
  add_v11_2 = _RAND_46[127:0];
  _RAND_47 = {4{`RANDOM}};
  add_v22_2 = _RAND_47[127:0];
  _RAND_48 = {3{`RANDOM}};
  add_ray_o_in_2 = _RAND_48[95:0];
  _RAND_49 = {3{`RANDOM}};
  add_ray_d_in_2 = _RAND_49[95:0];
  _RAND_50 = {1{`RANDOM}};
  add_enable_2 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  add_break_2 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  add_ray_aabb_1_2 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  add_ray_aabb_2_2 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  add_temp_0_2 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  add_temp_5_2 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  add2_nodeid_ist0_temp_2 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  add2_rayid_ist0_temp_2 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  add2_hitT_temp_2 = _RAND_58[31:0];
  _RAND_59 = {4{`RANDOM}};
  add2_v11_2 = _RAND_59[127:0];
  _RAND_60 = {4{`RANDOM}};
  add2_v22_2 = _RAND_60[127:0];
  _RAND_61 = {3{`RANDOM}};
  add2_ray_o_in_2 = _RAND_61[95:0];
  _RAND_62 = {3{`RANDOM}};
  add2_ray_d_in_2 = _RAND_62[95:0];
  _RAND_63 = {1{`RANDOM}};
  add2_enable_2 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  add2_break_2 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  add2_ray_aabb_1_2 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  add2_ray_aabb_2_2 = _RAND_66[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module lookupC(
  input  [5:0]  io_addr,
  output [23:0] io_out
);
  wire [9:0] _GEN_0 = io_addr == 6'h3f ? 10'h206 : 10'h0; // @[lookups.scala 386:43 lookups.scala 386:51 lookups.scala 387:27]
  wire [9:0] _GEN_1 = io_addr == 6'h3e ? 10'h212 : _GEN_0; // @[lookups.scala 385:43 lookups.scala 385:51]
  wire [9:0] _GEN_2 = io_addr == 6'h3d ? 10'h21f : _GEN_1; // @[lookups.scala 384:43 lookups.scala 384:51]
  wire [9:0] _GEN_3 = io_addr == 6'h3c ? 10'h22c : _GEN_2; // @[lookups.scala 383:43 lookups.scala 383:51]
  wire [9:0] _GEN_4 = io_addr == 6'h3b ? 10'h23a : _GEN_3; // @[lookups.scala 382:43 lookups.scala 382:51]
  wire [9:0] _GEN_5 = io_addr == 6'h3a ? 10'h248 : _GEN_4; // @[lookups.scala 381:43 lookups.scala 381:51]
  wire [9:0] _GEN_6 = io_addr == 6'h39 ? 10'h256 : _GEN_5; // @[lookups.scala 380:43 lookups.scala 380:51]
  wire [9:0] _GEN_7 = io_addr == 6'h38 ? 10'h265 : _GEN_6; // @[lookups.scala 379:43 lookups.scala 379:51]
  wire [9:0] _GEN_8 = io_addr == 6'h37 ? 10'h275 : _GEN_7; // @[lookups.scala 377:43 lookups.scala 377:51]
  wire [9:0] _GEN_9 = io_addr == 6'h36 ? 10'h285 : _GEN_8; // @[lookups.scala 376:43 lookups.scala 376:51]
  wire [9:0] _GEN_10 = io_addr == 6'h35 ? 10'h295 : _GEN_9; // @[lookups.scala 375:43 lookups.scala 375:51]
  wire [9:0] _GEN_11 = io_addr == 6'h34 ? 10'h2a7 : _GEN_10; // @[lookups.scala 374:43 lookups.scala 374:51]
  wire [9:0] _GEN_12 = io_addr == 6'h33 ? 10'h2b8 : _GEN_11; // @[lookups.scala 373:43 lookups.scala 373:51]
  wire [9:0] _GEN_13 = io_addr == 6'h32 ? 10'h2cb : _GEN_12; // @[lookups.scala 372:43 lookups.scala 372:51]
  wire [9:0] _GEN_14 = io_addr == 6'h31 ? 10'h2de : _GEN_13; // @[lookups.scala 371:43 lookups.scala 371:51]
  wire [9:0] _GEN_15 = io_addr == 6'h30 ? 10'h2f2 : _GEN_14; // @[lookups.scala 370:43 lookups.scala 370:51]
  wire [9:0] _GEN_16 = io_addr == 6'h2f ? 10'h306 : _GEN_15; // @[lookups.scala 368:43 lookups.scala 368:51]
  wire [9:0] _GEN_17 = io_addr == 6'h2e ? 10'h31b : _GEN_16; // @[lookups.scala 367:43 lookups.scala 367:51]
  wire [9:0] _GEN_18 = io_addr == 6'h2d ? 10'h331 : _GEN_17; // @[lookups.scala 366:43 lookups.scala 366:51]
  wire [9:0] _GEN_19 = io_addr == 6'h2c ? 10'h348 : _GEN_18; // @[lookups.scala 365:43 lookups.scala 365:51]
  wire [9:0] _GEN_20 = io_addr == 6'h2b ? 10'h360 : _GEN_19; // @[lookups.scala 364:43 lookups.scala 364:51]
  wire [9:0] _GEN_21 = io_addr == 6'h2a ? 10'h378 : _GEN_20; // @[lookups.scala 363:43 lookups.scala 363:51]
  wire [9:0] _GEN_22 = io_addr == 6'h29 ? 10'h392 : _GEN_21; // @[lookups.scala 362:43 lookups.scala 362:51]
  wire [9:0] _GEN_23 = io_addr == 6'h28 ? 10'h3ac : _GEN_22; // @[lookups.scala 361:43 lookups.scala 361:51]
  wire [9:0] _GEN_24 = io_addr == 6'h27 ? 10'h3c8 : _GEN_23; // @[lookups.scala 359:43 lookups.scala 359:51]
  wire [9:0] _GEN_25 = io_addr == 6'h26 ? 10'h3e5 : _GEN_24; // @[lookups.scala 358:43 lookups.scala 358:51]
  wire [10:0] _GEN_26 = io_addr == 6'h25 ? 11'h402 : {{1'd0}, _GEN_25}; // @[lookups.scala 357:43 lookups.scala 357:51]
  wire [10:0] _GEN_27 = io_addr == 6'h24 ? 11'h421 : _GEN_26; // @[lookups.scala 356:43 lookups.scala 356:51]
  wire [10:0] _GEN_28 = io_addr == 6'h23 ? 11'h442 : _GEN_27; // @[lookups.scala 355:43 lookups.scala 355:51]
  wire [10:0] _GEN_29 = io_addr == 6'h22 ? 11'h463 : _GEN_28; // @[lookups.scala 354:43 lookups.scala 354:51]
  wire [10:0] _GEN_30 = io_addr == 6'h21 ? 11'h486 : _GEN_29; // @[lookups.scala 353:43 lookups.scala 353:51]
  wire [10:0] _GEN_31 = io_addr == 6'h20 ? 11'h4aa : _GEN_30; // @[lookups.scala 352:43 lookups.scala 352:51]
  wire [10:0] _GEN_32 = io_addr == 6'h1f ? 11'h4d0 : _GEN_31; // @[lookups.scala 350:43 lookups.scala 350:51]
  wire [10:0] _GEN_33 = io_addr == 6'h1e ? 11'h4f8 : _GEN_32; // @[lookups.scala 349:43 lookups.scala 349:51]
  wire [10:0] _GEN_34 = io_addr == 6'h1d ? 11'h521 : _GEN_33; // @[lookups.scala 348:43 lookups.scala 348:51]
  wire [10:0] _GEN_35 = io_addr == 6'h1c ? 11'h54c : _GEN_34; // @[lookups.scala 347:43 lookups.scala 347:51]
  wire [10:0] _GEN_36 = io_addr == 6'h1b ? 11'h579 : _GEN_35; // @[lookups.scala 346:43 lookups.scala 346:51]
  wire [10:0] _GEN_37 = io_addr == 6'h1a ? 11'h5a8 : _GEN_36; // @[lookups.scala 345:43 lookups.scala 345:51]
  wire [10:0] _GEN_38 = io_addr == 6'h19 ? 11'h5d9 : _GEN_37; // @[lookups.scala 344:43 lookups.scala 344:51]
  wire [10:0] _GEN_39 = io_addr == 6'h18 ? 11'h60d : _GEN_38; // @[lookups.scala 343:43 lookups.scala 343:51]
  wire [10:0] _GEN_40 = io_addr == 6'h17 ? 11'h642 : _GEN_39; // @[lookups.scala 341:43 lookups.scala 341:51]
  wire [10:0] _GEN_41 = io_addr == 6'h16 ? 11'h67b : _GEN_40; // @[lookups.scala 340:43 lookups.scala 340:51]
  wire [10:0] _GEN_42 = io_addr == 6'h15 ? 11'h6b5 : _GEN_41; // @[lookups.scala 339:43 lookups.scala 339:51]
  wire [10:0] _GEN_43 = io_addr == 6'h14 ? 11'h6f3 : _GEN_42; // @[lookups.scala 338:43 lookups.scala 338:51]
  wire [10:0] _GEN_44 = io_addr == 6'h13 ? 11'h734 : _GEN_43; // @[lookups.scala 337:43 lookups.scala 337:51]
  wire [10:0] _GEN_45 = io_addr == 6'h12 ? 11'h778 : _GEN_44; // @[lookups.scala 336:43 lookups.scala 336:51]
  wire [10:0] _GEN_46 = io_addr == 6'h11 ? 11'h7bf : _GEN_45; // @[lookups.scala 335:43 lookups.scala 335:51]
  wire [11:0] _GEN_47 = io_addr == 6'h10 ? 12'h80a : {{1'd0}, _GEN_46}; // @[lookups.scala 334:43 lookups.scala 334:51]
  wire [11:0] _GEN_48 = io_addr == 6'hf ? 12'h859 : _GEN_47; // @[lookups.scala 332:43 lookups.scala 332:51]
  wire [11:0] _GEN_49 = io_addr == 6'he ? 12'h8ab : _GEN_48; // @[lookups.scala 331:43 lookups.scala 331:51]
  wire [11:0] _GEN_50 = io_addr == 6'hd ? 12'h902 : _GEN_49; // @[lookups.scala 330:43 lookups.scala 330:51]
  wire [11:0] _GEN_51 = io_addr == 6'hc ? 12'h95e : _GEN_50; // @[lookups.scala 329:43 lookups.scala 329:51]
  wire [11:0] _GEN_52 = io_addr == 6'hb ? 12'h9bf : _GEN_51; // @[lookups.scala 328:43 lookups.scala 328:51]
  wire [11:0] _GEN_53 = io_addr == 6'ha ? 12'ha24 : _GEN_52; // @[lookups.scala 327:43 lookups.scala 327:51]
  wire [11:0] _GEN_54 = io_addr == 6'h9 ? 12'ha90 : _GEN_53; // @[lookups.scala 326:43 lookups.scala 326:51]
  wire [11:0] _GEN_55 = io_addr == 6'h8 ? 12'hb01 : _GEN_54; // @[lookups.scala 325:43 lookups.scala 325:51]
  wire [11:0] _GEN_56 = io_addr == 6'h7 ? 12'hb79 : _GEN_55; // @[lookups.scala 323:43 lookups.scala 323:51]
  wire [11:0] _GEN_57 = io_addr == 6'h6 ? 12'hbf8 : _GEN_56; // @[lookups.scala 322:43 lookups.scala 322:51]
  wire [11:0] _GEN_58 = io_addr == 6'h5 ? 12'hc7e : _GEN_57; // @[lookups.scala 321:43 lookups.scala 321:51]
  wire [11:0] _GEN_59 = io_addr == 6'h4 ? 12'hd0c : _GEN_58; // @[lookups.scala 320:43 lookups.scala 320:51]
  wire [11:0] _GEN_60 = io_addr == 6'h3 ? 12'hda3 : _GEN_59; // @[lookups.scala 319:43 lookups.scala 319:51]
  wire [11:0] _GEN_61 = io_addr == 6'h2 ? 12'he43 : _GEN_60; // @[lookups.scala 318:43 lookups.scala 318:51]
  wire [11:0] _GEN_62 = io_addr == 6'h1 ? 12'heed : _GEN_61; // @[lookups.scala 317:43 lookups.scala 317:51]
  wire [11:0] _GEN_63 = io_addr == 6'h0 ? 12'hfa1 : _GEN_62; // @[lookups.scala 316:38 lookups.scala 316:46]
  assign io_out = {{12'd0}, _GEN_63}; // @[lookups.scala 316:38 lookups.scala 316:46]
endmodule
module lookupL(
  input  [5:0]  io_addr,
  output [26:0] io_out
);
  wire [26:0] _GEN_0 = io_addr == 6'h3f ? 27'h4081020 : 27'h0; // @[lookups.scala 134:43 lookups.scala 134:51 lookups.scala 135:27]
  wire [26:0] _GEN_1 = io_addr == 6'h3e ? 27'h4104104 : _GEN_0; // @[lookups.scala 133:43 lookups.scala 133:51]
  wire [26:0] _GEN_2 = io_addr == 6'h3d ? 27'h4189374 : _GEN_1; // @[lookups.scala 132:43 lookups.scala 132:51]
  wire [26:0] _GEN_3 = io_addr == 6'h3c ? 27'h4210842 : _GEN_2; // @[lookups.scala 131:43 lookups.scala 131:51]
  wire [26:0] _GEN_4 = io_addr == 6'h3b ? 27'h429a042 : _GEN_3; // @[lookups.scala 130:43 lookups.scala 130:51]
  wire [26:0] _GEN_5 = io_addr == 6'h3a ? 27'h4325c53 : _GEN_4; // @[lookups.scala 129:43 lookups.scala 129:51]
  wire [26:0] _GEN_6 = io_addr == 6'h39 ? 27'h43b3d5a : _GEN_5; // @[lookups.scala 128:43 lookups.scala 128:51]
  wire [26:0] _GEN_7 = io_addr == 6'h38 ? 27'h4444444 : _GEN_6; // @[lookups.scala 127:43 lookups.scala 127:51]
  wire [26:0] _GEN_8 = io_addr == 6'h37 ? 27'h44d7204 : _GEN_7; // @[lookups.scala 125:43 lookups.scala 125:51]
  wire [26:0] _GEN_9 = io_addr == 6'h36 ? 27'h456c797 : _GEN_8; // @[lookups.scala 124:43 lookups.scala 124:51]
  wire [26:0] _GEN_10 = io_addr == 6'h35 ? 27'h4604604 : _GEN_9; // @[lookups.scala 123:43 lookups.scala 123:51]
  wire [26:0] _GEN_11 = io_addr == 6'h34 ? 27'h469ee58 : _GEN_10; // @[lookups.scala 122:43 lookups.scala 122:51]
  wire [26:0] _GEN_12 = io_addr == 6'h33 ? 27'h473c1ab : _GEN_11; // @[lookups.scala 121:43 lookups.scala 121:51]
  wire [26:0] _GEN_13 = io_addr == 6'h32 ? 27'h47dc11f : _GEN_12; // @[lookups.scala 120:43 lookups.scala 120:51]
  wire [26:0] _GEN_14 = io_addr == 6'h31 ? 27'h487ede0 : _GEN_13; // @[lookups.scala 119:43 lookups.scala 119:51]
  wire [26:0] _GEN_15 = io_addr == 6'h30 ? 27'h4924924 : _GEN_14; // @[lookups.scala 118:43 lookups.scala 118:51]
  wire [26:0] _GEN_16 = io_addr == 6'h2f ? 27'h49cd42e : _GEN_15; // @[lookups.scala 116:43 lookups.scala 116:51]
  wire [26:0] _GEN_17 = io_addr == 6'h2e ? 27'h4a7904a : _GEN_16; // @[lookups.scala 115:43 lookups.scala 115:51]
  wire [26:0] _GEN_18 = io_addr == 6'h2d ? 27'h4b27ed3 : _GEN_17; // @[lookups.scala 114:43 lookups.scala 114:51]
  wire [26:0] _GEN_19 = io_addr == 6'h2c ? 27'h4bda12f : _GEN_18; // @[lookups.scala 113:43 lookups.scala 113:51]
  wire [26:0] _GEN_20 = io_addr == 6'h2b ? 27'h4c8f8d2 : _GEN_19; // @[lookups.scala 112:43 lookups.scala 112:51]
  wire [26:0] _GEN_21 = io_addr == 6'h2a ? 27'h4d4873e : _GEN_20; // @[lookups.scala 111:43 lookups.scala 111:51]
  wire [26:0] _GEN_22 = io_addr == 6'h29 ? 27'h4e04e04 : _GEN_21; // @[lookups.scala 110:43 lookups.scala 110:51]
  wire [26:0] _GEN_23 = io_addr == 6'h28 ? 27'h4ec4ec4 : _GEN_22; // @[lookups.scala 109:43 lookups.scala 109:51]
  wire [26:0] _GEN_24 = io_addr == 6'h27 ? 27'h4f88b2f : _GEN_23; // @[lookups.scala 107:43 lookups.scala 107:51]
  wire [26:0] _GEN_25 = io_addr == 6'h26 ? 27'h5050505 : _GEN_24; // @[lookups.scala 106:43 lookups.scala 106:51]
  wire [26:0] _GEN_26 = io_addr == 6'h25 ? 27'h511be19 : _GEN_25; // @[lookups.scala 105:43 lookups.scala 105:51]
  wire [26:0] _GEN_27 = io_addr == 6'h24 ? 27'h51eb851 : _GEN_26; // @[lookups.scala 104:43 lookups.scala 104:51]
  wire [26:0] _GEN_28 = io_addr == 6'h23 ? 27'h52bf5a8 : _GEN_27; // @[lookups.scala 103:43 lookups.scala 103:51]
  wire [26:0] _GEN_29 = io_addr == 6'h22 ? 27'h5397829 : _GEN_28; // @[lookups.scala 102:43 lookups.scala 102:51]
  wire [26:0] _GEN_30 = io_addr == 6'h21 ? 27'h54741fa : _GEN_29; // @[lookups.scala 101:43 lookups.scala 101:51]
  wire [26:0] _GEN_31 = io_addr == 6'h20 ? 27'h5555555 : _GEN_30; // @[lookups.scala 100:43 lookups.scala 100:51]
  wire [26:0] _GEN_32 = io_addr == 6'h1f ? 27'h563b48c : _GEN_31; // @[lookups.scala 98:43 lookups.scala 98:51]
  wire [26:0] _GEN_33 = io_addr == 6'h1e ? 27'h572620a : _GEN_32; // @[lookups.scala 97:43 lookups.scala 97:51]
  wire [26:0] _GEN_34 = io_addr == 6'h1d ? 27'h5816058 : _GEN_33; // @[lookups.scala 96:43 lookups.scala 96:51]
  wire [26:0] _GEN_35 = io_addr == 6'h1c ? 27'h590b216 : _GEN_34; // @[lookups.scala 95:43 lookups.scala 95:51]
  wire [26:0] _GEN_36 = io_addr == 6'h1b ? 27'h5a05a05 : _GEN_35; // @[lookups.scala 94:43 lookups.scala 94:51]
  wire [26:0] _GEN_37 = io_addr == 6'h1a ? 27'h5b05b05 : _GEN_36; // @[lookups.scala 93:43 lookups.scala 93:51]
  wire [26:0] _GEN_38 = io_addr == 6'h19 ? 27'h5c0b817 : _GEN_37; // @[lookups.scala 92:43 lookups.scala 92:51]
  wire [26:0] _GEN_39 = io_addr == 6'h18 ? 27'h5d1745d : _GEN_38; // @[lookups.scala 91:43 lookups.scala 91:51]
  wire [26:0] _GEN_40 = io_addr == 6'h17 ? 27'h5e29320 : _GEN_39; // @[lookups.scala 89:43 lookups.scala 89:51]
  wire [26:0] _GEN_41 = io_addr == 6'h16 ? 27'h5f417d0 : _GEN_40; // @[lookups.scala 88:43 lookups.scala 88:51]
  wire [26:0] _GEN_42 = io_addr == 6'h15 ? 27'h6060606 : _GEN_41; // @[lookups.scala 87:43 lookups.scala 87:51]
  wire [26:0] _GEN_43 = io_addr == 6'h14 ? 27'h6186186 : _GEN_42; // @[lookups.scala 86:43 lookups.scala 86:51]
  wire [26:0] _GEN_44 = io_addr == 6'h13 ? 27'h62b2e43 : _GEN_43; // @[lookups.scala 85:43 lookups.scala 85:51]
  wire [26:0] _GEN_45 = io_addr == 6'h12 ? 27'h63e7063 : _GEN_44; // @[lookups.scala 84:43 lookups.scala 84:51]
  wire [26:0] _GEN_46 = io_addr == 6'h11 ? 27'h6522c3f : _GEN_45; // @[lookups.scala 83:43 lookups.scala 83:51]
  wire [26:0] _GEN_47 = io_addr == 6'h10 ? 27'h6666666 : _GEN_46; // @[lookups.scala 82:43 lookups.scala 82:51]
  wire [26:0] _GEN_48 = io_addr == 6'hf ? 27'h67b23a5 : _GEN_47; // @[lookups.scala 80:43 lookups.scala 80:51]
  wire [26:0] _GEN_49 = io_addr == 6'he ? 27'h6906906 : _GEN_48; // @[lookups.scala 79:43 lookups.scala 79:51]
  wire [26:0] _GEN_50 = io_addr == 6'hd ? 27'h6a63bd8 : _GEN_49; // @[lookups.scala 78:43 lookups.scala 78:51]
  wire [26:0] _GEN_51 = io_addr == 6'hc ? 27'h6bca1af : _GEN_50; // @[lookups.scala 77:43 lookups.scala 77:51]
  wire [26:0] _GEN_52 = io_addr == 6'hb ? 27'h6d3a06d : _GEN_51; // @[lookups.scala 76:43 lookups.scala 76:51]
  wire [26:0] _GEN_53 = io_addr == 6'ha ? 27'h6eb3e45 : _GEN_52; // @[lookups.scala 75:43 lookups.scala 75:51]
  wire [26:0] _GEN_54 = io_addr == 6'h9 ? 27'h70381c0 : _GEN_53; // @[lookups.scala 74:43 lookups.scala 74:51]
  wire [26:0] _GEN_55 = io_addr == 6'h8 ? 27'h71c71c7 : _GEN_54; // @[lookups.scala 73:43 lookups.scala 73:51]
  wire [26:0] _GEN_56 = io_addr == 6'h7 ? 27'h73615a2 : _GEN_55; // @[lookups.scala 71:43 lookups.scala 71:51]
  wire [26:0] _GEN_57 = io_addr == 6'h6 ? 27'h7507507 : _GEN_56; // @[lookups.scala 70:43 lookups.scala 70:51]
  wire [26:0] _GEN_58 = io_addr == 6'h5 ? 27'h76b981d : _GEN_57; // @[lookups.scala 69:43 lookups.scala 69:51]
  wire [26:0] _GEN_59 = io_addr == 6'h4 ? 27'h7878787 : _GEN_58; // @[lookups.scala 68:43 lookups.scala 68:51]
  wire [26:0] _GEN_60 = io_addr == 6'h3 ? 27'h7a44c6a : _GEN_59; // @[lookups.scala 67:43 lookups.scala 67:51]
  wire [26:0] _GEN_61 = io_addr == 6'h2 ? 27'h7c1f07c : _GEN_60; // @[lookups.scala 66:43 lookups.scala 66:51]
  wire [26:0] _GEN_62 = io_addr == 6'h1 ? 27'h7e07e07 : _GEN_61; // @[lookups.scala 65:43 lookups.scala 65:51]
  assign io_out = io_addr == 6'h0 ? 27'h0 : _GEN_62; // @[lookups.scala 64:38 lookups.scala 64:46]
endmodule
module lookupJ(
  input  [5:0]  io_addr,
  output [22:0] io_out
);
  wire [15:0] _GEN_0 = io_addr == 6'h3f ? 16'h8205 : 16'h0; // @[lookups.scala 261:43 lookups.scala 261:51 lookups.scala 262:27]
  wire [15:0] _GEN_1 = io_addr == 6'h3e ? 16'h8417 : _GEN_0; // @[lookups.scala 260:43 lookups.scala 260:51]
  wire [15:0] _GEN_2 = io_addr == 6'h3d ? 16'h8636 : _GEN_1; // @[lookups.scala 259:43 lookups.scala 259:51]
  wire [15:0] _GEN_3 = io_addr == 6'h3c ? 16'h8863 : _GEN_2; // @[lookups.scala 258:43 lookups.scala 258:51]
  wire [15:0] _GEN_4 = io_addr == 6'h3b ? 16'h8a9d : _GEN_3; // @[lookups.scala 257:43 lookups.scala 257:51]
  wire [15:0] _GEN_5 = io_addr == 6'h3a ? 16'h8ce5 : _GEN_4; // @[lookups.scala 256:43 lookups.scala 256:51]
  wire [15:0] _GEN_6 = io_addr == 6'h39 ? 16'h8f3b : _GEN_5; // @[lookups.scala 255:43 lookups.scala 255:51]
  wire [15:0] _GEN_7 = io_addr == 6'h38 ? 16'h91a1 : _GEN_6; // @[lookups.scala 254:43 lookups.scala 254:51]
  wire [15:0] _GEN_8 = io_addr == 6'h37 ? 16'h9416 : _GEN_7; // @[lookups.scala 252:43 lookups.scala 252:51]
  wire [15:0] _GEN_9 = io_addr == 6'h36 ? 16'h969b : _GEN_8; // @[lookups.scala 251:43 lookups.scala 251:51]
  wire [15:0] _GEN_10 = io_addr == 6'h35 ? 16'h9931 : _GEN_9; // @[lookups.scala 250:43 lookups.scala 250:51]
  wire [15:0] _GEN_11 = io_addr == 6'h34 ? 16'h9bd8 : _GEN_10; // @[lookups.scala 249:43 lookups.scala 249:51]
  wire [15:0] _GEN_12 = io_addr == 6'h33 ? 16'h9e91 : _GEN_11; // @[lookups.scala 248:43 lookups.scala 248:51]
  wire [15:0] _GEN_13 = io_addr == 6'h32 ? 16'ha15c : _GEN_12; // @[lookups.scala 247:43 lookups.scala 247:51]
  wire [15:0] _GEN_14 = io_addr == 6'h31 ? 16'ha43b : _GEN_13; // @[lookups.scala 246:43 lookups.scala 246:51]
  wire [15:0] _GEN_15 = io_addr == 6'h30 ? 16'ha72d : _GEN_14; // @[lookups.scala 245:43 lookups.scala 245:51]
  wire [15:0] _GEN_16 = io_addr == 6'h2f ? 16'haa33 : _GEN_15; // @[lookups.scala 243:43 lookups.scala 243:51]
  wire [15:0] _GEN_17 = io_addr == 6'h2e ? 16'had4f : _GEN_16; // @[lookups.scala 242:43 lookups.scala 242:51]
  wire [15:0] _GEN_18 = io_addr == 6'h2d ? 16'hb081 : _GEN_17; // @[lookups.scala 241:43 lookups.scala 241:51]
  wire [15:0] _GEN_19 = io_addr == 6'h2c ? 16'hb3ca : _GEN_18; // @[lookups.scala 240:43 lookups.scala 240:51]
  wire [15:0] _GEN_20 = io_addr == 6'h2b ? 16'hb72a : _GEN_19; // @[lookups.scala 239:43 lookups.scala 239:51]
  wire [15:0] _GEN_21 = io_addr == 6'h2a ? 16'hbaa3 : _GEN_20; // @[lookups.scala 238:43 lookups.scala 238:51]
  wire [15:0] _GEN_22 = io_addr == 6'h29 ? 16'hbe35 : _GEN_21; // @[lookups.scala 237:43 lookups.scala 237:51]
  wire [15:0] _GEN_23 = io_addr == 6'h28 ? 16'hc1e2 : _GEN_22; // @[lookups.scala 236:43 lookups.scala 236:51]
  wire [15:0] _GEN_24 = io_addr == 6'h27 ? 16'hc5aa : _GEN_23; // @[lookups.scala 234:43 lookups.scala 234:51]
  wire [15:0] _GEN_25 = io_addr == 6'h26 ? 16'hc98f : _GEN_24; // @[lookups.scala 233:43 lookups.scala 233:51]
  wire [15:0] _GEN_26 = io_addr == 6'h25 ? 16'hcd92 : _GEN_25; // @[lookups.scala 232:43 lookups.scala 232:51]
  wire [15:0] _GEN_27 = io_addr == 6'h24 ? 16'hd1b4 : _GEN_26; // @[lookups.scala 231:43 lookups.scala 231:51]
  wire [15:0] _GEN_28 = io_addr == 6'h23 ? 16'hd5f6 : _GEN_27; // @[lookups.scala 230:43 lookups.scala 230:51]
  wire [15:0] _GEN_29 = io_addr == 6'h22 ? 16'hda59 : _GEN_28; // @[lookups.scala 229:43 lookups.scala 229:51]
  wire [15:0] _GEN_30 = io_addr == 6'h21 ? 16'hdee0 : _GEN_29; // @[lookups.scala 228:43 lookups.scala 228:51]
  wire [15:0] _GEN_31 = io_addr == 6'h20 ? 16'he38b : _GEN_30; // @[lookups.scala 227:43 lookups.scala 227:51]
  wire [15:0] _GEN_32 = io_addr == 6'h1f ? 16'he85b : _GEN_31; // @[lookups.scala 225:43 lookups.scala 225:51]
  wire [15:0] _GEN_33 = io_addr == 6'h1e ? 16'hed54 : _GEN_32; // @[lookups.scala 224:43 lookups.scala 224:51]
  wire [15:0] _GEN_34 = io_addr == 6'h1d ? 16'hf275 : _GEN_33; // @[lookups.scala 223:43 lookups.scala 223:51]
  wire [15:0] _GEN_35 = io_addr == 6'h1c ? 16'hf7c2 : _GEN_34; // @[lookups.scala 222:43 lookups.scala 222:51]
  wire [15:0] _GEN_36 = io_addr == 6'h1b ? 16'hfd3b : _GEN_35; // @[lookups.scala 221:43 lookups.scala 221:51]
  wire [16:0] _GEN_37 = io_addr == 6'h1a ? 17'h102e4 : {{1'd0}, _GEN_36}; // @[lookups.scala 220:43 lookups.scala 220:51]
  wire [16:0] _GEN_38 = io_addr == 6'h19 ? 17'h108bd : _GEN_37; // @[lookups.scala 219:43 lookups.scala 219:51]
  wire [16:0] _GEN_39 = io_addr == 6'h18 ? 17'h10eca : _GEN_38; // @[lookups.scala 218:43 lookups.scala 218:51]
  wire [16:0] _GEN_40 = io_addr == 6'h17 ? 17'h1150d : _GEN_39; // @[lookups.scala 216:43 lookups.scala 216:51]
  wire [16:0] _GEN_41 = io_addr == 6'h16 ? 17'h11b88 : _GEN_40; // @[lookups.scala 215:43 lookups.scala 215:51]
  wire [16:0] _GEN_42 = io_addr == 6'h15 ? 17'h1223e : _GEN_41; // @[lookups.scala 214:43 lookups.scala 214:51]
  wire [16:0] _GEN_43 = io_addr == 6'h14 ? 17'h12931 : _GEN_42; // @[lookups.scala 213:43 lookups.scala 213:51]
  wire [16:0] _GEN_44 = io_addr == 6'h13 ? 17'h13066 : _GEN_43; // @[lookups.scala 212:43 lookups.scala 212:51]
  wire [16:0] _GEN_45 = io_addr == 6'h12 ? 17'h137de : _GEN_44; // @[lookups.scala 211:43 lookups.scala 211:51]
  wire [16:0] _GEN_46 = io_addr == 6'h11 ? 17'h13f9d : _GEN_45; // @[lookups.scala 210:43 lookups.scala 210:51]
  wire [16:0] _GEN_47 = io_addr == 6'h10 ? 17'h147a7 : _GEN_46; // @[lookups.scala 209:43 lookups.scala 209:51]
  wire [16:0] _GEN_48 = io_addr == 6'hf ? 17'h15000 : _GEN_47; // @[lookups.scala 207:43 lookups.scala 207:51]
  wire [16:0] _GEN_49 = io_addr == 6'he ? 17'h158ab : _GEN_48; // @[lookups.scala 206:43 lookups.scala 206:51]
  wire [16:0] _GEN_50 = io_addr == 6'hd ? 17'h161ae : _GEN_49; // @[lookups.scala 205:43 lookups.scala 205:51]
  wire [16:0] _GEN_51 = io_addr == 6'hc ? 17'h16b0c : _GEN_50; // @[lookups.scala 204:43 lookups.scala 204:51]
  wire [16:0] _GEN_52 = io_addr == 6'hb ? 17'h174cb : _GEN_51; // @[lookups.scala 203:43 lookups.scala 203:51]
  wire [16:0] _GEN_53 = io_addr == 6'ha ? 17'h17eef : _GEN_52; // @[lookups.scala 202:43 lookups.scala 202:51]
  wire [16:0] _GEN_54 = io_addr == 6'h9 ? 17'h1897f : _GEN_53; // @[lookups.scala 201:43 lookups.scala 201:51]
  wire [16:0] _GEN_55 = io_addr == 6'h8 ? 17'h19481 : _GEN_54; // @[lookups.scala 200:43 lookups.scala 200:51]
  wire [16:0] _GEN_56 = io_addr == 6'h7 ? 17'h19ffa : _GEN_55; // @[lookups.scala 198:43 lookups.scala 198:51]
  wire [16:0] _GEN_57 = io_addr == 6'h6 ? 17'h1abf2 : _GEN_56; // @[lookups.scala 197:43 lookups.scala 197:51]
  wire [16:0] _GEN_58 = io_addr == 6'h5 ? 17'h1b870 : _GEN_57; // @[lookups.scala 196:43 lookups.scala 196:51]
  wire [16:0] _GEN_59 = io_addr == 6'h4 ? 17'h1c57d : _GEN_58; // @[lookups.scala 195:43 lookups.scala 195:51]
  wire [16:0] _GEN_60 = io_addr == 6'h3 ? 17'h1d31f : _GEN_59; // @[lookups.scala 194:43 lookups.scala 194:51]
  wire [16:0] _GEN_61 = io_addr == 6'h2 ? 17'h1e162 : _GEN_60; // @[lookups.scala 193:43 lookups.scala 193:51]
  wire [16:0] _GEN_62 = io_addr == 6'h1 ? 17'h1f04f : _GEN_61; // @[lookups.scala 192:43 lookups.scala 192:51]
  wire [16:0] _GEN_63 = io_addr == 6'h0 ? 17'h1fff0 : _GEN_62; // @[lookups.scala 191:38 lookups.scala 191:46]
  assign io_out = {{6'd0}, _GEN_63}; // @[lookups.scala 191:38 lookups.scala 191:46]
endmodule
module VarSizeMul(
  input  [22:0] io_in1,
  input  [16:0] io_in2,
  output [23:0] io_out
);
  wire [22:0] _GEN_0 = {{6'd0}, io_in2}; // @[VarSizeMul.scala 20:26]
  wire [39:0] result = io_in1 * _GEN_0; // @[VarSizeMul.scala 20:26]
  assign io_out = result[39:16]; // @[VarSizeMul.scala 22:25]
endmodule
module mul2(
  input  [23:0] io_in1,
  input  [16:0] io_in2,
  output [28:0] io_out
);
  wire [23:0] _GEN_0 = {{7'd0}, io_in2}; // @[VarSizeMul.scala 37:26]
  wire [40:0] result = io_in1 * _GEN_0; // @[VarSizeMul.scala 37:26]
  assign io_out = result[40:12]; // @[VarSizeMul.scala 38:25]
endmodule
module VarSizeSub(
  input  [26:0] io_in1,
  input  [26:0] io_in2,
  output [26:0] io_out
);
  assign io_out = io_in1 + io_in2; // @[VarSizeAdder.scala 36:27]
endmodule
module VarSizeAdder(
  input  [28:0] io_in1,
  input  [28:0] io_in2,
  output [24:0] io_out
);
  wire [28:0] _T_1 = io_in1 + io_in2; // @[VarSizeAdder.scala 21:27]
  assign io_out = _T_1[28:4]; // @[VarSizeAdder.scala 21:36]
endmodule
module mul3(
  input  [22:0] io_in1,
  input  [24:0] io_in2,
  output [23:0] io_out
);
  wire [24:0] _GEN_0 = {{2'd0}, io_in1}; // @[VarSizeMul.scala 54:26]
  wire [47:0] result = _GEN_0 * io_in2; // @[VarSizeMul.scala 54:26]
  assign io_out = result[47:24]; // @[VarSizeMul.scala 55:25]
endmodule
module fpInverter(
  input         clock,
  input         reset,
  input  [22:0] io_in1,
  output [23:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire [5:0] tableC_io_addr; // @[fpInverter.scala 19:28]
  wire [23:0] tableC_io_out; // @[fpInverter.scala 19:28]
  wire [5:0] tableL_io_addr; // @[fpInverter.scala 20:28]
  wire [26:0] tableL_io_out; // @[fpInverter.scala 20:28]
  wire [5:0] tableJ_io_addr; // @[fpInverter.scala 21:28]
  wire [22:0] tableJ_io_out; // @[fpInverter.scala 21:28]
  wire [22:0] mul1_io_in1; // @[fpInverter.scala 32:26]
  wire [16:0] mul1_io_in2; // @[fpInverter.scala 32:26]
  wire [23:0] mul1_io_out; // @[fpInverter.scala 32:26]
  wire [23:0] mul2_io_in1; // @[fpInverter.scala 37:26]
  wire [16:0] mul2_io_in2; // @[fpInverter.scala 37:26]
  wire [28:0] mul2_io_out; // @[fpInverter.scala 37:26]
  wire [26:0] sub2_io_in1; // @[fpInverter.scala 65:30]
  wire [26:0] sub2_io_in2; // @[fpInverter.scala 65:30]
  wire [26:0] sub2_io_out; // @[fpInverter.scala 65:30]
  wire [28:0] adder_io_in1; // @[fpInverter.scala 74:31]
  wire [28:0] adder_io_in2; // @[fpInverter.scala 74:31]
  wire [24:0] adder_io_out; // @[fpInverter.scala 74:31]
  wire [22:0] mul3_io_in1; // @[fpInverter.scala 89:30]
  wire [24:0] mul3_io_in2; // @[fpInverter.scala 89:30]
  wire [23:0] mul3_io_out; // @[fpInverter.scala 89:30]
  wire [22:0] _T = io_in1 ^ 23'h7fffff; // @[fpInverter.scala 30:28]
  wire [33:0] _T_5 = io_in1[16:0] * io_in1[16:0]; // @[fpInverter.scala 39:42]
  reg [22:0] w_sub1_reg; // @[fpInverter.scala 43:41]
  reg [23:0] w_mul1_reg; // @[fpInverter.scala 44:41]
  reg [28:0] w_mul2_reg; // @[fpInverter.scala 45:41]
  reg [26:0] tableL_out_reg; // @[fpInverter.scala 57:37]
  reg [22:0] sub1_out_reg1; // @[fpInverter.scala 59:37]
  reg [23:0] mul1_out_reg; // @[fpInverter.scala 60:37]
  reg [28:0] mul2_out_reg; // @[fpInverter.scala 61:37]
  wire [23:0] _T_7 = mul1_out_reg ^ 24'hffffff; // @[fpInverter.scala 66:38]
  wire [23:0] sub2_in2 = _T_7 + 24'h1; // @[fpInverter.scala 66:71]
  wire [25:0] temp4 = {sub2_in2,1'h0,1'h0}; // @[Cat.scala 30:58]
  wire [27:0] temp1 = {sub2_io_out,1'h0}; // @[Cat.scala 30:58]
  reg [22:0] sub1_out_reg2; // @[fpInverter.scala 82:36]
  reg [24:0] adder_out_reg; // @[fpInverter.scala 85:36]
  reg [24:0] adder_out_reg_2; // @[fpInverter.scala 87:38]
  lookupC tableC ( // @[fpInverter.scala 19:28]
    .io_addr(tableC_io_addr),
    .io_out(tableC_io_out)
  );
  lookupL tableL ( // @[fpInverter.scala 20:28]
    .io_addr(tableL_io_addr),
    .io_out(tableL_io_out)
  );
  lookupJ tableJ ( // @[fpInverter.scala 21:28]
    .io_addr(tableJ_io_addr),
    .io_out(tableJ_io_out)
  );
  VarSizeMul mul1 ( // @[fpInverter.scala 32:26]
    .io_in1(mul1_io_in1),
    .io_in2(mul1_io_in2),
    .io_out(mul1_io_out)
  );
  mul2 mul2 ( // @[fpInverter.scala 37:26]
    .io_in1(mul2_io_in1),
    .io_in2(mul2_io_in2),
    .io_out(mul2_io_out)
  );
  VarSizeSub sub2 ( // @[fpInverter.scala 65:30]
    .io_in1(sub2_io_in1),
    .io_in2(sub2_io_in2),
    .io_out(sub2_io_out)
  );
  VarSizeAdder adder ( // @[fpInverter.scala 74:31]
    .io_in1(adder_io_in1),
    .io_in2(adder_io_in2),
    .io_out(adder_io_out)
  );
  mul3 mul3 ( // @[fpInverter.scala 89:30]
    .io_in1(mul3_io_in1),
    .io_in2(mul3_io_in2),
    .io_out(mul3_io_out)
  );
  assign io_out = mul3_io_out; // @[fpInverter.scala 97:16]
  assign tableC_io_addr = io_in1[22:17]; // @[fpInverter.scala 25:33]
  assign tableL_io_addr = io_in1[22:17]; // @[fpInverter.scala 25:33]
  assign tableJ_io_addr = io_in1[22:17]; // @[fpInverter.scala 25:33]
  assign mul1_io_in1 = tableJ_io_out; // @[fpInverter.scala 33:21]
  assign mul1_io_in2 = io_in1[16:0]; // @[fpInverter.scala 34:30]
  assign mul2_io_in1 = tableC_io_out; // @[fpInverter.scala 38:21]
  assign mul2_io_in2 = _T_5[33:17]; // @[fpInverter.scala 39:61]
  assign sub2_io_in1 = tableL_out_reg; // @[fpInverter.scala 70:21]
  assign sub2_io_in2 = {temp4,1'h0}; // @[Cat.scala 30:58]
  assign adder_io_in1 = {temp1,1'h0}; // @[Cat.scala 30:58]
  assign adder_io_in2 = mul2_out_reg; // @[fpInverter.scala 78:22]
  assign mul3_io_in1 = sub1_out_reg2; // @[fpInverter.scala 91:21]
  assign mul3_io_in2 = adder_out_reg_2; // @[fpInverter.scala 92:21]
  always @(posedge clock) begin
    w_sub1_reg <= _T + 23'h1; // @[fpInverter.scala 30:60]
    w_mul1_reg <= mul1_io_out; // @[fpInverter.scala 44:41]
    w_mul2_reg <= mul2_io_out; // @[fpInverter.scala 45:41]
    tableL_out_reg <= tableL_io_out; // @[fpInverter.scala 57:37]
    sub1_out_reg1 <= w_sub1_reg; // @[fpInverter.scala 59:37]
    mul1_out_reg <= w_mul1_reg; // @[fpInverter.scala 60:37]
    mul2_out_reg <= w_mul2_reg; // @[fpInverter.scala 61:37]
    sub1_out_reg2 <= sub1_out_reg1; // @[fpInverter.scala 82:36]
    if (reset) begin // @[fpInverter.scala 85:36]
      adder_out_reg <= 25'h0; // @[fpInverter.scala 85:36]
    end else begin
      adder_out_reg <= adder_io_out; // @[fpInverter.scala 86:25]
    end
    if (reset) begin // @[fpInverter.scala 87:38]
      adder_out_reg_2 <= 25'h0; // @[fpInverter.scala 87:38]
    end else begin
      adder_out_reg_2 <= adder_out_reg; // @[fpInverter.scala 88:25]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  w_sub1_reg = _RAND_0[22:0];
  _RAND_1 = {1{`RANDOM}};
  w_mul1_reg = _RAND_1[23:0];
  _RAND_2 = {1{`RANDOM}};
  w_mul2_reg = _RAND_2[28:0];
  _RAND_3 = {1{`RANDOM}};
  tableL_out_reg = _RAND_3[26:0];
  _RAND_4 = {1{`RANDOM}};
  sub1_out_reg1 = _RAND_4[22:0];
  _RAND_5 = {1{`RANDOM}};
  mul1_out_reg = _RAND_5[23:0];
  _RAND_6 = {1{`RANDOM}};
  mul2_out_reg = _RAND_6[28:0];
  _RAND_7 = {1{`RANDOM}};
  sub1_out_reg2 = _RAND_7[22:0];
  _RAND_8 = {1{`RANDOM}};
  adder_out_reg = _RAND_8[24:0];
  _RAND_9 = {1{`RANDOM}};
  adder_out_reg_2 = _RAND_9[24:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module fp_inverter(
  input         clock,
  input         reset,
  input  [31:0] io_in1,
  output [31:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire  inverter_clock; // @[FP_inverter.scala 14:29]
  wire  inverter_reset; // @[FP_inverter.scala 14:29]
  wire [22:0] inverter_io_in1; // @[FP_inverter.scala 14:29]
  wire [23:0] inverter_io_out; // @[FP_inverter.scala 14:29]
  reg [7:0] in2ExpReg0; // @[FP_inverter.scala 18:42]
  reg  in2SignReg0; // @[FP_inverter.scala 20:42]
  reg [7:0] in2ExpReg1; // @[FP_inverter.scala 22:35]
  reg  in2SignReg1; // @[FP_inverter.scala 24:42]
  reg [7:0] in2ExpReg2; // @[FP_inverter.scala 27:35]
  reg  in2SignReg2; // @[FP_inverter.scala 29:42]
  reg [7:0] in2ExpReg3; // @[FP_inverter.scala 32:35]
  reg  in2SignReg3; // @[FP_inverter.scala 34:42]
  reg [23:0] invMant; // @[FP_inverter.scala 37:42]
  wire [23:0] _T_3 = inverter_io_out; // @[FP_inverter.scala 38:67]
  wire [7:0] negExpTmp = 8'hfe - in2ExpReg3; // @[FP_inverter.scala 41:35]
  wire [7:0] _T_7 = negExpTmp - 8'h1; // @[FP_inverter.scala 42:71]
  wire [7:0] negExp = invMant == 24'h0 ? negExpTmp : _T_7; // @[FP_inverter.scala 42:32]
  wire [22:0] lo = invMant[23:1]; // @[FP_inverter.scala 43:77]
  wire [8:0] hi = {in2SignReg3,negExp}; // @[Cat.scala 30:58]
  fpInverter inverter ( // @[FP_inverter.scala 14:29]
    .clock(inverter_clock),
    .reset(inverter_reset),
    .io_in1(inverter_io_in1),
    .io_out(inverter_io_out)
  );
  assign io_out = {hi,lo}; // @[Cat.scala 30:58]
  assign inverter_clock = clock;
  assign inverter_reset = reset;
  assign inverter_io_in1 = io_in1[22:0]; // @[FP_inverter.scala 16:30]
  always @(posedge clock) begin
    if (reset) begin // @[FP_inverter.scala 18:42]
      in2ExpReg0 <= 8'h0; // @[FP_inverter.scala 18:42]
    end else begin
      in2ExpReg0 <= io_in1[30:23]; // @[FP_inverter.scala 19:44]
    end
    if (reset) begin // @[FP_inverter.scala 20:42]
      in2SignReg0 <= 1'h0; // @[FP_inverter.scala 20:42]
    end else begin
      in2SignReg0 <= io_in1[31]; // @[FP_inverter.scala 21:43]
    end
    if (reset) begin // @[FP_inverter.scala 22:35]
      in2ExpReg1 <= 8'h0; // @[FP_inverter.scala 22:35]
    end else begin
      in2ExpReg1 <= in2ExpReg0; // @[FP_inverter.scala 23:43]
    end
    if (reset) begin // @[FP_inverter.scala 24:42]
      in2SignReg1 <= 1'h0; // @[FP_inverter.scala 24:42]
    end else begin
      in2SignReg1 <= in2SignReg0; // @[FP_inverter.scala 25:43]
    end
    if (reset) begin // @[FP_inverter.scala 27:35]
      in2ExpReg2 <= 8'h0; // @[FP_inverter.scala 27:35]
    end else begin
      in2ExpReg2 <= in2ExpReg1; // @[FP_inverter.scala 28:43]
    end
    if (reset) begin // @[FP_inverter.scala 29:42]
      in2SignReg2 <= 1'h0; // @[FP_inverter.scala 29:42]
    end else begin
      in2SignReg2 <= in2SignReg1; // @[FP_inverter.scala 30:43]
    end
    if (reset) begin // @[FP_inverter.scala 32:35]
      in2ExpReg3 <= 8'h0; // @[FP_inverter.scala 32:35]
    end else begin
      in2ExpReg3 <= in2ExpReg2; // @[FP_inverter.scala 33:43]
    end
    if (reset) begin // @[FP_inverter.scala 34:42]
      in2SignReg3 <= 1'h0; // @[FP_inverter.scala 34:42]
    end else begin
      in2SignReg3 <= in2SignReg2; // @[FP_inverter.scala 35:43]
    end
    if (reset) begin // @[FP_inverter.scala 37:42]
      invMant <= 24'h0; // @[FP_inverter.scala 37:42]
    end else begin
      invMant <= _T_3; // @[FP_inverter.scala 38:49]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  in2ExpReg0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  in2SignReg0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  in2ExpReg1 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  in2SignReg1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  in2ExpReg2 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  in2SignReg2 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  in2ExpReg3 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  in2SignReg3 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  invMant = _RAND_8[23:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Schedule_unit(
  input         clock,
  input         reset,
  input  [31:0] io_invDz_div,
  input         io_valid_in,
  input  [31:0] io_v11_x,
  input  [31:0] io_v11_y,
  input  [31:0] io_v11_z,
  input  [31:0] io_v11_w,
  input  [31:0] io_v22_x,
  input  [31:0] io_v22_y,
  input  [31:0] io_v22_z,
  input  [31:0] io_v22_w,
  input  [31:0] io_ray_in,
  input  [31:0] io_Oz,
  input  [31:0] io_ray_o_in_x,
  input  [31:0] io_ray_o_in_y,
  input  [31:0] io_ray_o_in_z,
  input  [31:0] io_ray_d_in_x,
  input  [31:0] io_ray_d_in_y,
  input  [31:0] io_ray_d_in_z,
  input  [31:0] io_node_id_in,
  input  [31:0] io_hitT_in,
  input         io_break_in,
  input         io_RAY_AABB_1,
  input         io_RAY_AABB_2,
  output [31:0] io_fdiv_out,
  output        io_valid_out,
  output [31:0] io_v11_out_x,
  output [31:0] io_v11_out_y,
  output [31:0] io_v11_out_z,
  output [31:0] io_v11_out_w,
  output [31:0] io_v22_out_x,
  output [31:0] io_v22_out_y,
  output [31:0] io_v22_out_z,
  output [31:0] io_v22_out_w,
  output [31:0] io_ray_out,
  output [31:0] io_Oz_out,
  output [31:0] io_ray_o_out_x,
  output [31:0] io_ray_o_out_y,
  output [31:0] io_ray_o_out_z,
  output [31:0] io_ray_d_out_x,
  output [31:0] io_ray_d_out_y,
  output [31:0] io_ray_d_out_z,
  output [31:0] io_node_id_out,
  output [31:0] io_hitT_out,
  output [31:0] io_counter_fdiv,
  output        io_break_out,
  output        io_RAY_AABB_1_out,
  output        io_RAY_AABB_2_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [95:0] _RAND_4;
  reg [95:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [127:0] _RAND_12;
  reg [127:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [95:0] _RAND_16;
  reg [95:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [127:0] _RAND_24;
  reg [127:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [95:0] _RAND_28;
  reg [95:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [127:0] _RAND_36;
  reg [127:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [95:0] _RAND_40;
  reg [95:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [63:0] _RAND_48;
`endif // RANDOMIZE_REG_INIT
  wire  FP_inverter_clock; // @[Schedule_unit_1.scala 39:39]
  wire  FP_inverter_reset; // @[Schedule_unit_1.scala 39:39]
  wire [31:0] FP_inverter_io_in1; // @[Schedule_unit_1.scala 39:39]
  wire [31:0] FP_inverter_io_out; // @[Schedule_unit_1.scala 39:39]
  reg [127:0] v11_temp_1; // @[Schedule_unit_1.scala 44:38]
  reg [127:0] v22_temp_1; // @[Schedule_unit_1.scala 45:42]
  reg [31:0] ray_temp_1; // @[Schedule_unit_1.scala 46:43]
  reg [31:0] Oz_temp_1; // @[Schedule_unit_1.scala 47:43]
  reg [95:0] ray_o_temp_1; // @[Schedule_unit_1.scala 48:40]
  reg [95:0] ray_d_temp_1; // @[Schedule_unit_1.scala 49:40]
  reg [31:0] node_id_temp_1; // @[Schedule_unit_1.scala 50:37]
  reg [31:0] hitT_temp_1; // @[Schedule_unit_1.scala 51:43]
  reg  inValid_1; // @[Schedule_unit_1.scala 52:61]
  reg  break_1; // @[Schedule_unit_1.scala 53:45]
  reg  ray_aabb_1; // @[Schedule_unit_1.scala 54:46]
  reg  ray_aabb_2; // @[Schedule_unit_1.scala 55:46]
  wire [127:0] _T = {io_v11_w,io_v11_z,io_v11_y,io_v11_x}; // @[Cat.scala 30:58]
  wire [127:0] _T_1 = {io_v22_w,io_v22_z,io_v22_y,io_v22_x}; // @[Cat.scala 30:58]
  wire [95:0] _T_2 = {io_ray_o_in_z,io_ray_o_in_y,io_ray_o_in_x}; // @[Cat.scala 30:58]
  wire [95:0] _T_3 = {io_ray_d_in_z,io_ray_d_in_y,io_ray_d_in_x}; // @[Cat.scala 30:58]
  reg [127:0] v11_temp_2; // @[Schedule_unit_1.scala 70:42]
  reg [127:0] v22_temp_2; // @[Schedule_unit_1.scala 71:42]
  reg [31:0] ray_temp_2; // @[Schedule_unit_1.scala 72:43]
  reg [31:0] Oz_temp_2; // @[Schedule_unit_1.scala 73:43]
  reg [95:0] ray_o_temp_2; // @[Schedule_unit_1.scala 74:40]
  reg [95:0] ray_d_temp_2; // @[Schedule_unit_1.scala 75:40]
  reg [31:0] node_id_temp_2; // @[Schedule_unit_1.scala 76:37]
  reg [31:0] hitT_temp_2; // @[Schedule_unit_1.scala 77:43]
  reg  inValid_2; // @[Schedule_unit_1.scala 78:61]
  reg  break_2; // @[Schedule_unit_1.scala 79:45]
  reg  ray_aabb_1_2; // @[Schedule_unit_1.scala 80:43]
  reg  ray_aabb_2_2; // @[Schedule_unit_1.scala 81:43]
  reg [127:0] v11_temp_3; // @[Schedule_unit_1.scala 96:42]
  reg [127:0] v22_temp_3; // @[Schedule_unit_1.scala 97:42]
  reg [31:0] ray_temp_3; // @[Schedule_unit_1.scala 98:43]
  reg [31:0] Oz_temp_3; // @[Schedule_unit_1.scala 99:43]
  reg [95:0] ray_o_temp_3; // @[Schedule_unit_1.scala 100:40]
  reg [95:0] ray_d_temp_3; // @[Schedule_unit_1.scala 101:40]
  reg [31:0] node_id_temp_3; // @[Schedule_unit_1.scala 102:37]
  reg [31:0] hitT_temp_3; // @[Schedule_unit_1.scala 103:43]
  reg  inValid_3; // @[Schedule_unit_1.scala 104:61]
  reg  break_3; // @[Schedule_unit_1.scala 105:45]
  reg  ray_aabb_1_3; // @[Schedule_unit_1.scala 106:43]
  reg  ray_aabb_2_3; // @[Schedule_unit_1.scala 107:43]
  reg [127:0] v11_temp_4; // @[Schedule_unit_1.scala 121:38]
  reg [127:0] v22_temp_4; // @[Schedule_unit_1.scala 122:42]
  reg [31:0] ray_temp_4; // @[Schedule_unit_1.scala 123:43]
  reg [31:0] Oz_temp_4; // @[Schedule_unit_1.scala 124:43]
  reg [95:0] ray_o_temp_4; // @[Schedule_unit_1.scala 125:40]
  reg [95:0] ray_d_temp_4; // @[Schedule_unit_1.scala 126:40]
  reg [31:0] node_id_temp_4; // @[Schedule_unit_1.scala 127:37]
  reg [31:0] hitT_temp_4; // @[Schedule_unit_1.scala 128:43]
  reg  inValid_4; // @[Schedule_unit_1.scala 129:61]
  reg  break_4; // @[Schedule_unit_1.scala 130:45]
  reg  ray_aabb_1_4; // @[Schedule_unit_1.scala 131:43]
  reg  ray_aabb_2_4; // @[Schedule_unit_1.scala 132:43]
  reg [63:0] count; // @[Schedule_unit_1.scala 171:46]
  wire [63:0] _T_19 = count + 64'h1; // @[Schedule_unit_1.scala 191:26]
  fp_inverter FP_inverter ( // @[Schedule_unit_1.scala 39:39]
    .clock(FP_inverter_clock),
    .reset(FP_inverter_reset),
    .io_in1(FP_inverter_io_in1),
    .io_out(FP_inverter_io_out)
  );
  assign io_fdiv_out = FP_inverter_io_out; // @[Schedule_unit_1.scala 42:45]
  assign io_valid_out = inValid_4; // @[Schedule_unit_1.scala 147:65]
  assign io_v11_out_x = v11_temp_4[31:0]; // @[Schedule_unit_1.scala 148:61]
  assign io_v11_out_y = v11_temp_4[63:32]; // @[Schedule_unit_1.scala 149:61]
  assign io_v11_out_z = v11_temp_4[95:64]; // @[Schedule_unit_1.scala 150:61]
  assign io_v11_out_w = v11_temp_4[127:96]; // @[Schedule_unit_1.scala 151:60]
  assign io_v22_out_x = v22_temp_4[31:0]; // @[Schedule_unit_1.scala 152:61]
  assign io_v22_out_y = v22_temp_4[63:32]; // @[Schedule_unit_1.scala 153:61]
  assign io_v22_out_z = v22_temp_4[95:64]; // @[Schedule_unit_1.scala 154:61]
  assign io_v22_out_w = v22_temp_4[127:96]; // @[Schedule_unit_1.scala 155:59]
  assign io_ray_out = ray_temp_4; // @[Schedule_unit_1.scala 157:50]
  assign io_Oz_out = Oz_temp_4; // @[Schedule_unit_1.scala 158:50]
  assign io_ray_o_out_x = ray_o_temp_4[31:0]; // @[Schedule_unit_1.scala 159:60]
  assign io_ray_o_out_y = ray_o_temp_4[63:32]; // @[Schedule_unit_1.scala 160:60]
  assign io_ray_o_out_z = ray_o_temp_4[95:64]; // @[Schedule_unit_1.scala 161:60]
  assign io_ray_d_out_x = ray_d_temp_4[31:0]; // @[Schedule_unit_1.scala 162:60]
  assign io_ray_d_out_y = ray_d_temp_4[63:32]; // @[Schedule_unit_1.scala 163:60]
  assign io_ray_d_out_z = ray_d_temp_4[95:64]; // @[Schedule_unit_1.scala 164:60]
  assign io_node_id_out = node_id_temp_4; // @[Schedule_unit_1.scala 165:59]
  assign io_hitT_out = hitT_temp_4; // @[Schedule_unit_1.scala 166:73]
  assign io_counter_fdiv = count[31:0]; // @[Schedule_unit_1.scala 196:21]
  assign io_break_out = break_4; // @[Schedule_unit_1.scala 167:42]
  assign io_RAY_AABB_1_out = ray_aabb_1_4; // @[Schedule_unit_1.scala 168:33]
  assign io_RAY_AABB_2_out = ray_aabb_2_4; // @[Schedule_unit_1.scala 169:33]
  assign FP_inverter_clock = clock;
  assign FP_inverter_reset = reset;
  assign FP_inverter_io_in1 = io_invDz_div; // @[Schedule_unit_1.scala 41:37]
  always @(posedge clock) begin
    if (reset) begin // @[Schedule_unit_1.scala 44:38]
      v11_temp_1 <= 128'h0; // @[Schedule_unit_1.scala 44:38]
    end else begin
      v11_temp_1 <= _T; // @[Schedule_unit_1.scala 57:48]
    end
    if (reset) begin // @[Schedule_unit_1.scala 45:42]
      v22_temp_1 <= 128'h0; // @[Schedule_unit_1.scala 45:42]
    end else begin
      v22_temp_1 <= _T_1; // @[Schedule_unit_1.scala 58:48]
    end
    if (reset) begin // @[Schedule_unit_1.scala 46:43]
      ray_temp_1 <= 32'h0; // @[Schedule_unit_1.scala 46:43]
    end else begin
      ray_temp_1 <= io_ray_in; // @[Schedule_unit_1.scala 59:49]
    end
    if (reset) begin // @[Schedule_unit_1.scala 47:43]
      Oz_temp_1 <= 32'h0; // @[Schedule_unit_1.scala 47:43]
    end else begin
      Oz_temp_1 <= io_Oz; // @[Schedule_unit_1.scala 60:49]
    end
    if (reset) begin // @[Schedule_unit_1.scala 48:40]
      ray_o_temp_1 <= 96'h0; // @[Schedule_unit_1.scala 48:40]
    end else begin
      ray_o_temp_1 <= _T_2; // @[Schedule_unit_1.scala 61:46]
    end
    if (reset) begin // @[Schedule_unit_1.scala 49:40]
      ray_d_temp_1 <= 96'h0; // @[Schedule_unit_1.scala 49:40]
    end else begin
      ray_d_temp_1 <= _T_3; // @[Schedule_unit_1.scala 62:46]
    end
    if (reset) begin // @[Schedule_unit_1.scala 50:37]
      node_id_temp_1 <= 32'sh0; // @[Schedule_unit_1.scala 50:37]
    end else begin
      node_id_temp_1 <= io_node_id_in; // @[Schedule_unit_1.scala 63:43]
    end
    if (reset) begin // @[Schedule_unit_1.scala 51:43]
      hitT_temp_1 <= 32'h0; // @[Schedule_unit_1.scala 51:43]
    end else begin
      hitT_temp_1 <= io_hitT_in; // @[Schedule_unit_1.scala 64:49]
    end
    if (reset) begin // @[Schedule_unit_1.scala 52:61]
      inValid_1 <= 1'h0; // @[Schedule_unit_1.scala 52:61]
    end else begin
      inValid_1 <= io_valid_in; // @[Schedule_unit_1.scala 65:50]
    end
    if (reset) begin // @[Schedule_unit_1.scala 53:45]
      break_1 <= 1'h0; // @[Schedule_unit_1.scala 53:45]
    end else begin
      break_1 <= io_break_in; // @[Schedule_unit_1.scala 66:51]
    end
    if (reset) begin // @[Schedule_unit_1.scala 54:46]
      ray_aabb_1 <= 1'h0; // @[Schedule_unit_1.scala 54:46]
    end else begin
      ray_aabb_1 <= io_RAY_AABB_1; // @[Schedule_unit_1.scala 67:40]
    end
    if (reset) begin // @[Schedule_unit_1.scala 55:46]
      ray_aabb_2 <= 1'h0; // @[Schedule_unit_1.scala 55:46]
    end else begin
      ray_aabb_2 <= io_RAY_AABB_2; // @[Schedule_unit_1.scala 68:40]
    end
    if (reset) begin // @[Schedule_unit_1.scala 70:42]
      v11_temp_2 <= 128'h0; // @[Schedule_unit_1.scala 70:42]
    end else begin
      v11_temp_2 <= v11_temp_1; // @[Schedule_unit_1.scala 83:57]
    end
    if (reset) begin // @[Schedule_unit_1.scala 71:42]
      v22_temp_2 <= 128'h0; // @[Schedule_unit_1.scala 71:42]
    end else begin
      v22_temp_2 <= v22_temp_1; // @[Schedule_unit_1.scala 84:57]
    end
    if (reset) begin // @[Schedule_unit_1.scala 72:43]
      ray_temp_2 <= 32'h0; // @[Schedule_unit_1.scala 72:43]
    end else begin
      ray_temp_2 <= ray_temp_1; // @[Schedule_unit_1.scala 85:58]
    end
    if (reset) begin // @[Schedule_unit_1.scala 73:43]
      Oz_temp_2 <= 32'h0; // @[Schedule_unit_1.scala 73:43]
    end else begin
      Oz_temp_2 <= Oz_temp_1; // @[Schedule_unit_1.scala 86:54]
    end
    if (reset) begin // @[Schedule_unit_1.scala 74:40]
      ray_o_temp_2 <= 96'h0; // @[Schedule_unit_1.scala 74:40]
    end else begin
      ray_o_temp_2 <= ray_o_temp_1; // @[Schedule_unit_1.scala 87:39]
    end
    if (reset) begin // @[Schedule_unit_1.scala 75:40]
      ray_d_temp_2 <= 96'h0; // @[Schedule_unit_1.scala 75:40]
    end else begin
      ray_d_temp_2 <= ray_d_temp_1; // @[Schedule_unit_1.scala 88:39]
    end
    if (reset) begin // @[Schedule_unit_1.scala 76:37]
      node_id_temp_2 <= 32'sh0; // @[Schedule_unit_1.scala 76:37]
    end else begin
      node_id_temp_2 <= node_id_temp_1; // @[Schedule_unit_1.scala 89:35]
    end
    if (reset) begin // @[Schedule_unit_1.scala 77:43]
      hitT_temp_2 <= 32'h0; // @[Schedule_unit_1.scala 77:43]
    end else begin
      hitT_temp_2 <= hitT_temp_1; // @[Schedule_unit_1.scala 90:57]
    end
    if (reset) begin // @[Schedule_unit_1.scala 78:61]
      inValid_2 <= 1'h0; // @[Schedule_unit_1.scala 78:61]
    end else begin
      inValid_2 <= inValid_1; // @[Schedule_unit_1.scala 91:66]
    end
    if (reset) begin // @[Schedule_unit_1.scala 79:45]
      break_2 <= 1'h0; // @[Schedule_unit_1.scala 79:45]
    end else begin
      break_2 <= break_1; // @[Schedule_unit_1.scala 92:39]
    end
    if (reset) begin // @[Schedule_unit_1.scala 80:43]
      ray_aabb_1_2 <= 1'h0; // @[Schedule_unit_1.scala 80:43]
    end else begin
      ray_aabb_1_2 <= ray_aabb_1; // @[Schedule_unit_1.scala 93:37]
    end
    if (reset) begin // @[Schedule_unit_1.scala 81:43]
      ray_aabb_2_2 <= 1'h0; // @[Schedule_unit_1.scala 81:43]
    end else begin
      ray_aabb_2_2 <= ray_aabb_2; // @[Schedule_unit_1.scala 94:37]
    end
    if (reset) begin // @[Schedule_unit_1.scala 96:42]
      v11_temp_3 <= 128'h0; // @[Schedule_unit_1.scala 96:42]
    end else begin
      v11_temp_3 <= v11_temp_2; // @[Schedule_unit_1.scala 109:57]
    end
    if (reset) begin // @[Schedule_unit_1.scala 97:42]
      v22_temp_3 <= 128'h0; // @[Schedule_unit_1.scala 97:42]
    end else begin
      v22_temp_3 <= v22_temp_2; // @[Schedule_unit_1.scala 110:57]
    end
    if (reset) begin // @[Schedule_unit_1.scala 98:43]
      ray_temp_3 <= 32'h0; // @[Schedule_unit_1.scala 98:43]
    end else begin
      ray_temp_3 <= ray_temp_2; // @[Schedule_unit_1.scala 111:58]
    end
    if (reset) begin // @[Schedule_unit_1.scala 99:43]
      Oz_temp_3 <= 32'h0; // @[Schedule_unit_1.scala 99:43]
    end else begin
      Oz_temp_3 <= Oz_temp_2; // @[Schedule_unit_1.scala 112:54]
    end
    if (reset) begin // @[Schedule_unit_1.scala 100:40]
      ray_o_temp_3 <= 96'h0; // @[Schedule_unit_1.scala 100:40]
    end else begin
      ray_o_temp_3 <= ray_o_temp_2; // @[Schedule_unit_1.scala 113:39]
    end
    if (reset) begin // @[Schedule_unit_1.scala 101:40]
      ray_d_temp_3 <= 96'h0; // @[Schedule_unit_1.scala 101:40]
    end else begin
      ray_d_temp_3 <= ray_d_temp_2; // @[Schedule_unit_1.scala 114:39]
    end
    if (reset) begin // @[Schedule_unit_1.scala 102:37]
      node_id_temp_3 <= 32'sh0; // @[Schedule_unit_1.scala 102:37]
    end else begin
      node_id_temp_3 <= node_id_temp_2; // @[Schedule_unit_1.scala 115:35]
    end
    if (reset) begin // @[Schedule_unit_1.scala 103:43]
      hitT_temp_3 <= 32'h0; // @[Schedule_unit_1.scala 103:43]
    end else begin
      hitT_temp_3 <= hitT_temp_2; // @[Schedule_unit_1.scala 116:49]
    end
    if (reset) begin // @[Schedule_unit_1.scala 104:61]
      inValid_3 <= 1'h0; // @[Schedule_unit_1.scala 104:61]
    end else begin
      inValid_3 <= inValid_2; // @[Schedule_unit_1.scala 117:66]
    end
    if (reset) begin // @[Schedule_unit_1.scala 105:45]
      break_3 <= 1'h0; // @[Schedule_unit_1.scala 105:45]
    end else begin
      break_3 <= break_2; // @[Schedule_unit_1.scala 118:39]
    end
    if (reset) begin // @[Schedule_unit_1.scala 106:43]
      ray_aabb_1_3 <= 1'h0; // @[Schedule_unit_1.scala 106:43]
    end else begin
      ray_aabb_1_3 <= ray_aabb_1_2; // @[Schedule_unit_1.scala 119:37]
    end
    if (reset) begin // @[Schedule_unit_1.scala 107:43]
      ray_aabb_2_3 <= 1'h0; // @[Schedule_unit_1.scala 107:43]
    end else begin
      ray_aabb_2_3 <= ray_aabb_2_2; // @[Schedule_unit_1.scala 120:37]
    end
    if (reset) begin // @[Schedule_unit_1.scala 121:38]
      v11_temp_4 <= 128'h0; // @[Schedule_unit_1.scala 121:38]
    end else begin
      v11_temp_4 <= v11_temp_3; // @[Schedule_unit_1.scala 134:57]
    end
    if (reset) begin // @[Schedule_unit_1.scala 122:42]
      v22_temp_4 <= 128'h0; // @[Schedule_unit_1.scala 122:42]
    end else begin
      v22_temp_4 <= v22_temp_3; // @[Schedule_unit_1.scala 135:57]
    end
    if (reset) begin // @[Schedule_unit_1.scala 123:43]
      ray_temp_4 <= 32'h0; // @[Schedule_unit_1.scala 123:43]
    end else begin
      ray_temp_4 <= ray_temp_3; // @[Schedule_unit_1.scala 136:58]
    end
    if (reset) begin // @[Schedule_unit_1.scala 124:43]
      Oz_temp_4 <= 32'h0; // @[Schedule_unit_1.scala 124:43]
    end else begin
      Oz_temp_4 <= Oz_temp_3; // @[Schedule_unit_1.scala 137:54]
    end
    if (reset) begin // @[Schedule_unit_1.scala 125:40]
      ray_o_temp_4 <= 96'h0; // @[Schedule_unit_1.scala 125:40]
    end else begin
      ray_o_temp_4 <= ray_o_temp_3; // @[Schedule_unit_1.scala 138:39]
    end
    if (reset) begin // @[Schedule_unit_1.scala 126:40]
      ray_d_temp_4 <= 96'h0; // @[Schedule_unit_1.scala 126:40]
    end else begin
      ray_d_temp_4 <= ray_d_temp_3; // @[Schedule_unit_1.scala 139:39]
    end
    if (reset) begin // @[Schedule_unit_1.scala 127:37]
      node_id_temp_4 <= 32'sh0; // @[Schedule_unit_1.scala 127:37]
    end else begin
      node_id_temp_4 <= node_id_temp_3; // @[Schedule_unit_1.scala 140:35]
    end
    if (reset) begin // @[Schedule_unit_1.scala 128:43]
      hitT_temp_4 <= 32'h0; // @[Schedule_unit_1.scala 128:43]
    end else begin
      hitT_temp_4 <= hitT_temp_3; // @[Schedule_unit_1.scala 141:49]
    end
    if (reset) begin // @[Schedule_unit_1.scala 129:61]
      inValid_4 <= 1'h0; // @[Schedule_unit_1.scala 129:61]
    end else begin
      inValid_4 <= inValid_3; // @[Schedule_unit_1.scala 142:66]
    end
    if (reset) begin // @[Schedule_unit_1.scala 130:45]
      break_4 <= 1'h0; // @[Schedule_unit_1.scala 130:45]
    end else begin
      break_4 <= break_3; // @[Schedule_unit_1.scala 143:39]
    end
    if (reset) begin // @[Schedule_unit_1.scala 131:43]
      ray_aabb_1_4 <= 1'h0; // @[Schedule_unit_1.scala 131:43]
    end else begin
      ray_aabb_1_4 <= ray_aabb_1_3; // @[Schedule_unit_1.scala 144:37]
    end
    if (reset) begin // @[Schedule_unit_1.scala 132:43]
      ray_aabb_2_4 <= 1'h0; // @[Schedule_unit_1.scala 132:43]
    end else begin
      ray_aabb_2_4 <= ray_aabb_2_3; // @[Schedule_unit_1.scala 145:37]
    end
    if (reset) begin // @[Schedule_unit_1.scala 171:46]
      count <= 64'h0; // @[Schedule_unit_1.scala 171:46]
    end else if (io_valid_in) begin // @[Schedule_unit_1.scala 190:22]
      count <= _T_19; // @[Schedule_unit_1.scala 191:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  v11_temp_1 = _RAND_0[127:0];
  _RAND_1 = {4{`RANDOM}};
  v22_temp_1 = _RAND_1[127:0];
  _RAND_2 = {1{`RANDOM}};
  ray_temp_1 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  Oz_temp_1 = _RAND_3[31:0];
  _RAND_4 = {3{`RANDOM}};
  ray_o_temp_1 = _RAND_4[95:0];
  _RAND_5 = {3{`RANDOM}};
  ray_d_temp_1 = _RAND_5[95:0];
  _RAND_6 = {1{`RANDOM}};
  node_id_temp_1 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  hitT_temp_1 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  inValid_1 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  break_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  ray_aabb_1 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ray_aabb_2 = _RAND_11[0:0];
  _RAND_12 = {4{`RANDOM}};
  v11_temp_2 = _RAND_12[127:0];
  _RAND_13 = {4{`RANDOM}};
  v22_temp_2 = _RAND_13[127:0];
  _RAND_14 = {1{`RANDOM}};
  ray_temp_2 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  Oz_temp_2 = _RAND_15[31:0];
  _RAND_16 = {3{`RANDOM}};
  ray_o_temp_2 = _RAND_16[95:0];
  _RAND_17 = {3{`RANDOM}};
  ray_d_temp_2 = _RAND_17[95:0];
  _RAND_18 = {1{`RANDOM}};
  node_id_temp_2 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  hitT_temp_2 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  inValid_2 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  break_2 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  ray_aabb_1_2 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  ray_aabb_2_2 = _RAND_23[0:0];
  _RAND_24 = {4{`RANDOM}};
  v11_temp_3 = _RAND_24[127:0];
  _RAND_25 = {4{`RANDOM}};
  v22_temp_3 = _RAND_25[127:0];
  _RAND_26 = {1{`RANDOM}};
  ray_temp_3 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  Oz_temp_3 = _RAND_27[31:0];
  _RAND_28 = {3{`RANDOM}};
  ray_o_temp_3 = _RAND_28[95:0];
  _RAND_29 = {3{`RANDOM}};
  ray_d_temp_3 = _RAND_29[95:0];
  _RAND_30 = {1{`RANDOM}};
  node_id_temp_3 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  hitT_temp_3 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  inValid_3 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  break_3 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  ray_aabb_1_3 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  ray_aabb_2_3 = _RAND_35[0:0];
  _RAND_36 = {4{`RANDOM}};
  v11_temp_4 = _RAND_36[127:0];
  _RAND_37 = {4{`RANDOM}};
  v22_temp_4 = _RAND_37[127:0];
  _RAND_38 = {1{`RANDOM}};
  ray_temp_4 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  Oz_temp_4 = _RAND_39[31:0];
  _RAND_40 = {3{`RANDOM}};
  ray_o_temp_4 = _RAND_40[95:0];
  _RAND_41 = {3{`RANDOM}};
  ray_d_temp_4 = _RAND_41[95:0];
  _RAND_42 = {1{`RANDOM}};
  node_id_temp_4 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  hitT_temp_4 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  inValid_4 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  break_4 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  ray_aabb_1_4 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  ray_aabb_2_4 = _RAND_47[0:0];
  _RAND_48 = {2{`RANDOM}};
  count = _RAND_48[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IST1(
  input         clock,
  input         reset,
  input         io_enable_IST1,
  input  [31:0] io_nodeid_leaf_1,
  input  [31:0] io_rayid_leaf_1,
  input  [31:0] io_hiT_in,
  input  [31:0] io_Oz,
  input  [31:0] io_invDz,
  input  [31:0] io_v11_in_x,
  input  [31:0] io_v11_in_y,
  input  [31:0] io_v11_in_z,
  input  [31:0] io_v11_in_w,
  input  [31:0] io_v22_in_x,
  input  [31:0] io_v22_in_y,
  input  [31:0] io_v22_in_z,
  input  [31:0] io_v22_in_w,
  input  [31:0] io_ray_o_in_x,
  input  [31:0] io_ray_o_in_y,
  input  [31:0] io_ray_o_in_z,
  input  [31:0] io_ray_d_in_x,
  input  [31:0] io_ray_d_in_y,
  input  [31:0] io_ray_d_in_z,
  input         io_break_in,
  input         io_RAY_AABB_1,
  input         io_RAY_AABB_2,
  output [31:0] io_nodeid_ist1_out,
  output [31:0] io_rayid_ist1_out,
  output [31:0] io_hiT_out,
  output [31:0] io_t,
  output        io_pop_1,
  output [31:0] io_v11_out_x,
  output [31:0] io_v11_out_y,
  output [31:0] io_v11_out_z,
  output [31:0] io_v11_out_w,
  output [31:0] io_v22_out_x,
  output [31:0] io_v22_out_y,
  output [31:0] io_v22_out_z,
  output [31:0] io_v22_out_w,
  output [31:0] io_ray_o_out_x,
  output [31:0] io_ray_o_out_y,
  output [31:0] io_ray_o_out_z,
  output [31:0] io_ray_d_out_x,
  output [31:0] io_ray_d_out_y,
  output [31:0] io_ray_d_out_z,
  output        io_enable_IST2,
  output        io_break_out,
  output        io_break_ist1,
  output        io_RAY_AABB_1_out,
  output        io_RAY_AABB_2_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [127:0] _RAND_5;
  reg [127:0] _RAND_6;
  reg [95:0] _RAND_7;
  reg [95:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [127:0] _RAND_16;
  reg [127:0] _RAND_17;
  reg [95:0] _RAND_18;
  reg [95:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [127:0] _RAND_29;
  reg [127:0] _RAND_30;
  reg [95:0] _RAND_31;
  reg [95:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
`endif // RANDOMIZE_REG_INIT
  wire  FMUL_6_clock; // @[IST1.scala 69:24]
  wire  FMUL_6_reset; // @[IST1.scala 69:24]
  wire [31:0] FMUL_6_io_a; // @[IST1.scala 69:24]
  wire [31:0] FMUL_6_io_b; // @[IST1.scala 69:24]
  wire [31:0] FMUL_6_io_out; // @[IST1.scala 69:24]
  wire [31:0] FCMP_21_io_a; // @[IST1.scala 131:25]
  wire [31:0] FCMP_21_io_b; // @[IST1.scala 131:25]
  wire  FCMP_21_io_actual_out; // @[IST1.scala 131:25]
  wire [31:0] FCMP_22_io_a; // @[IST1.scala 141:25]
  wire [31:0] FCMP_22_io_b; // @[IST1.scala 141:25]
  wire  FCMP_22_io_actual_out; // @[IST1.scala 141:25]
  reg  enable_1; // @[IST1.scala 45:52]
  reg [31:0] nodeid_ist1_temp_1; // @[IST1.scala 46:38]
  reg [31:0] rayid_ist1_temp_1; // @[IST1.scala 47:41]
  reg [31:0] hitT_temp_1; // @[IST1.scala 48:47]
  reg [31:0] t_1; // @[IST1.scala 49:59]
  reg [127:0] v11_1; // @[IST1.scala 50:56]
  reg [127:0] v22_1; // @[IST1.scala 51:56]
  reg [95:0] ray_o_in_1; // @[IST1.scala 52:50]
  reg [95:0] ray_d_in_1; // @[IST1.scala 53:50]
  reg  break_1; // @[IST1.scala 54:54]
  reg  ray_aabb_1; // @[IST1.scala 55:46]
  reg  ray_aabb_2; // @[IST1.scala 56:46]
  wire [127:0] _T = {io_v11_in_w,io_v11_in_z,io_v11_in_y,io_v11_in_x}; // @[Cat.scala 30:58]
  wire [127:0] _T_1 = {io_v22_in_w,io_v22_in_z,io_v22_in_y,io_v22_in_x}; // @[Cat.scala 30:58]
  wire [95:0] _T_2 = {io_ray_o_in_z,io_ray_o_in_y,io_ray_o_in_x}; // @[Cat.scala 30:58]
  wire [95:0] _T_3 = {io_ray_d_in_z,io_ray_d_in_y,io_ray_d_in_x}; // @[Cat.scala 30:58]
  reg  mul_enable_1; // @[IST1.scala 78:56]
  reg [31:0] mul_nodeid_ist1_temp_1; // @[IST1.scala 79:42]
  reg [31:0] mul_rayid_ist1_temp_1; // @[IST1.scala 80:45]
  reg [31:0] mul_hitT_temp_1; // @[IST1.scala 81:51]
  reg [127:0] mul_v11_1; // @[IST1.scala 83:60]
  reg [127:0] mul_v22_1; // @[IST1.scala 84:60]
  reg [95:0] mul_ray_o_in_1; // @[IST1.scala 85:54]
  reg [95:0] mul_ray_d_in_1; // @[IST1.scala 86:54]
  reg  mul_break_1; // @[IST1.scala 87:58]
  reg  mul_ray_aabb_1; // @[IST1.scala 88:50]
  reg  mul_ray_aabb_2; // @[IST1.scala 89:50]
  reg [31:0] nodeid_ist1_temp_2; // @[IST1.scala 104:38]
  reg [31:0] rayid_ist1_temp_2; // @[IST1.scala 105:41]
  reg [31:0] hitT_temp_2; // @[IST1.scala 106:47]
  reg [31:0] t_2; // @[IST1.scala 107:59]
  reg  t_min; // @[IST1.scala 108:54]
  reg  t_hitT; // @[IST1.scala 109:55]
  reg [127:0] v11_2; // @[IST1.scala 110:56]
  reg [127:0] v22_2; // @[IST1.scala 111:56]
  reg [95:0] ray_o_in_2; // @[IST1.scala 112:50]
  reg [95:0] ray_d_in_2; // @[IST1.scala 113:50]
  reg  enable_2; // @[IST1.scala 114:50]
  reg  break_2; // @[IST1.scala 115:52]
  reg  ray_aabb_1_2; // @[IST1.scala 116:43]
  reg  ray_aabb_2_2; // @[IST1.scala 117:43]
  wire  _T_4 = FCMP_21_io_actual_out > 1'h0; // @[IST1.scala 136:36]
  wire  _T_5 = FCMP_22_io_actual_out > 1'h0; // @[IST1.scala 146:36]
  wire  _T_20 = t_min & t_hitT; // @[IST1.scala 173:19]
  wire  _T_23 = t_min & t_hitT & enable_2; // @[IST1.scala 173:36]
  wire  _T_24 = ~break_2; // @[IST1.scala 173:64]
  wire  _T_29 = ~_T_20 & enable_2; // @[IST1.scala 178:41]
  wire  _T_31 = ~_T_20 & enable_2 & _T_24; // @[IST1.scala 178:59]
  wire  _T_37 = _T_23 & break_2; // @[IST1.scala 183:59]
  wire  _T_43 = _T_29 & break_2; // @[IST1.scala 188:59]
  wire  _GEN_6 = _T_23 & break_2 ? 1'h0 : _T_43; // @[IST1.scala 183:77 IST1.scala 187:31]
  wire  _GEN_7 = ~_T_20 & enable_2 & _T_24 ? 1'h0 : _T_37; // @[IST1.scala 178:77 IST1.scala 179:28]
  wire  _GEN_9 = ~_T_20 & enable_2 & _T_24 ? 1'h0 : _GEN_6; // @[IST1.scala 178:77 IST1.scala 182:31]
  MY_MUL FMUL_6 ( // @[IST1.scala 69:24]
    .clock(FMUL_6_clock),
    .reset(FMUL_6_reset),
    .io_a(FMUL_6_io_a),
    .io_b(FMUL_6_io_b),
    .io_out(FMUL_6_io_out)
  );
  ValExec_CompareRecF32_lt FCMP_21 ( // @[IST1.scala 131:25]
    .io_a(FCMP_21_io_a),
    .io_b(FCMP_21_io_b),
    .io_actual_out(FCMP_21_io_actual_out)
  );
  ValExec_CompareRecF32_lt FCMP_22 ( // @[IST1.scala 141:25]
    .io_a(FCMP_22_io_a),
    .io_b(FCMP_22_io_b),
    .io_actual_out(FCMP_22_io_actual_out)
  );
  assign io_nodeid_ist1_out = nodeid_ist1_temp_2; // @[IST1.scala 160:39]
  assign io_rayid_ist1_out = rayid_ist1_temp_2; // @[IST1.scala 161:42]
  assign io_hiT_out = hitT_temp_2; // @[IST1.scala 163:49]
  assign io_t = t_2; // @[IST1.scala 162:58]
  assign io_pop_1 = t_min & t_hitT & enable_2 & ~break_2 ? 1'h0 : _T_31; // @[IST1.scala 173:72 IST1.scala 175:35]
  assign io_v11_out_x = v11_2[31:0]; // @[IST1.scala 152:52]
  assign io_v11_out_y = v11_2[63:32]; // @[IST1.scala 153:52]
  assign io_v11_out_z = v11_2[95:64]; // @[IST1.scala 154:52]
  assign io_v11_out_w = v11_2[127:96]; // @[IST1.scala 155:51]
  assign io_v22_out_x = v22_2[31:0]; // @[IST1.scala 156:56]
  assign io_v22_out_y = v22_2[63:32]; // @[IST1.scala 157:56]
  assign io_v22_out_z = v22_2[95:64]; // @[IST1.scala 158:56]
  assign io_v22_out_w = v22_2[127:96]; // @[IST1.scala 159:54]
  assign io_ray_o_out_x = ray_o_in_2[31:0]; // @[IST1.scala 164:58]
  assign io_ray_o_out_y = ray_o_in_2[63:32]; // @[IST1.scala 165:58]
  assign io_ray_o_out_z = ray_o_in_2[95:64]; // @[IST1.scala 166:58]
  assign io_ray_d_out_x = ray_d_in_2[31:0]; // @[IST1.scala 167:58]
  assign io_ray_d_out_y = ray_d_in_2[63:32]; // @[IST1.scala 168:58]
  assign io_ray_d_out_z = ray_d_in_2[95:64]; // @[IST1.scala 169:58]
  assign io_enable_IST2 = t_min & t_hitT & enable_2 & ~break_2 | _GEN_7; // @[IST1.scala 173:72 IST1.scala 174:28]
  assign io_break_out = t_min & t_hitT & enable_2 & ~break_2 ? 1'h0 : _GEN_9; // @[IST1.scala 173:72 IST1.scala 177:31]
  assign io_break_ist1 = break_2; // @[IST1.scala 170:47]
  assign io_RAY_AABB_1_out = ray_aabb_1_2; // @[IST1.scala 171:36]
  assign io_RAY_AABB_2_out = ray_aabb_2_2; // @[IST1.scala 172:36]
  assign FMUL_6_clock = clock;
  assign FMUL_6_reset = reset;
  assign FMUL_6_io_a = io_Oz; // @[IST1.scala 70:21]
  assign FMUL_6_io_b = io_invDz; // @[IST1.scala 71:21]
  assign FCMP_21_io_a = 32'h0; // @[IST1.scala 132:22]
  assign FCMP_21_io_b = t_1; // @[IST1.scala 133:22]
  assign FCMP_22_io_a = t_1; // @[IST1.scala 142:22]
  assign FCMP_22_io_b = mul_hitT_temp_1; // @[IST1.scala 143:22]
  always @(posedge clock) begin
    if (reset) begin // @[IST1.scala 45:52]
      enable_1 <= 1'h0; // @[IST1.scala 45:52]
    end else begin
      enable_1 <= io_enable_IST1; // @[IST1.scala 65:43]
    end
    if (reset) begin // @[IST1.scala 46:38]
      nodeid_ist1_temp_1 <= 32'sh0; // @[IST1.scala 46:38]
    end else begin
      nodeid_ist1_temp_1 <= io_nodeid_leaf_1; // @[IST1.scala 58:29]
    end
    if (reset) begin // @[IST1.scala 47:41]
      rayid_ist1_temp_1 <= 32'h0; // @[IST1.scala 47:41]
    end else begin
      rayid_ist1_temp_1 <= io_rayid_leaf_1; // @[IST1.scala 59:32]
    end
    if (reset) begin // @[IST1.scala 48:47]
      hitT_temp_1 <= 32'h0; // @[IST1.scala 48:47]
    end else begin
      hitT_temp_1 <= io_hiT_in; // @[IST1.scala 60:38]
    end
    if (reset) begin // @[IST1.scala 49:59]
      t_1 <= 32'h0; // @[IST1.scala 49:59]
    end else begin
      t_1 <= FMUL_6_io_out; // @[IST1.scala 76:46]
    end
    if (reset) begin // @[IST1.scala 50:56]
      v11_1 <= 128'h0; // @[IST1.scala 50:56]
    end else begin
      v11_1 <= _T; // @[IST1.scala 61:46]
    end
    if (reset) begin // @[IST1.scala 51:56]
      v22_1 <= 128'h0; // @[IST1.scala 51:56]
    end else begin
      v22_1 <= _T_1; // @[IST1.scala 62:46]
    end
    if (reset) begin // @[IST1.scala 52:50]
      ray_o_in_1 <= 96'h0; // @[IST1.scala 52:50]
    end else begin
      ray_o_in_1 <= _T_2; // @[IST1.scala 63:40]
    end
    if (reset) begin // @[IST1.scala 53:50]
      ray_d_in_1 <= 96'h0; // @[IST1.scala 53:50]
    end else begin
      ray_d_in_1 <= _T_3; // @[IST1.scala 64:40]
    end
    if (reset) begin // @[IST1.scala 54:54]
      break_1 <= 1'h0; // @[IST1.scala 54:54]
    end else begin
      break_1 <= io_break_in; // @[IST1.scala 66:45]
    end
    if (reset) begin // @[IST1.scala 55:46]
      ray_aabb_1 <= 1'h0; // @[IST1.scala 55:46]
    end else begin
      ray_aabb_1 <= io_RAY_AABB_1; // @[IST1.scala 67:40]
    end
    if (reset) begin // @[IST1.scala 56:46]
      ray_aabb_2 <= 1'h0; // @[IST1.scala 56:46]
    end else begin
      ray_aabb_2 <= io_RAY_AABB_2; // @[IST1.scala 68:40]
    end
    if (reset) begin // @[IST1.scala 78:56]
      mul_enable_1 <= 1'h0; // @[IST1.scala 78:56]
    end else begin
      mul_enable_1 <= enable_1; // @[IST1.scala 98:47]
    end
    if (reset) begin // @[IST1.scala 79:42]
      mul_nodeid_ist1_temp_1 <= 32'sh0; // @[IST1.scala 79:42]
    end else begin
      mul_nodeid_ist1_temp_1 <= nodeid_ist1_temp_1; // @[IST1.scala 91:33]
    end
    if (reset) begin // @[IST1.scala 80:45]
      mul_rayid_ist1_temp_1 <= 32'h0; // @[IST1.scala 80:45]
    end else begin
      mul_rayid_ist1_temp_1 <= rayid_ist1_temp_1; // @[IST1.scala 92:36]
    end
    if (reset) begin // @[IST1.scala 81:51]
      mul_hitT_temp_1 <= 32'h0; // @[IST1.scala 81:51]
    end else begin
      mul_hitT_temp_1 <= hitT_temp_1; // @[IST1.scala 93:42]
    end
    if (reset) begin // @[IST1.scala 83:60]
      mul_v11_1 <= 128'h0; // @[IST1.scala 83:60]
    end else begin
      mul_v11_1 <= v11_1; // @[IST1.scala 94:50]
    end
    if (reset) begin // @[IST1.scala 84:60]
      mul_v22_1 <= 128'h0; // @[IST1.scala 84:60]
    end else begin
      mul_v22_1 <= v22_1; // @[IST1.scala 95:50]
    end
    if (reset) begin // @[IST1.scala 85:54]
      mul_ray_o_in_1 <= 96'h0; // @[IST1.scala 85:54]
    end else begin
      mul_ray_o_in_1 <= ray_o_in_1; // @[IST1.scala 96:44]
    end
    if (reset) begin // @[IST1.scala 86:54]
      mul_ray_d_in_1 <= 96'h0; // @[IST1.scala 86:54]
    end else begin
      mul_ray_d_in_1 <= ray_d_in_1; // @[IST1.scala 97:44]
    end
    if (reset) begin // @[IST1.scala 87:58]
      mul_break_1 <= 1'h0; // @[IST1.scala 87:58]
    end else begin
      mul_break_1 <= break_1; // @[IST1.scala 99:49]
    end
    if (reset) begin // @[IST1.scala 88:50]
      mul_ray_aabb_1 <= 1'h0; // @[IST1.scala 88:50]
    end else begin
      mul_ray_aabb_1 <= ray_aabb_1; // @[IST1.scala 100:45]
    end
    if (reset) begin // @[IST1.scala 89:50]
      mul_ray_aabb_2 <= 1'h0; // @[IST1.scala 89:50]
    end else begin
      mul_ray_aabb_2 <= ray_aabb_2; // @[IST1.scala 101:46]
    end
    if (reset) begin // @[IST1.scala 104:38]
      nodeid_ist1_temp_2 <= 32'sh0; // @[IST1.scala 104:38]
    end else begin
      nodeid_ist1_temp_2 <= mul_nodeid_ist1_temp_1; // @[IST1.scala 119:29]
    end
    if (reset) begin // @[IST1.scala 105:41]
      rayid_ist1_temp_2 <= 32'h0; // @[IST1.scala 105:41]
    end else begin
      rayid_ist1_temp_2 <= mul_rayid_ist1_temp_1; // @[IST1.scala 120:32]
    end
    if (reset) begin // @[IST1.scala 106:47]
      hitT_temp_2 <= 32'h0; // @[IST1.scala 106:47]
    end else begin
      hitT_temp_2 <= mul_hitT_temp_1; // @[IST1.scala 121:38]
    end
    if (reset) begin // @[IST1.scala 107:59]
      t_2 <= 32'h0; // @[IST1.scala 107:59]
    end else begin
      t_2 <= t_1; // @[IST1.scala 122:50]
    end
    if (reset) begin // @[IST1.scala 108:54]
      t_min <= 1'h0; // @[IST1.scala 108:54]
    end else begin
      t_min <= _T_4;
    end
    if (reset) begin // @[IST1.scala 109:55]
      t_hitT <= 1'h0; // @[IST1.scala 109:55]
    end else begin
      t_hitT <= _T_5;
    end
    if (reset) begin // @[IST1.scala 110:56]
      v11_2 <= 128'h0; // @[IST1.scala 110:56]
    end else begin
      v11_2 <= mul_v11_1; // @[IST1.scala 123:46]
    end
    if (reset) begin // @[IST1.scala 111:56]
      v22_2 <= 128'h0; // @[IST1.scala 111:56]
    end else begin
      v22_2 <= mul_v22_1; // @[IST1.scala 124:46]
    end
    if (reset) begin // @[IST1.scala 112:50]
      ray_o_in_2 <= 96'h0; // @[IST1.scala 112:50]
    end else begin
      ray_o_in_2 <= mul_ray_o_in_1; // @[IST1.scala 125:40]
    end
    if (reset) begin // @[IST1.scala 113:50]
      ray_d_in_2 <= 96'h0; // @[IST1.scala 113:50]
    end else begin
      ray_d_in_2 <= mul_ray_d_in_1; // @[IST1.scala 126:40]
    end
    if (reset) begin // @[IST1.scala 114:50]
      enable_2 <= 1'h0; // @[IST1.scala 114:50]
    end else begin
      enable_2 <= mul_enable_1; // @[IST1.scala 127:42]
    end
    if (reset) begin // @[IST1.scala 115:52]
      break_2 <= 1'h0; // @[IST1.scala 115:52]
    end else begin
      break_2 <= mul_break_1; // @[IST1.scala 128:44]
    end
    if (reset) begin // @[IST1.scala 116:43]
      ray_aabb_1_2 <= 1'h0; // @[IST1.scala 116:43]
    end else begin
      ray_aabb_1_2 <= mul_ray_aabb_1; // @[IST1.scala 129:37]
    end
    if (reset) begin // @[IST1.scala 117:43]
      ray_aabb_2_2 <= 1'h0; // @[IST1.scala 117:43]
    end else begin
      ray_aabb_2_2 <= mul_ray_aabb_2; // @[IST1.scala 130:37]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_1 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  nodeid_ist1_temp_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  rayid_ist1_temp_1 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  hitT_temp_1 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  t_1 = _RAND_4[31:0];
  _RAND_5 = {4{`RANDOM}};
  v11_1 = _RAND_5[127:0];
  _RAND_6 = {4{`RANDOM}};
  v22_1 = _RAND_6[127:0];
  _RAND_7 = {3{`RANDOM}};
  ray_o_in_1 = _RAND_7[95:0];
  _RAND_8 = {3{`RANDOM}};
  ray_d_in_1 = _RAND_8[95:0];
  _RAND_9 = {1{`RANDOM}};
  break_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  ray_aabb_1 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ray_aabb_2 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  mul_enable_1 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  mul_nodeid_ist1_temp_1 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  mul_rayid_ist1_temp_1 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  mul_hitT_temp_1 = _RAND_15[31:0];
  _RAND_16 = {4{`RANDOM}};
  mul_v11_1 = _RAND_16[127:0];
  _RAND_17 = {4{`RANDOM}};
  mul_v22_1 = _RAND_17[127:0];
  _RAND_18 = {3{`RANDOM}};
  mul_ray_o_in_1 = _RAND_18[95:0];
  _RAND_19 = {3{`RANDOM}};
  mul_ray_d_in_1 = _RAND_19[95:0];
  _RAND_20 = {1{`RANDOM}};
  mul_break_1 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  mul_ray_aabb_1 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  mul_ray_aabb_2 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  nodeid_ist1_temp_2 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  rayid_ist1_temp_2 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  hitT_temp_2 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  t_2 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  t_min = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  t_hitT = _RAND_28[0:0];
  _RAND_29 = {4{`RANDOM}};
  v11_2 = _RAND_29[127:0];
  _RAND_30 = {4{`RANDOM}};
  v22_2 = _RAND_30[127:0];
  _RAND_31 = {3{`RANDOM}};
  ray_o_in_2 = _RAND_31[95:0];
  _RAND_32 = {3{`RANDOM}};
  ray_d_in_2 = _RAND_32[95:0];
  _RAND_33 = {1{`RANDOM}};
  enable_2 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  break_2 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  ray_aabb_1_2 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  ray_aabb_2_2 = _RAND_36[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IST2(
  input         clock,
  input         reset,
  input         io_enable_IST2,
  input  [31:0] io_nodeid_leaf_2,
  input  [31:0] io_rayid_leaf_2,
  input  [31:0] io_hiT_in,
  input  [31:0] io_v11_in_x,
  input  [31:0] io_v11_in_y,
  input  [31:0] io_v11_in_z,
  input  [31:0] io_v11_in_w,
  input  [31:0] io_v22_in_x,
  input  [31:0] io_v22_in_y,
  input  [31:0] io_v22_in_z,
  input  [31:0] io_v22_in_w,
  input  [31:0] io_ray_o_in_x,
  input  [31:0] io_ray_o_in_y,
  input  [31:0] io_ray_o_in_z,
  input  [31:0] io_ray_d_in_x,
  input  [31:0] io_ray_d_in_y,
  input  [31:0] io_ray_d_in_z,
  input  [31:0] io_t,
  input         io_break_in,
  input         io_RAY_AABB_1,
  input         io_RAY_AABB_2,
  output [31:0] io_nodeid_ist2_out,
  output [31:0] io_rayid_ist2_out,
  output [31:0] io_hiT_out,
  output [31:0] io_u,
  output        io_pop_2,
  output [31:0] io_t_out,
  output [31:0] io_v22_out_x,
  output [31:0] io_v22_out_y,
  output [31:0] io_v22_out_z,
  output [31:0] io_v22_out_w,
  output [31:0] io_ray_o_out_x,
  output [31:0] io_ray_o_out_y,
  output [31:0] io_ray_o_out_z,
  output [31:0] io_ray_d_out_x,
  output [31:0] io_ray_d_out_y,
  output [31:0] io_ray_d_out_z,
  output        io_enable_IST3,
  output        io_break_ist2,
  output        io_break_out,
  output        io_RAY_AABB_1_out,
  output        io_RAY_AABB_2_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [127:0] _RAND_10;
  reg [95:0] _RAND_11;
  reg [95:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [127:0] _RAND_21;
  reg [95:0] _RAND_22;
  reg [95:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [127:0] _RAND_32;
  reg [95:0] _RAND_33;
  reg [95:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [127:0] _RAND_49;
  reg [95:0] _RAND_50;
  reg [95:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [127:0] _RAND_60;
  reg [95:0] _RAND_61;
  reg [95:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [127:0] _RAND_73;
  reg [95:0] _RAND_74;
  reg [95:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [127:0] _RAND_85;
  reg [95:0] _RAND_86;
  reg [95:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [127:0] _RAND_96;
  reg [95:0] _RAND_97;
  reg [95:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
`endif // RANDOMIZE_REG_INIT
  wire  FADD_MUL_14_clock; // @[IST2.scala 74:33]
  wire  FADD_MUL_14_reset; // @[IST2.scala 74:33]
  wire [31:0] FADD_MUL_14_io_a; // @[IST2.scala 74:33]
  wire [31:0] FADD_MUL_14_io_b; // @[IST2.scala 74:33]
  wire [31:0] FADD_MUL_14_io_c; // @[IST2.scala 74:33]
  wire [31:0] FADD_MUL_14_io_out; // @[IST2.scala 74:33]
  wire  FMUL_7_clock; // @[IST2.scala 84:24]
  wire  FMUL_7_reset; // @[IST2.scala 84:24]
  wire [31:0] FMUL_7_io_a; // @[IST2.scala 84:24]
  wire [31:0] FMUL_7_io_b; // @[IST2.scala 84:24]
  wire [31:0] FMUL_7_io_out; // @[IST2.scala 84:24]
  wire  FMUL_8_clock; // @[IST2.scala 93:24]
  wire  FMUL_8_reset; // @[IST2.scala 93:24]
  wire [31:0] FMUL_8_io_a; // @[IST2.scala 93:24]
  wire [31:0] FMUL_8_io_b; // @[IST2.scala 93:24]
  wire [31:0] FMUL_8_io_out; // @[IST2.scala 93:24]
  wire  FMUL_9_clock; // @[IST2.scala 102:24]
  wire  FMUL_9_reset; // @[IST2.scala 102:24]
  wire [31:0] FMUL_9_io_a; // @[IST2.scala 102:24]
  wire [31:0] FMUL_9_io_b; // @[IST2.scala 102:24]
  wire [31:0] FMUL_9_io_out; // @[IST2.scala 102:24]
  wire  FMUL_10_clock; // @[IST2.scala 111:25]
  wire  FMUL_10_reset; // @[IST2.scala 111:25]
  wire [31:0] FMUL_10_io_a; // @[IST2.scala 111:25]
  wire [31:0] FMUL_10_io_b; // @[IST2.scala 111:25]
  wire [31:0] FMUL_10_io_out; // @[IST2.scala 111:25]
  wire  FMUL_11_clock; // @[IST2.scala 120:25]
  wire  FMUL_11_reset; // @[IST2.scala 120:25]
  wire [31:0] FMUL_11_io_a; // @[IST2.scala 120:25]
  wire [31:0] FMUL_11_io_b; // @[IST2.scala 120:25]
  wire [31:0] FMUL_11_io_out; // @[IST2.scala 120:25]
  wire  FADD_5_clock; // @[IST2.scala 192:24]
  wire  FADD_5_reset; // @[IST2.scala 192:24]
  wire [31:0] FADD_5_io_a; // @[IST2.scala 192:24]
  wire [31:0] FADD_5_io_b; // @[IST2.scala 192:24]
  wire [31:0] FADD_5_io_out; // @[IST2.scala 192:24]
  wire  FADD_6_clock; // @[IST2.scala 201:24]
  wire  FADD_6_reset; // @[IST2.scala 201:24]
  wire [31:0] FADD_6_io_a; // @[IST2.scala 201:24]
  wire [31:0] FADD_6_io_b; // @[IST2.scala 201:24]
  wire [31:0] FADD_6_io_out; // @[IST2.scala 201:24]
  wire  FADD_7_clock; // @[IST2.scala 264:24]
  wire  FADD_7_reset; // @[IST2.scala 264:24]
  wire [31:0] FADD_7_io_a; // @[IST2.scala 264:24]
  wire [31:0] FADD_7_io_b; // @[IST2.scala 264:24]
  wire [31:0] FADD_7_io_out; // @[IST2.scala 264:24]
  wire  FADD_8_clock; // @[IST2.scala 273:24]
  wire  FADD_8_reset; // @[IST2.scala 273:24]
  wire [31:0] FADD_8_io_a; // @[IST2.scala 273:24]
  wire [31:0] FADD_8_io_b; // @[IST2.scala 273:24]
  wire [31:0] FADD_8_io_out; // @[IST2.scala 273:24]
  wire  FADD_MUL_15_clock; // @[IST2.scala 332:33]
  wire  FADD_MUL_15_reset; // @[IST2.scala 332:33]
  wire [31:0] FADD_MUL_15_io_a; // @[IST2.scala 332:33]
  wire [31:0] FADD_MUL_15_io_b; // @[IST2.scala 332:33]
  wire [31:0] FADD_MUL_15_io_c; // @[IST2.scala 332:33]
  wire [31:0] FADD_MUL_15_io_out; // @[IST2.scala 332:33]
  wire [31:0] FCMP_23_io_a; // @[IST2.scala 384:25]
  wire [31:0] FCMP_23_io_b; // @[IST2.scala 384:25]
  wire  FCMP_23_io_actual_out; // @[IST2.scala 384:25]
  reg [31:0] temp_0; // @[IST2.scala 44:33]
  reg [31:0] temp_1; // @[IST2.scala 45:33]
  reg [31:0] temp_2; // @[IST2.scala 46:33]
  reg [31:0] temp_3; // @[IST2.scala 47:33]
  reg [31:0] temp_4; // @[IST2.scala 48:33]
  reg [31:0] temp_5; // @[IST2.scala 49:33]
  reg [31:0] nodeid_ist2_temp_1_temp; // @[IST2.scala 51:42]
  reg [31:0] rayid_ist2_temp_1_temp; // @[IST2.scala 52:46]
  reg [31:0] t_temp_1_temp; // @[IST2.scala 53:56]
  reg [31:0] hitT_temp_1_temp; // @[IST2.scala 54:52]
  reg [127:0] v22_1_temp; // @[IST2.scala 55:60]
  reg [95:0] ray_o_in_1_temp; // @[IST2.scala 56:55]
  reg [95:0] ray_d_in_1_temp; // @[IST2.scala 57:55]
  reg  enable_1_temp; // @[IST2.scala 58:57]
  reg  break_1_temp; // @[IST2.scala 59:58]
  reg  ray_aabb_1_temp; // @[IST2.scala 60:51]
  reg  ray_aabb_2_temp; // @[IST2.scala 61:51]
  wire [127:0] _T = {io_v22_in_w,io_v22_in_z,io_v22_in_y,io_v22_in_x}; // @[Cat.scala 30:58]
  wire [95:0] _T_1 = {io_ray_o_in_z,io_ray_o_in_y,io_ray_o_in_x}; // @[Cat.scala 30:58]
  wire [95:0] _T_2 = {io_ray_d_in_z,io_ray_d_in_y,io_ray_d_in_x}; // @[Cat.scala 30:58]
  reg [31:0] nodeid_ist2_temp_1; // @[IST2.scala 129:37]
  reg [31:0] rayid_ist2_temp_1; // @[IST2.scala 130:41]
  reg [31:0] t_temp_1; // @[IST2.scala 131:51]
  reg [31:0] hitT_temp_1; // @[IST2.scala 132:47]
  reg [127:0] v22_1; // @[IST2.scala 133:55]
  reg [95:0] ray_o_in_1; // @[IST2.scala 134:50]
  reg [95:0] ray_d_in_1; // @[IST2.scala 135:50]
  reg  enable_1; // @[IST2.scala 136:52]
  reg  break_1; // @[IST2.scala 137:53]
  reg  ray_aabb_1; // @[IST2.scala 138:46]
  reg  ray_aabb_2; // @[IST2.scala 139:46]
  reg [31:0] nodeid_ist2_temp_2_temp; // @[IST2.scala 155:43]
  reg [31:0] rayid_ist2_temp_2_temp; // @[IST2.scala 156:46]
  reg [31:0] t_temp_2_temp; // @[IST2.scala 157:56]
  reg [31:0] hitT_temp_2_temp; // @[IST2.scala 158:52]
  reg [127:0] v22_2_temp; // @[IST2.scala 159:60]
  reg [95:0] ray_o_in_2_temp; // @[IST2.scala 160:55]
  reg [95:0] ray_d_in_2_temp; // @[IST2.scala 161:55]
  reg  enable_2_temp; // @[IST2.scala 162:55]
  reg  break_2_temp; // @[IST2.scala 163:58]
  reg  ray_aabb_1_2_temp; // @[IST2.scala 164:48]
  reg  ray_aabb_2_2_temp; // @[IST2.scala 165:48]
  reg [31:0] temp_6; // @[IST2.scala 179:50]
  reg [31:0] temp_7; // @[IST2.scala 180:50]
  reg [31:0] temp_0_2; // @[IST2.scala 181:47]
  reg [31:0] temp_0_3; // @[IST2.scala 182:47]
  reg [31:0] temp_5_2; // @[IST2.scala 184:46]
  reg [31:0] temp_5_3; // @[IST2.scala 185:46]
  reg [31:0] nodeid_ist2_temp_2; // @[IST2.scala 210:38]
  reg [31:0] rayid_ist2_temp_2; // @[IST2.scala 211:41]
  reg [31:0] t_temp_2; // @[IST2.scala 212:51]
  reg [31:0] hitT_temp_2; // @[IST2.scala 213:47]
  reg [127:0] v22_2; // @[IST2.scala 214:55]
  reg [95:0] ray_o_in_2; // @[IST2.scala 215:50]
  reg [95:0] ray_d_in_2; // @[IST2.scala 216:50]
  reg  enable_2; // @[IST2.scala 217:50]
  reg  break_2; // @[IST2.scala 218:53]
  reg  ray_aabb_1_2; // @[IST2.scala 219:43]
  reg  ray_aabb_2_2; // @[IST2.scala 220:43]
  reg [31:0] nodeid_ist2_temp_3_temp; // @[IST2.scala 236:43]
  reg [31:0] rayid_ist2_temp_3_temp; // @[IST2.scala 237:46]
  reg [31:0] t_temp_3_temp; // @[IST2.scala 238:56]
  reg [31:0] hitT_temp_3_temp; // @[IST2.scala 239:52]
  reg [127:0] v22_3_temp; // @[IST2.scala 240:60]
  reg [95:0] ray_o_in_3_temp; // @[IST2.scala 241:55]
  reg [95:0] ray_d_in_3_temp; // @[IST2.scala 242:55]
  reg  enable_3_temp; // @[IST2.scala 243:55]
  reg  break_3_temp; // @[IST2.scala 244:58]
  reg  ray_aabb_1_3_temp; // @[IST2.scala 245:48]
  reg  ray_aabb_2_3_temp; // @[IST2.scala 246:48]
  reg [31:0] Ox; // @[IST2.scala 261:58]
  reg [31:0] Dx; // @[IST2.scala 262:58]
  reg [31:0] nodeid_ist2_temp_3; // @[IST2.scala 282:38]
  reg [31:0] rayid_ist2_temp_3; // @[IST2.scala 283:41]
  reg [31:0] t_temp_3; // @[IST2.scala 284:51]
  reg [31:0] hitT_temp_3; // @[IST2.scala 285:47]
  reg [127:0] v22_3; // @[IST2.scala 286:55]
  reg [95:0] ray_o_in_3; // @[IST2.scala 287:50]
  reg [95:0] ray_d_in_3; // @[IST2.scala 288:50]
  reg  enable_3; // @[IST2.scala 289:50]
  reg  break_3; // @[IST2.scala 290:53]
  reg  ray_aabb_1_3; // @[IST2.scala 291:43]
  reg  ray_aabb_2_3; // @[IST2.scala 292:43]
  reg [31:0] nodeid_ist2_temp_4_temp; // @[IST2.scala 307:43]
  reg [31:0] rayid_ist2_temp_4_temp; // @[IST2.scala 308:46]
  reg [31:0] temp_u; // @[IST2.scala 309:53]
  reg [31:0] t_temp_4_temp; // @[IST2.scala 311:56]
  reg [31:0] hitT_temp_4_temp; // @[IST2.scala 312:52]
  reg [127:0] v22_4_temp; // @[IST2.scala 313:60]
  reg [95:0] ray_o_in_4_temp; // @[IST2.scala 314:55]
  reg [95:0] ray_d_in_4_temp; // @[IST2.scala 315:55]
  reg  enable_4_temp; // @[IST2.scala 316:55]
  reg  break_4_temp; // @[IST2.scala 317:58]
  reg  ray_aabb_1_4_temp; // @[IST2.scala 318:48]
  reg  ray_aabb_2_4_temp; // @[IST2.scala 319:48]
  reg [31:0] nodeid_ist2_temp_4; // @[IST2.scala 342:38]
  reg [31:0] rayid_ist2_temp_4; // @[IST2.scala 343:41]
  reg [31:0] t_temp_4; // @[IST2.scala 345:51]
  reg [31:0] hitT_temp_4; // @[IST2.scala 346:47]
  reg [127:0] v22_4; // @[IST2.scala 347:55]
  reg [95:0] ray_o_in_4; // @[IST2.scala 348:50]
  reg [95:0] ray_d_in_4; // @[IST2.scala 349:50]
  reg  enable_4; // @[IST2.scala 350:50]
  reg  break_4; // @[IST2.scala 351:53]
  reg  ray_aabb_1_4; // @[IST2.scala 352:43]
  reg  ray_aabb_2_4; // @[IST2.scala 353:43]
  wire  _T_15 = FCMP_23_io_actual_out > 1'h0 & enable_4; // @[IST2.scala 389:41]
  wire  _T_16 = ~break_4; // @[IST2.scala 389:69]
  wire  _T_20 = FCMP_23_io_actual_out < 1'h1 & enable_4; // @[IST2.scala 395:47]
  wire  _T_22 = FCMP_23_io_actual_out < 1'h1 & enable_4 & _T_16; // @[IST2.scala 395:65]
  wire  _T_27 = _T_15 & break_4; // @[IST2.scala 401:65]
  wire  _T_32 = _T_20 & break_4; // @[IST2.scala 407:65]
  wire  _GEN_6 = _T_15 & break_4 ? 1'h0 : _T_32; // @[IST2.scala 401:83 IST2.scala 406:34]
  wire  _GEN_9 = FCMP_23_io_actual_out < 1'h1 & enable_4 & _T_16 ? 1'h0 : _T_27; // @[IST2.scala 395:84 IST2.scala 399:32]
  wire  _GEN_10 = FCMP_23_io_actual_out < 1'h1 & enable_4 & _T_16 ? 1'h0 : _GEN_6; // @[IST2.scala 395:84 IST2.scala 400:34]
  MY_MULADD FADD_MUL_14 ( // @[IST2.scala 74:33]
    .clock(FADD_MUL_14_clock),
    .reset(FADD_MUL_14_reset),
    .io_a(FADD_MUL_14_io_a),
    .io_b(FADD_MUL_14_io_b),
    .io_c(FADD_MUL_14_io_c),
    .io_out(FADD_MUL_14_io_out)
  );
  MY_MUL FMUL_7 ( // @[IST2.scala 84:24]
    .clock(FMUL_7_clock),
    .reset(FMUL_7_reset),
    .io_a(FMUL_7_io_a),
    .io_b(FMUL_7_io_b),
    .io_out(FMUL_7_io_out)
  );
  MY_MUL FMUL_8 ( // @[IST2.scala 93:24]
    .clock(FMUL_8_clock),
    .reset(FMUL_8_reset),
    .io_a(FMUL_8_io_a),
    .io_b(FMUL_8_io_b),
    .io_out(FMUL_8_io_out)
  );
  MY_MUL FMUL_9 ( // @[IST2.scala 102:24]
    .clock(FMUL_9_clock),
    .reset(FMUL_9_reset),
    .io_a(FMUL_9_io_a),
    .io_b(FMUL_9_io_b),
    .io_out(FMUL_9_io_out)
  );
  MY_MUL FMUL_10 ( // @[IST2.scala 111:25]
    .clock(FMUL_10_clock),
    .reset(FMUL_10_reset),
    .io_a(FMUL_10_io_a),
    .io_b(FMUL_10_io_b),
    .io_out(FMUL_10_io_out)
  );
  MY_MUL FMUL_11 ( // @[IST2.scala 120:25]
    .clock(FMUL_11_clock),
    .reset(FMUL_11_reset),
    .io_a(FMUL_11_io_a),
    .io_b(FMUL_11_io_b),
    .io_out(FMUL_11_io_out)
  );
  MY_ADD FADD_5 ( // @[IST2.scala 192:24]
    .clock(FADD_5_clock),
    .reset(FADD_5_reset),
    .io_a(FADD_5_io_a),
    .io_b(FADD_5_io_b),
    .io_out(FADD_5_io_out)
  );
  MY_ADD FADD_6 ( // @[IST2.scala 201:24]
    .clock(FADD_6_clock),
    .reset(FADD_6_reset),
    .io_a(FADD_6_io_a),
    .io_b(FADD_6_io_b),
    .io_out(FADD_6_io_out)
  );
  MY_ADD FADD_7 ( // @[IST2.scala 264:24]
    .clock(FADD_7_clock),
    .reset(FADD_7_reset),
    .io_a(FADD_7_io_a),
    .io_b(FADD_7_io_b),
    .io_out(FADD_7_io_out)
  );
  MY_ADD FADD_8 ( // @[IST2.scala 273:24]
    .clock(FADD_8_clock),
    .reset(FADD_8_reset),
    .io_a(FADD_8_io_a),
    .io_b(FADD_8_io_b),
    .io_out(FADD_8_io_out)
  );
  MY_MULADD FADD_MUL_15 ( // @[IST2.scala 332:33]
    .clock(FADD_MUL_15_clock),
    .reset(FADD_MUL_15_reset),
    .io_a(FADD_MUL_15_io_a),
    .io_b(FADD_MUL_15_io_b),
    .io_c(FADD_MUL_15_io_c),
    .io_out(FADD_MUL_15_io_out)
  );
  ValExec_CompareRecF32_lt FCMP_23 ( // @[IST2.scala 384:25]
    .io_a(FCMP_23_io_a),
    .io_b(FCMP_23_io_b),
    .io_actual_out(FCMP_23_io_actual_out)
  );
  assign io_nodeid_ist2_out = nodeid_ist2_temp_4; // @[IST2.scala 367:37]
  assign io_rayid_ist2_out = rayid_ist2_temp_4; // @[IST2.scala 368:40]
  assign io_hiT_out = hitT_temp_4; // @[IST2.scala 370:47]
  assign io_u = temp_u; // @[IST2.scala 389:77 IST2.scala 390:45]
  assign io_pop_2 = FCMP_23_io_actual_out > 1'h0 & enable_4 & ~break_4 ? 1'h0 : _T_22; // @[IST2.scala 389:77 IST2.scala 392:38]
  assign io_t_out = t_temp_4; // @[IST2.scala 369:50]
  assign io_v22_out_x = v22_4[31:0]; // @[IST2.scala 371:53]
  assign io_v22_out_y = v22_4[63:32]; // @[IST2.scala 372:53]
  assign io_v22_out_z = v22_4[95:64]; // @[IST2.scala 373:53]
  assign io_v22_out_w = v22_4[127:96]; // @[IST2.scala 374:52]
  assign io_ray_o_out_x = ray_o_in_4[31:0]; // @[IST2.scala 375:54]
  assign io_ray_o_out_y = ray_o_in_4[63:32]; // @[IST2.scala 376:54]
  assign io_ray_o_out_z = ray_o_in_4[95:64]; // @[IST2.scala 377:54]
  assign io_ray_d_out_x = ray_d_in_4[31:0]; // @[IST2.scala 378:54]
  assign io_ray_d_out_y = ray_d_in_4[63:32]; // @[IST2.scala 379:54]
  assign io_ray_d_out_z = ray_d_in_4[95:64]; // @[IST2.scala 380:54]
  assign io_enable_IST3 = FCMP_23_io_actual_out > 1'h0 & enable_4 & ~break_4 | _GEN_9; // @[IST2.scala 389:77 IST2.scala 393:32]
  assign io_break_ist2 = break_4; // @[IST2.scala 381:43]
  assign io_break_out = FCMP_23_io_actual_out > 1'h0 & enable_4 & ~break_4 ? 1'h0 : _GEN_10; // @[IST2.scala 389:77 IST2.scala 394:34]
  assign io_RAY_AABB_1_out = ray_aabb_1_4; // @[IST2.scala 382:33]
  assign io_RAY_AABB_2_out = ray_aabb_2_4; // @[IST2.scala 383:33]
  assign FADD_MUL_14_clock = clock;
  assign FADD_MUL_14_reset = reset;
  assign FADD_MUL_14_io_a = io_ray_o_in_x; // @[IST2.scala 75:26]
  assign FADD_MUL_14_io_b = io_v11_in_x; // @[IST2.scala 76:26]
  assign FADD_MUL_14_io_c = io_v11_in_w; // @[IST2.scala 77:26]
  assign FMUL_7_clock = clock;
  assign FMUL_7_reset = reset;
  assign FMUL_7_io_a = io_ray_o_in_y; // @[IST2.scala 85:21]
  assign FMUL_7_io_b = io_v11_in_y; // @[IST2.scala 86:21]
  assign FMUL_8_clock = clock;
  assign FMUL_8_reset = reset;
  assign FMUL_8_io_a = io_ray_o_in_z; // @[IST2.scala 94:21]
  assign FMUL_8_io_b = io_v11_in_z; // @[IST2.scala 95:21]
  assign FMUL_9_clock = clock;
  assign FMUL_9_reset = reset;
  assign FMUL_9_io_a = io_ray_d_in_x; // @[IST2.scala 103:21]
  assign FMUL_9_io_b = io_v11_in_x; // @[IST2.scala 104:21]
  assign FMUL_10_clock = clock;
  assign FMUL_10_reset = reset;
  assign FMUL_10_io_a = io_ray_d_in_y; // @[IST2.scala 112:22]
  assign FMUL_10_io_b = io_v11_in_y; // @[IST2.scala 113:22]
  assign FMUL_11_clock = clock;
  assign FMUL_11_reset = reset;
  assign FMUL_11_io_a = io_ray_d_in_z; // @[IST2.scala 121:22]
  assign FMUL_11_io_b = io_v11_in_z; // @[IST2.scala 122:22]
  assign FADD_5_clock = clock;
  assign FADD_5_reset = reset;
  assign FADD_5_io_a = temp_1; // @[IST2.scala 193:21]
  assign FADD_5_io_b = temp_2; // @[IST2.scala 194:21]
  assign FADD_6_clock = clock;
  assign FADD_6_reset = reset;
  assign FADD_6_io_a = temp_3; // @[IST2.scala 202:21]
  assign FADD_6_io_b = temp_4; // @[IST2.scala 203:21]
  assign FADD_7_clock = clock;
  assign FADD_7_reset = reset;
  assign FADD_7_io_a = temp_0_3; // @[IST2.scala 265:21]
  assign FADD_7_io_b = temp_6; // @[IST2.scala 266:21]
  assign FADD_8_clock = clock;
  assign FADD_8_reset = reset;
  assign FADD_8_io_a = temp_5_3; // @[IST2.scala 274:21]
  assign FADD_8_io_b = temp_7; // @[IST2.scala 275:21]
  assign FADD_MUL_15_clock = clock;
  assign FADD_MUL_15_reset = reset;
  assign FADD_MUL_15_io_a = t_temp_3; // @[IST2.scala 333:26]
  assign FADD_MUL_15_io_b = Dx; // @[IST2.scala 334:26]
  assign FADD_MUL_15_io_c = Ox; // @[IST2.scala 335:26]
  assign FCMP_23_io_a = 32'h0; // @[IST2.scala 385:22]
  assign FCMP_23_io_b = temp_u; // @[IST2.scala 386:22]
  always @(posedge clock) begin
    if (reset) begin // @[IST2.scala 44:33]
      temp_0 <= 32'h0; // @[IST2.scala 44:33]
    end else begin
      temp_0 <= FADD_MUL_14_io_out; // @[IST2.scala 82:42]
    end
    if (reset) begin // @[IST2.scala 45:33]
      temp_1 <= 32'h0; // @[IST2.scala 45:33]
    end else begin
      temp_1 <= FMUL_7_io_out; // @[IST2.scala 91:42]
    end
    if (reset) begin // @[IST2.scala 46:33]
      temp_2 <= 32'h0; // @[IST2.scala 46:33]
    end else begin
      temp_2 <= FMUL_8_io_out; // @[IST2.scala 100:42]
    end
    if (reset) begin // @[IST2.scala 47:33]
      temp_3 <= 32'h0; // @[IST2.scala 47:33]
    end else begin
      temp_3 <= FMUL_9_io_out; // @[IST2.scala 109:42]
    end
    if (reset) begin // @[IST2.scala 48:33]
      temp_4 <= 32'h0; // @[IST2.scala 48:33]
    end else begin
      temp_4 <= FMUL_10_io_out; // @[IST2.scala 118:42]
    end
    if (reset) begin // @[IST2.scala 49:33]
      temp_5 <= 32'h0; // @[IST2.scala 49:33]
    end else begin
      temp_5 <= FMUL_11_io_out; // @[IST2.scala 127:42]
    end
    if (reset) begin // @[IST2.scala 51:42]
      nodeid_ist2_temp_1_temp <= 32'sh0; // @[IST2.scala 51:42]
    end else begin
      nodeid_ist2_temp_1_temp <= io_nodeid_leaf_2; // @[IST2.scala 63:34]
    end
    if (reset) begin // @[IST2.scala 52:46]
      rayid_ist2_temp_1_temp <= 32'h0; // @[IST2.scala 52:46]
    end else begin
      rayid_ist2_temp_1_temp <= io_rayid_leaf_2; // @[IST2.scala 64:37]
    end
    if (reset) begin // @[IST2.scala 53:56]
      t_temp_1_temp <= 32'h0; // @[IST2.scala 53:56]
    end else begin
      t_temp_1_temp <= io_t; // @[IST2.scala 65:47]
    end
    if (reset) begin // @[IST2.scala 54:52]
      hitT_temp_1_temp <= 32'h0; // @[IST2.scala 54:52]
    end else begin
      hitT_temp_1_temp <= io_hiT_in; // @[IST2.scala 66:43]
    end
    if (reset) begin // @[IST2.scala 55:60]
      v22_1_temp <= 128'h0; // @[IST2.scala 55:60]
    end else begin
      v22_1_temp <= _T; // @[IST2.scala 67:51]
    end
    if (reset) begin // @[IST2.scala 56:55]
      ray_o_in_1_temp <= 96'h0; // @[IST2.scala 56:55]
    end else begin
      ray_o_in_1_temp <= _T_1; // @[IST2.scala 68:45]
    end
    if (reset) begin // @[IST2.scala 57:55]
      ray_d_in_1_temp <= 96'h0; // @[IST2.scala 57:55]
    end else begin
      ray_d_in_1_temp <= _T_2; // @[IST2.scala 69:45]
    end
    if (reset) begin // @[IST2.scala 58:57]
      enable_1_temp <= 1'h0; // @[IST2.scala 58:57]
    end else begin
      enable_1_temp <= io_enable_IST2; // @[IST2.scala 70:48]
    end
    if (reset) begin // @[IST2.scala 59:58]
      break_1_temp <= 1'h0; // @[IST2.scala 59:58]
    end else begin
      break_1_temp <= io_break_in; // @[IST2.scala 71:50]
    end
    if (reset) begin // @[IST2.scala 60:51]
      ray_aabb_1_temp <= 1'h0; // @[IST2.scala 60:51]
    end else begin
      ray_aabb_1_temp <= io_RAY_AABB_1; // @[IST2.scala 72:45]
    end
    if (reset) begin // @[IST2.scala 61:51]
      ray_aabb_2_temp <= 1'h0; // @[IST2.scala 61:51]
    end else begin
      ray_aabb_2_temp <= io_RAY_AABB_2; // @[IST2.scala 73:45]
    end
    if (reset) begin // @[IST2.scala 129:37]
      nodeid_ist2_temp_1 <= 32'sh0; // @[IST2.scala 129:37]
    end else begin
      nodeid_ist2_temp_1 <= nodeid_ist2_temp_1_temp; // @[IST2.scala 141:29]
    end
    if (reset) begin // @[IST2.scala 130:41]
      rayid_ist2_temp_1 <= 32'h0; // @[IST2.scala 130:41]
    end else begin
      rayid_ist2_temp_1 <= rayid_ist2_temp_1_temp; // @[IST2.scala 142:32]
    end
    if (reset) begin // @[IST2.scala 131:51]
      t_temp_1 <= 32'h0; // @[IST2.scala 131:51]
    end else begin
      t_temp_1 <= t_temp_1_temp; // @[IST2.scala 143:42]
    end
    if (reset) begin // @[IST2.scala 132:47]
      hitT_temp_1 <= 32'h0; // @[IST2.scala 132:47]
    end else begin
      hitT_temp_1 <= hitT_temp_1_temp; // @[IST2.scala 144:38]
    end
    if (reset) begin // @[IST2.scala 133:55]
      v22_1 <= 128'h0; // @[IST2.scala 133:55]
    end else begin
      v22_1 <= v22_1_temp; // @[IST2.scala 145:46]
    end
    if (reset) begin // @[IST2.scala 134:50]
      ray_o_in_1 <= 96'h0; // @[IST2.scala 134:50]
    end else begin
      ray_o_in_1 <= ray_o_in_1_temp; // @[IST2.scala 146:40]
    end
    if (reset) begin // @[IST2.scala 135:50]
      ray_d_in_1 <= 96'h0; // @[IST2.scala 135:50]
    end else begin
      ray_d_in_1 <= ray_d_in_1_temp; // @[IST2.scala 147:40]
    end
    if (reset) begin // @[IST2.scala 136:52]
      enable_1 <= 1'h0; // @[IST2.scala 136:52]
    end else begin
      enable_1 <= enable_1_temp; // @[IST2.scala 148:43]
    end
    if (reset) begin // @[IST2.scala 137:53]
      break_1 <= 1'h0; // @[IST2.scala 137:53]
    end else begin
      break_1 <= break_1_temp; // @[IST2.scala 149:45]
    end
    if (reset) begin // @[IST2.scala 138:46]
      ray_aabb_1 <= 1'h0; // @[IST2.scala 138:46]
    end else begin
      ray_aabb_1 <= ray_aabb_1_temp; // @[IST2.scala 150:40]
    end
    if (reset) begin // @[IST2.scala 139:46]
      ray_aabb_2 <= 1'h0; // @[IST2.scala 139:46]
    end else begin
      ray_aabb_2 <= ray_aabb_2_temp; // @[IST2.scala 151:40]
    end
    if (reset) begin // @[IST2.scala 155:43]
      nodeid_ist2_temp_2_temp <= 32'sh0; // @[IST2.scala 155:43]
    end else begin
      nodeid_ist2_temp_2_temp <= nodeid_ist2_temp_1; // @[IST2.scala 167:34]
    end
    if (reset) begin // @[IST2.scala 156:46]
      rayid_ist2_temp_2_temp <= 32'h0; // @[IST2.scala 156:46]
    end else begin
      rayid_ist2_temp_2_temp <= rayid_ist2_temp_1; // @[IST2.scala 168:37]
    end
    if (reset) begin // @[IST2.scala 157:56]
      t_temp_2_temp <= 32'h0; // @[IST2.scala 157:56]
    end else begin
      t_temp_2_temp <= t_temp_1; // @[IST2.scala 169:47]
    end
    if (reset) begin // @[IST2.scala 158:52]
      hitT_temp_2_temp <= 32'h0; // @[IST2.scala 158:52]
    end else begin
      hitT_temp_2_temp <= hitT_temp_1; // @[IST2.scala 170:43]
    end
    if (reset) begin // @[IST2.scala 159:60]
      v22_2_temp <= 128'h0; // @[IST2.scala 159:60]
    end else begin
      v22_2_temp <= v22_1; // @[IST2.scala 171:51]
    end
    if (reset) begin // @[IST2.scala 160:55]
      ray_o_in_2_temp <= 96'h0; // @[IST2.scala 160:55]
    end else begin
      ray_o_in_2_temp <= ray_o_in_1; // @[IST2.scala 172:45]
    end
    if (reset) begin // @[IST2.scala 161:55]
      ray_d_in_2_temp <= 96'h0; // @[IST2.scala 161:55]
    end else begin
      ray_d_in_2_temp <= ray_d_in_1; // @[IST2.scala 173:45]
    end
    if (reset) begin // @[IST2.scala 162:55]
      enable_2_temp <= 1'h0; // @[IST2.scala 162:55]
    end else begin
      enable_2_temp <= enable_1; // @[IST2.scala 174:47]
    end
    if (reset) begin // @[IST2.scala 163:58]
      break_2_temp <= 1'h0; // @[IST2.scala 163:58]
    end else begin
      break_2_temp <= break_1; // @[IST2.scala 175:50]
    end
    if (reset) begin // @[IST2.scala 164:48]
      ray_aabb_1_2_temp <= 1'h0; // @[IST2.scala 164:48]
    end else begin
      ray_aabb_1_2_temp <= ray_aabb_1; // @[IST2.scala 176:41]
    end
    if (reset) begin // @[IST2.scala 165:48]
      ray_aabb_2_2_temp <= 1'h0; // @[IST2.scala 165:48]
    end else begin
      ray_aabb_2_2_temp <= ray_aabb_2; // @[IST2.scala 177:41]
    end
    if (reset) begin // @[IST2.scala 179:50]
      temp_6 <= 32'h0; // @[IST2.scala 179:50]
    end else begin
      temp_6 <= FADD_5_io_out; // @[IST2.scala 199:26]
    end
    if (reset) begin // @[IST2.scala 180:50]
      temp_7 <= 32'h0; // @[IST2.scala 180:50]
    end else begin
      temp_7 <= FADD_6_io_out; // @[IST2.scala 208:26]
    end
    if (reset) begin // @[IST2.scala 181:47]
      temp_0_2 <= 32'h0; // @[IST2.scala 181:47]
    end else begin
      temp_0_2 <= temp_0; // @[IST2.scala 186:41]
    end
    if (reset) begin // @[IST2.scala 182:47]
      temp_0_3 <= 32'h0; // @[IST2.scala 182:47]
    end else begin
      temp_0_3 <= temp_0_2; // @[IST2.scala 187:41]
    end
    if (reset) begin // @[IST2.scala 184:46]
      temp_5_2 <= 32'h0; // @[IST2.scala 184:46]
    end else begin
      temp_5_2 <= temp_5; // @[IST2.scala 188:41]
    end
    if (reset) begin // @[IST2.scala 185:46]
      temp_5_3 <= 32'h0; // @[IST2.scala 185:46]
    end else begin
      temp_5_3 <= temp_5_2; // @[IST2.scala 189:41]
    end
    if (reset) begin // @[IST2.scala 210:38]
      nodeid_ist2_temp_2 <= 32'sh0; // @[IST2.scala 210:38]
    end else begin
      nodeid_ist2_temp_2 <= nodeid_ist2_temp_2_temp; // @[IST2.scala 222:29]
    end
    if (reset) begin // @[IST2.scala 211:41]
      rayid_ist2_temp_2 <= 32'h0; // @[IST2.scala 211:41]
    end else begin
      rayid_ist2_temp_2 <= rayid_ist2_temp_2_temp; // @[IST2.scala 223:32]
    end
    if (reset) begin // @[IST2.scala 212:51]
      t_temp_2 <= 32'h0; // @[IST2.scala 212:51]
    end else begin
      t_temp_2 <= t_temp_2_temp; // @[IST2.scala 224:42]
    end
    if (reset) begin // @[IST2.scala 213:47]
      hitT_temp_2 <= 32'h0; // @[IST2.scala 213:47]
    end else begin
      hitT_temp_2 <= hitT_temp_2_temp; // @[IST2.scala 225:38]
    end
    if (reset) begin // @[IST2.scala 214:55]
      v22_2 <= 128'h0; // @[IST2.scala 214:55]
    end else begin
      v22_2 <= v22_2_temp; // @[IST2.scala 226:46]
    end
    if (reset) begin // @[IST2.scala 215:50]
      ray_o_in_2 <= 96'h0; // @[IST2.scala 215:50]
    end else begin
      ray_o_in_2 <= ray_o_in_2_temp; // @[IST2.scala 227:40]
    end
    if (reset) begin // @[IST2.scala 216:50]
      ray_d_in_2 <= 96'h0; // @[IST2.scala 216:50]
    end else begin
      ray_d_in_2 <= ray_d_in_2_temp; // @[IST2.scala 228:40]
    end
    if (reset) begin // @[IST2.scala 217:50]
      enable_2 <= 1'h0; // @[IST2.scala 217:50]
    end else begin
      enable_2 <= enable_2_temp; // @[IST2.scala 229:42]
    end
    if (reset) begin // @[IST2.scala 218:53]
      break_2 <= 1'h0; // @[IST2.scala 218:53]
    end else begin
      break_2 <= break_2_temp; // @[IST2.scala 230:45]
    end
    if (reset) begin // @[IST2.scala 219:43]
      ray_aabb_1_2 <= 1'h0; // @[IST2.scala 219:43]
    end else begin
      ray_aabb_1_2 <= ray_aabb_1_2_temp; // @[IST2.scala 231:37]
    end
    if (reset) begin // @[IST2.scala 220:43]
      ray_aabb_2_2 <= 1'h0; // @[IST2.scala 220:43]
    end else begin
      ray_aabb_2_2 <= ray_aabb_2_2_temp; // @[IST2.scala 232:37]
    end
    if (reset) begin // @[IST2.scala 236:43]
      nodeid_ist2_temp_3_temp <= 32'sh0; // @[IST2.scala 236:43]
    end else begin
      nodeid_ist2_temp_3_temp <= nodeid_ist2_temp_2; // @[IST2.scala 248:37]
    end
    if (reset) begin // @[IST2.scala 237:46]
      rayid_ist2_temp_3_temp <= 32'h0; // @[IST2.scala 237:46]
    end else begin
      rayid_ist2_temp_3_temp <= rayid_ist2_temp_2; // @[IST2.scala 249:40]
    end
    if (reset) begin // @[IST2.scala 238:56]
      t_temp_3_temp <= 32'h0; // @[IST2.scala 238:56]
    end else begin
      t_temp_3_temp <= t_temp_2; // @[IST2.scala 250:50]
    end
    if (reset) begin // @[IST2.scala 239:52]
      hitT_temp_3_temp <= 32'h0; // @[IST2.scala 239:52]
    end else begin
      hitT_temp_3_temp <= hitT_temp_2; // @[IST2.scala 251:46]
    end
    if (reset) begin // @[IST2.scala 240:60]
      v22_3_temp <= 128'h0; // @[IST2.scala 240:60]
    end else begin
      v22_3_temp <= v22_2; // @[IST2.scala 252:54]
    end
    if (reset) begin // @[IST2.scala 241:55]
      ray_o_in_3_temp <= 96'h0; // @[IST2.scala 241:55]
    end else begin
      ray_o_in_3_temp <= ray_o_in_2; // @[IST2.scala 253:45]
    end
    if (reset) begin // @[IST2.scala 242:55]
      ray_d_in_3_temp <= 96'h0; // @[IST2.scala 242:55]
    end else begin
      ray_d_in_3_temp <= ray_d_in_2; // @[IST2.scala 254:45]
    end
    if (reset) begin // @[IST2.scala 243:55]
      enable_3_temp <= 1'h0; // @[IST2.scala 243:55]
    end else begin
      enable_3_temp <= enable_2; // @[IST2.scala 255:47]
    end
    if (reset) begin // @[IST2.scala 244:58]
      break_3_temp <= 1'h0; // @[IST2.scala 244:58]
    end else begin
      break_3_temp <= break_2; // @[IST2.scala 256:49]
    end
    if (reset) begin // @[IST2.scala 245:48]
      ray_aabb_1_3_temp <= 1'h0; // @[IST2.scala 245:48]
    end else begin
      ray_aabb_1_3_temp <= ray_aabb_1_2; // @[IST2.scala 257:41]
    end
    if (reset) begin // @[IST2.scala 246:48]
      ray_aabb_2_3_temp <= 1'h0; // @[IST2.scala 246:48]
    end else begin
      ray_aabb_2_3_temp <= ray_aabb_2_2; // @[IST2.scala 258:41]
    end
    if (reset) begin // @[IST2.scala 261:58]
      Ox <= 32'h0; // @[IST2.scala 261:58]
    end else begin
      Ox <= FADD_7_io_out; // @[IST2.scala 271:26]
    end
    if (reset) begin // @[IST2.scala 262:58]
      Dx <= 32'h0; // @[IST2.scala 262:58]
    end else begin
      Dx <= FADD_8_io_out; // @[IST2.scala 280:26]
    end
    if (reset) begin // @[IST2.scala 282:38]
      nodeid_ist2_temp_3 <= 32'sh0; // @[IST2.scala 282:38]
    end else begin
      nodeid_ist2_temp_3 <= nodeid_ist2_temp_3_temp; // @[IST2.scala 294:32]
    end
    if (reset) begin // @[IST2.scala 283:41]
      rayid_ist2_temp_3 <= 32'h0; // @[IST2.scala 283:41]
    end else begin
      rayid_ist2_temp_3 <= rayid_ist2_temp_3_temp; // @[IST2.scala 295:35]
    end
    if (reset) begin // @[IST2.scala 284:51]
      t_temp_3 <= 32'h0; // @[IST2.scala 284:51]
    end else begin
      t_temp_3 <= t_temp_3_temp; // @[IST2.scala 296:45]
    end
    if (reset) begin // @[IST2.scala 285:47]
      hitT_temp_3 <= 32'h0; // @[IST2.scala 285:47]
    end else begin
      hitT_temp_3 <= hitT_temp_3_temp; // @[IST2.scala 297:41]
    end
    if (reset) begin // @[IST2.scala 286:55]
      v22_3 <= 128'h0; // @[IST2.scala 286:55]
    end else begin
      v22_3 <= v22_3_temp; // @[IST2.scala 298:49]
    end
    if (reset) begin // @[IST2.scala 287:50]
      ray_o_in_3 <= 96'h0; // @[IST2.scala 287:50]
    end else begin
      ray_o_in_3 <= ray_o_in_3_temp; // @[IST2.scala 299:40]
    end
    if (reset) begin // @[IST2.scala 288:50]
      ray_d_in_3 <= 96'h0; // @[IST2.scala 288:50]
    end else begin
      ray_d_in_3 <= ray_d_in_3_temp; // @[IST2.scala 300:40]
    end
    if (reset) begin // @[IST2.scala 289:50]
      enable_3 <= 1'h0; // @[IST2.scala 289:50]
    end else begin
      enable_3 <= enable_3_temp; // @[IST2.scala 301:42]
    end
    if (reset) begin // @[IST2.scala 290:53]
      break_3 <= 1'h0; // @[IST2.scala 290:53]
    end else begin
      break_3 <= break_3_temp; // @[IST2.scala 302:44]
    end
    if (reset) begin // @[IST2.scala 291:43]
      ray_aabb_1_3 <= 1'h0; // @[IST2.scala 291:43]
    end else begin
      ray_aabb_1_3 <= ray_aabb_1_3_temp; // @[IST2.scala 303:37]
    end
    if (reset) begin // @[IST2.scala 292:43]
      ray_aabb_2_3 <= 1'h0; // @[IST2.scala 292:43]
    end else begin
      ray_aabb_2_3 <= ray_aabb_2_3_temp; // @[IST2.scala 304:37]
    end
    if (reset) begin // @[IST2.scala 307:43]
      nodeid_ist2_temp_4_temp <= 32'sh0; // @[IST2.scala 307:43]
    end else begin
      nodeid_ist2_temp_4_temp <= nodeid_ist2_temp_3; // @[IST2.scala 321:37]
    end
    if (reset) begin // @[IST2.scala 308:46]
      rayid_ist2_temp_4_temp <= 32'h0; // @[IST2.scala 308:46]
    end else begin
      rayid_ist2_temp_4_temp <= rayid_ist2_temp_3; // @[IST2.scala 322:40]
    end
    if (reset) begin // @[IST2.scala 309:53]
      temp_u <= 32'h0; // @[IST2.scala 309:53]
    end else begin
      temp_u <= FADD_MUL_15_io_out; // @[IST2.scala 340:42]
    end
    if (reset) begin // @[IST2.scala 311:56]
      t_temp_4_temp <= 32'h0; // @[IST2.scala 311:56]
    end else begin
      t_temp_4_temp <= t_temp_3; // @[IST2.scala 323:50]
    end
    if (reset) begin // @[IST2.scala 312:52]
      hitT_temp_4_temp <= 32'h0; // @[IST2.scala 312:52]
    end else begin
      hitT_temp_4_temp <= hitT_temp_3; // @[IST2.scala 324:46]
    end
    if (reset) begin // @[IST2.scala 313:60]
      v22_4_temp <= 128'h0; // @[IST2.scala 313:60]
    end else begin
      v22_4_temp <= v22_3; // @[IST2.scala 325:54]
    end
    if (reset) begin // @[IST2.scala 314:55]
      ray_o_in_4_temp <= 96'h0; // @[IST2.scala 314:55]
    end else begin
      ray_o_in_4_temp <= ray_o_in_3; // @[IST2.scala 327:45]
    end
    if (reset) begin // @[IST2.scala 315:55]
      ray_d_in_4_temp <= 96'h0; // @[IST2.scala 315:55]
    end else begin
      ray_d_in_4_temp <= ray_d_in_3; // @[IST2.scala 326:45]
    end
    if (reset) begin // @[IST2.scala 316:55]
      enable_4_temp <= 1'h0; // @[IST2.scala 316:55]
    end else begin
      enable_4_temp <= enable_3; // @[IST2.scala 328:47]
    end
    if (reset) begin // @[IST2.scala 317:58]
      break_4_temp <= 1'h0; // @[IST2.scala 317:58]
    end else begin
      break_4_temp <= break_3; // @[IST2.scala 329:48]
    end
    if (reset) begin // @[IST2.scala 318:48]
      ray_aabb_1_4_temp <= 1'h0; // @[IST2.scala 318:48]
    end else begin
      ray_aabb_1_4_temp <= ray_aabb_1_3; // @[IST2.scala 330:42]
    end
    if (reset) begin // @[IST2.scala 319:48]
      ray_aabb_2_4_temp <= 1'h0; // @[IST2.scala 319:48]
    end else begin
      ray_aabb_2_4_temp <= ray_aabb_2_3; // @[IST2.scala 331:42]
    end
    if (reset) begin // @[IST2.scala 342:38]
      nodeid_ist2_temp_4 <= 32'sh0; // @[IST2.scala 342:38]
    end else begin
      nodeid_ist2_temp_4 <= nodeid_ist2_temp_4_temp; // @[IST2.scala 355:32]
    end
    if (reset) begin // @[IST2.scala 343:41]
      rayid_ist2_temp_4 <= 32'h0; // @[IST2.scala 343:41]
    end else begin
      rayid_ist2_temp_4 <= rayid_ist2_temp_4_temp; // @[IST2.scala 356:35]
    end
    if (reset) begin // @[IST2.scala 345:51]
      t_temp_4 <= 32'h0; // @[IST2.scala 345:51]
    end else begin
      t_temp_4 <= t_temp_4_temp; // @[IST2.scala 357:45]
    end
    if (reset) begin // @[IST2.scala 346:47]
      hitT_temp_4 <= 32'h0; // @[IST2.scala 346:47]
    end else begin
      hitT_temp_4 <= hitT_temp_4_temp; // @[IST2.scala 358:41]
    end
    if (reset) begin // @[IST2.scala 347:55]
      v22_4 <= 128'h0; // @[IST2.scala 347:55]
    end else begin
      v22_4 <= v22_4_temp; // @[IST2.scala 359:49]
    end
    if (reset) begin // @[IST2.scala 348:50]
      ray_o_in_4 <= 96'h0; // @[IST2.scala 348:50]
    end else begin
      ray_o_in_4 <= ray_o_in_4_temp; // @[IST2.scala 361:40]
    end
    if (reset) begin // @[IST2.scala 349:50]
      ray_d_in_4 <= 96'h0; // @[IST2.scala 349:50]
    end else begin
      ray_d_in_4 <= ray_d_in_4_temp; // @[IST2.scala 360:40]
    end
    if (reset) begin // @[IST2.scala 350:50]
      enable_4 <= 1'h0; // @[IST2.scala 350:50]
    end else begin
      enable_4 <= enable_4_temp; // @[IST2.scala 362:42]
    end
    if (reset) begin // @[IST2.scala 351:53]
      break_4 <= 1'h0; // @[IST2.scala 351:53]
    end else begin
      break_4 <= break_4_temp; // @[IST2.scala 363:43]
    end
    if (reset) begin // @[IST2.scala 352:43]
      ray_aabb_1_4 <= 1'h0; // @[IST2.scala 352:43]
    end else begin
      ray_aabb_1_4 <= ray_aabb_1_4_temp; // @[IST2.scala 364:37]
    end
    if (reset) begin // @[IST2.scala 353:43]
      ray_aabb_2_4 <= 1'h0; // @[IST2.scala 353:43]
    end else begin
      ray_aabb_2_4 <= ray_aabb_2_4_temp; // @[IST2.scala 365:37]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  temp_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  temp_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  temp_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  temp_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  temp_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  temp_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  nodeid_ist2_temp_1_temp = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  rayid_ist2_temp_1_temp = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  t_temp_1_temp = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  hitT_temp_1_temp = _RAND_9[31:0];
  _RAND_10 = {4{`RANDOM}};
  v22_1_temp = _RAND_10[127:0];
  _RAND_11 = {3{`RANDOM}};
  ray_o_in_1_temp = _RAND_11[95:0];
  _RAND_12 = {3{`RANDOM}};
  ray_d_in_1_temp = _RAND_12[95:0];
  _RAND_13 = {1{`RANDOM}};
  enable_1_temp = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  break_1_temp = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  ray_aabb_1_temp = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  ray_aabb_2_temp = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  nodeid_ist2_temp_1 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  rayid_ist2_temp_1 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  t_temp_1 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  hitT_temp_1 = _RAND_20[31:0];
  _RAND_21 = {4{`RANDOM}};
  v22_1 = _RAND_21[127:0];
  _RAND_22 = {3{`RANDOM}};
  ray_o_in_1 = _RAND_22[95:0];
  _RAND_23 = {3{`RANDOM}};
  ray_d_in_1 = _RAND_23[95:0];
  _RAND_24 = {1{`RANDOM}};
  enable_1 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  break_1 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  ray_aabb_1 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  ray_aabb_2 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  nodeid_ist2_temp_2_temp = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  rayid_ist2_temp_2_temp = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  t_temp_2_temp = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  hitT_temp_2_temp = _RAND_31[31:0];
  _RAND_32 = {4{`RANDOM}};
  v22_2_temp = _RAND_32[127:0];
  _RAND_33 = {3{`RANDOM}};
  ray_o_in_2_temp = _RAND_33[95:0];
  _RAND_34 = {3{`RANDOM}};
  ray_d_in_2_temp = _RAND_34[95:0];
  _RAND_35 = {1{`RANDOM}};
  enable_2_temp = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  break_2_temp = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  ray_aabb_1_2_temp = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  ray_aabb_2_2_temp = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  temp_6 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  temp_7 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  temp_0_2 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  temp_0_3 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  temp_5_2 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  temp_5_3 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  nodeid_ist2_temp_2 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  rayid_ist2_temp_2 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  t_temp_2 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  hitT_temp_2 = _RAND_48[31:0];
  _RAND_49 = {4{`RANDOM}};
  v22_2 = _RAND_49[127:0];
  _RAND_50 = {3{`RANDOM}};
  ray_o_in_2 = _RAND_50[95:0];
  _RAND_51 = {3{`RANDOM}};
  ray_d_in_2 = _RAND_51[95:0];
  _RAND_52 = {1{`RANDOM}};
  enable_2 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  break_2 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  ray_aabb_1_2 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  ray_aabb_2_2 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  nodeid_ist2_temp_3_temp = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  rayid_ist2_temp_3_temp = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  t_temp_3_temp = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  hitT_temp_3_temp = _RAND_59[31:0];
  _RAND_60 = {4{`RANDOM}};
  v22_3_temp = _RAND_60[127:0];
  _RAND_61 = {3{`RANDOM}};
  ray_o_in_3_temp = _RAND_61[95:0];
  _RAND_62 = {3{`RANDOM}};
  ray_d_in_3_temp = _RAND_62[95:0];
  _RAND_63 = {1{`RANDOM}};
  enable_3_temp = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  break_3_temp = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  ray_aabb_1_3_temp = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  ray_aabb_2_3_temp = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  Ox = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  Dx = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  nodeid_ist2_temp_3 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  rayid_ist2_temp_3 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  t_temp_3 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  hitT_temp_3 = _RAND_72[31:0];
  _RAND_73 = {4{`RANDOM}};
  v22_3 = _RAND_73[127:0];
  _RAND_74 = {3{`RANDOM}};
  ray_o_in_3 = _RAND_74[95:0];
  _RAND_75 = {3{`RANDOM}};
  ray_d_in_3 = _RAND_75[95:0];
  _RAND_76 = {1{`RANDOM}};
  enable_3 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  break_3 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  ray_aabb_1_3 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  ray_aabb_2_3 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  nodeid_ist2_temp_4_temp = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  rayid_ist2_temp_4_temp = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  temp_u = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  t_temp_4_temp = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  hitT_temp_4_temp = _RAND_84[31:0];
  _RAND_85 = {4{`RANDOM}};
  v22_4_temp = _RAND_85[127:0];
  _RAND_86 = {3{`RANDOM}};
  ray_o_in_4_temp = _RAND_86[95:0];
  _RAND_87 = {3{`RANDOM}};
  ray_d_in_4_temp = _RAND_87[95:0];
  _RAND_88 = {1{`RANDOM}};
  enable_4_temp = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  break_4_temp = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  ray_aabb_1_4_temp = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  ray_aabb_2_4_temp = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  nodeid_ist2_temp_4 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  rayid_ist2_temp_4 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  t_temp_4 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  hitT_temp_4 = _RAND_95[31:0];
  _RAND_96 = {4{`RANDOM}};
  v22_4 = _RAND_96[127:0];
  _RAND_97 = {3{`RANDOM}};
  ray_o_in_4 = _RAND_97[95:0];
  _RAND_98 = {3{`RANDOM}};
  ray_d_in_4 = _RAND_98[95:0];
  _RAND_99 = {1{`RANDOM}};
  enable_4 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  break_4 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  ray_aabb_1_4 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  ray_aabb_2_4 = _RAND_102[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IST3(
  input         clock,
  input         reset,
  input         io_enable_IST3,
  input  [31:0] io_nodeid_leaf_3,
  input  [31:0] io_rayid_leaf_3,
  input  [31:0] io_hiT_in,
  input  [31:0] io_t_in,
  input  [31:0] io_v22_in_x,
  input  [31:0] io_v22_in_y,
  input  [31:0] io_v22_in_z,
  input  [31:0] io_v22_in_w,
  input  [31:0] io_ray_o_in_x,
  input  [31:0] io_ray_o_in_y,
  input  [31:0] io_ray_o_in_z,
  input  [31:0] io_ray_d_in_x,
  input  [31:0] io_ray_d_in_y,
  input  [31:0] io_ray_d_in_z,
  input  [31:0] io_u_in,
  input         io_break_in,
  input         io_RAY_AABB_1,
  input         io_RAY_AABB_2,
  output [31:0] io_nodeid_ist3_out,
  output [31:0] io_rayid_ist3_out,
  output [31:0] io_hiT_out,
  output        io_hitT_en,
  output        io_pop_3,
  output [31:0] io_hitIndex,
  output        io_hitIndex_en,
  output        io_break_out,
  output        io_RAY_AABB_1_out,
  output        io_RAY_AABB_2_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
`endif // RANDOMIZE_REG_INIT
  wire  FADD_MUL_16_clock; // @[IST3.scala 70:33]
  wire  FADD_MUL_16_reset; // @[IST3.scala 70:33]
  wire [31:0] FADD_MUL_16_io_a; // @[IST3.scala 70:33]
  wire [31:0] FADD_MUL_16_io_b; // @[IST3.scala 70:33]
  wire [31:0] FADD_MUL_16_io_c; // @[IST3.scala 70:33]
  wire [31:0] FADD_MUL_16_io_out; // @[IST3.scala 70:33]
  wire  FMUL_12_clock; // @[IST3.scala 80:25]
  wire  FMUL_12_reset; // @[IST3.scala 80:25]
  wire [31:0] FMUL_12_io_a; // @[IST3.scala 80:25]
  wire [31:0] FMUL_12_io_b; // @[IST3.scala 80:25]
  wire [31:0] FMUL_12_io_out; // @[IST3.scala 80:25]
  wire  FMUL_13_clock; // @[IST3.scala 89:25]
  wire  FMUL_13_reset; // @[IST3.scala 89:25]
  wire [31:0] FMUL_13_io_a; // @[IST3.scala 89:25]
  wire [31:0] FMUL_13_io_b; // @[IST3.scala 89:25]
  wire [31:0] FMUL_13_io_out; // @[IST3.scala 89:25]
  wire  FMUL_14_clock; // @[IST3.scala 98:25]
  wire  FMUL_14_reset; // @[IST3.scala 98:25]
  wire [31:0] FMUL_14_io_a; // @[IST3.scala 98:25]
  wire [31:0] FMUL_14_io_b; // @[IST3.scala 98:25]
  wire [31:0] FMUL_14_io_out; // @[IST3.scala 98:25]
  wire  FMUL_15_clock; // @[IST3.scala 107:25]
  wire  FMUL_15_reset; // @[IST3.scala 107:25]
  wire [31:0] FMUL_15_io_a; // @[IST3.scala 107:25]
  wire [31:0] FMUL_15_io_b; // @[IST3.scala 107:25]
  wire [31:0] FMUL_15_io_out; // @[IST3.scala 107:25]
  wire  FMUL_16_clock; // @[IST3.scala 116:25]
  wire  FMUL_16_reset; // @[IST3.scala 116:25]
  wire [31:0] FMUL_16_io_a; // @[IST3.scala 116:25]
  wire [31:0] FMUL_16_io_b; // @[IST3.scala 116:25]
  wire [31:0] FMUL_16_io_out; // @[IST3.scala 116:25]
  wire  FADD_9_clock; // @[IST3.scala 178:24]
  wire  FADD_9_reset; // @[IST3.scala 178:24]
  wire [31:0] FADD_9_io_a; // @[IST3.scala 178:24]
  wire [31:0] FADD_9_io_b; // @[IST3.scala 178:24]
  wire [31:0] FADD_9_io_out; // @[IST3.scala 178:24]
  wire  FADD_10_clock; // @[IST3.scala 187:25]
  wire  FADD_10_reset; // @[IST3.scala 187:25]
  wire [31:0] FADD_10_io_a; // @[IST3.scala 187:25]
  wire [31:0] FADD_10_io_b; // @[IST3.scala 187:25]
  wire [31:0] FADD_10_io_out; // @[IST3.scala 187:25]
  wire  FADD_11_clock; // @[IST3.scala 238:25]
  wire  FADD_11_reset; // @[IST3.scala 238:25]
  wire [31:0] FADD_11_io_a; // @[IST3.scala 238:25]
  wire [31:0] FADD_11_io_b; // @[IST3.scala 238:25]
  wire [31:0] FADD_11_io_out; // @[IST3.scala 238:25]
  wire  FADD_12_clock; // @[IST3.scala 247:25]
  wire  FADD_12_reset; // @[IST3.scala 247:25]
  wire [31:0] FADD_12_io_a; // @[IST3.scala 247:25]
  wire [31:0] FADD_12_io_b; // @[IST3.scala 247:25]
  wire [31:0] FADD_12_io_out; // @[IST3.scala 247:25]
  wire  FADD_MUL_17_clock; // @[IST3.scala 299:33]
  wire  FADD_MUL_17_reset; // @[IST3.scala 299:33]
  wire [31:0] FADD_MUL_17_io_a; // @[IST3.scala 299:33]
  wire [31:0] FADD_MUL_17_io_b; // @[IST3.scala 299:33]
  wire [31:0] FADD_MUL_17_io_c; // @[IST3.scala 299:33]
  wire [31:0] FADD_MUL_17_io_out; // @[IST3.scala 299:33]
  wire [31:0] FCMP_24_io_a; // @[IST3.scala 350:25]
  wire [31:0] FCMP_24_io_b; // @[IST3.scala 350:25]
  wire  FCMP_24_io_actual_out; // @[IST3.scala 350:25]
  wire  FADD_13_clock; // @[IST3.scala 364:25]
  wire  FADD_13_reset; // @[IST3.scala 364:25]
  wire [31:0] FADD_13_io_a; // @[IST3.scala 364:25]
  wire [31:0] FADD_13_io_b; // @[IST3.scala 364:25]
  wire [31:0] FADD_13_io_out; // @[IST3.scala 364:25]
  wire [31:0] FCMP_25_io_a; // @[IST3.scala 398:25]
  wire [31:0] FCMP_25_io_b; // @[IST3.scala 398:25]
  wire  FCMP_25_io_actual_out; // @[IST3.scala 398:25]
  reg [31:0] temp_0; // @[IST3.scala 44:33]
  reg [31:0] temp_1; // @[IST3.scala 45:33]
  reg [31:0] temp_2; // @[IST3.scala 46:33]
  reg [31:0] temp_3; // @[IST3.scala 47:33]
  reg [31:0] temp_4; // @[IST3.scala 48:33]
  reg [31:0] temp_5; // @[IST3.scala 49:33]
  reg [31:0] nodeid_ist3_temp_1_temp; // @[IST3.scala 51:42]
  reg [31:0] rayid_ist3_temp_1_temp; // @[IST3.scala 52:46]
  reg [31:0] t_temp_1_temp; // @[IST3.scala 53:56]
  reg [31:0] u_temp_1_temp; // @[IST3.scala 54:54]
  reg [31:0] hitT_temp_1_temp; // @[IST3.scala 55:52]
  reg  enable_1_temp; // @[IST3.scala 56:55]
  reg  break_1_temp; // @[IST3.scala 57:56]
  reg  ray_aabb_1_temp; // @[IST3.scala 58:51]
  reg  ray_aabb_2_temp; // @[IST3.scala 59:51]
  reg [31:0] nodeid_ist3_temp_1; // @[IST3.scala 126:37]
  reg [31:0] rayid_ist3_temp_1; // @[IST3.scala 127:41]
  reg [31:0] t_temp_1; // @[IST3.scala 128:51]
  reg [31:0] u_temp_1; // @[IST3.scala 129:49]
  reg [31:0] hitT_temp_1; // @[IST3.scala 130:47]
  reg  enable_1; // @[IST3.scala 131:50]
  reg  break_1; // @[IST3.scala 132:51]
  reg  ray_aabb_1; // @[IST3.scala 133:46]
  reg  ray_aabb_2; // @[IST3.scala 134:46]
  reg [31:0] nodeid_ist3_temp_2_temp; // @[IST3.scala 145:43]
  reg [31:0] rayid_ist3_temp_2_temp; // @[IST3.scala 146:46]
  reg [31:0] t_temp_2_temp; // @[IST3.scala 147:56]
  reg [31:0] u_temp_2_temp; // @[IST3.scala 148:55]
  reg [31:0] hitT_temp_2_temp; // @[IST3.scala 149:52]
  reg  enable_2_temp; // @[IST3.scala 150:55]
  reg  break_2_temp; // @[IST3.scala 151:56]
  reg  ray_aabb_1_2_temp; // @[IST3.scala 152:48]
  reg  ray_aabb_2_2_temp; // @[IST3.scala 153:48]
  reg [31:0] temp_6; // @[IST3.scala 164:50]
  reg [31:0] temp_7; // @[IST3.scala 165:50]
  reg [31:0] temp_0_2; // @[IST3.scala 166:47]
  reg [31:0] temp_0_3; // @[IST3.scala 167:47]
  reg [31:0] temp_5_2; // @[IST3.scala 168:46]
  reg [31:0] temp_5_3; // @[IST3.scala 169:46]
  reg [31:0] nodeid_ist3_temp_2; // @[IST3.scala 196:38]
  reg [31:0] rayid_ist3_temp_2; // @[IST3.scala 197:41]
  reg [31:0] t_temp_2; // @[IST3.scala 198:51]
  reg [31:0] u_temp_2; // @[IST3.scala 199:50]
  reg [31:0] hitT_temp_2; // @[IST3.scala 200:47]
  reg  enable_2; // @[IST3.scala 201:50]
  reg  break_2; // @[IST3.scala 202:51]
  reg  ray_aabb_1_2; // @[IST3.scala 203:44]
  reg  ray_aabb_2_2; // @[IST3.scala 204:43]
  reg [31:0] nodeid_ist3_temp_3_temp; // @[IST3.scala 217:43]
  reg [31:0] rayid_ist3_temp_3_temp; // @[IST3.scala 218:46]
  reg [31:0] t_temp_3_temp; // @[IST3.scala 219:56]
  reg [31:0] u_temp_3_temp; // @[IST3.scala 220:55]
  reg [31:0] hitT_temp_3_temp; // @[IST3.scala 221:52]
  reg  enable_3_temp; // @[IST3.scala 222:55]
  reg  break_3_temp; // @[IST3.scala 223:56]
  reg  ray_aabb_1_3_temp; // @[IST3.scala 224:48]
  reg  ray_aabb_2_3_temp; // @[IST3.scala 225:48]
  reg [31:0] Oy; // @[IST3.scala 235:58]
  reg [31:0] Dy; // @[IST3.scala 236:58]
  reg [31:0] nodeid_ist3_temp_3; // @[IST3.scala 258:38]
  reg [31:0] rayid_ist3_temp_3; // @[IST3.scala 259:41]
  reg [31:0] t_temp_3; // @[IST3.scala 260:51]
  reg [31:0] u_temp_3; // @[IST3.scala 261:50]
  reg [31:0] hitT_temp_3; // @[IST3.scala 262:47]
  reg  enable_3; // @[IST3.scala 263:50]
  reg  break_3; // @[IST3.scala 264:51]
  reg  ray_aabb_1_3; // @[IST3.scala 265:43]
  reg  ray_aabb_2_3; // @[IST3.scala 266:43]
  reg [31:0] nodeid_ist3_temp_4_temp; // @[IST3.scala 279:47]
  reg [31:0] rayid_ist3_temp_4_temp; // @[IST3.scala 280:50]
  reg [31:0] t_temp_4_temp; // @[IST3.scala 281:60]
  reg [31:0] u_temp_4_temp; // @[IST3.scala 282:59]
  reg [31:0] hitT_temp_4_temp; // @[IST3.scala 283:56]
  reg  enable_4_temp; // @[IST3.scala 284:59]
  reg  break_4_temp; // @[IST3.scala 285:60]
  reg  ray_aabb_1_4_temp; // @[IST3.scala 286:52]
  reg  ray_aabb_2_4_temp; // @[IST3.scala 287:52]
  reg [31:0] temp_v; // @[IST3.scala 297:67]
  reg [31:0] nodeid_ist3_temp_4; // @[IST3.scala 309:42]
  reg [31:0] rayid_ist3_temp_4; // @[IST3.scala 310:45]
  reg [31:0] t_temp_4; // @[IST3.scala 311:55]
  reg [31:0] u_temp_4; // @[IST3.scala 312:54]
  reg [31:0] hitT_temp_4; // @[IST3.scala 313:51]
  reg  enable_4; // @[IST3.scala 314:54]
  reg  break_4; // @[IST3.scala 315:55]
  reg  ray_aabb_1_4; // @[IST3.scala 316:47]
  reg  ray_aabb_2_4; // @[IST3.scala 317:47]
  reg [31:0] u_add_v; // @[IST3.scala 331:52]
  reg [31:0] nodeid_ist3_temp_5_temp; // @[IST3.scala 332:43]
  reg [31:0] rayid_ist3_temp_5_temp; // @[IST3.scala 333:46]
  reg [31:0] t_temp_5_temp; // @[IST3.scala 334:56]
  reg  v_cmp_0_0; // @[IST3.scala 335:61]
  reg [31:0] hitT_temp_5_temp; // @[IST3.scala 336:52]
  reg  enable_5_temp; // @[IST3.scala 337:55]
  reg  break_5_temp; // @[IST3.scala 339:56]
  reg  ray_aabb_1_5_temp; // @[IST3.scala 340:48]
  reg  ray_aabb_2_5_temp; // @[IST3.scala 341:48]
  wire  _T = FCMP_24_io_actual_out > 1'h0; // @[IST3.scala 355:36]
  reg  v_cmp_0; // @[IST3.scala 361:52]
  reg [31:0] nodeid_ist3_temp_5; // @[IST3.scala 377:38]
  reg [31:0] rayid_ist3_temp_5; // @[IST3.scala 378:41]
  reg [31:0] t_temp_5; // @[IST3.scala 379:51]
  reg [31:0] hitT_temp_5; // @[IST3.scala 382:47]
  reg  enable_5; // @[IST3.scala 383:50]
  reg  break_5; // @[IST3.scala 385:51]
  reg  ray_aabb_1_5; // @[IST3.scala 386:43]
  reg  ray_aabb_2_5; // @[IST3.scala 387:43]
  wire  _T_3 = FCMP_25_io_actual_out & enable_5; // @[IST3.scala 403:43]
  wire  _T_5 = FCMP_25_io_actual_out & enable_5 & v_cmp_0; // @[IST3.scala 403:61]
  wire  _T_6 = ~break_5; // @[IST3.scala 403:90]
  wire  _T_10 = ~FCMP_25_io_actual_out & enable_5; // @[IST3.scala 411:49]
  wire  _T_12 = ~FCMP_25_io_actual_out & enable_5 & v_cmp_0; // @[IST3.scala 411:67]
  wire  _T_18 = ~v_cmp_0; // @[IST3.scala 419:78]
  wire  _T_19 = _T_10 & ~v_cmp_0; // @[IST3.scala 419:67]
  wire  _T_26 = _T_3 & _T_18; // @[IST3.scala 427:67]
  wire  _T_28 = _T_3 & _T_18 & _T_6; // @[IST3.scala 427:86]
  wire  _T_35 = _T_5 & break_5; // @[IST3.scala 435:86]
  wire  _T_56 = _T_26 & break_5; // @[IST3.scala 459:86]
  wire [31:0] _GEN_1 = _T_26 & break_5 ? hitT_temp_5 : 32'h0; // @[IST3.scala 459:104 IST3.scala 460:45 IST3.scala 468:45]
  wire [32:0] _GEN_2 = _T_26 & break_5 ? $signed(33'shbf800000) : $signed(33'sh0); // @[IST3.scala 459:104 IST3.scala 461:45 IST3.scala 469:45]
  wire [31:0] _GEN_4 = _T_26 & break_5 ? rayid_ist3_temp_5 : 32'h0; // @[IST3.scala 459:104 IST3.scala 463:38 IST3.scala 471:38]
  wire [31:0] _GEN_6 = _T_19 & break_5 ? hitT_temp_5 : _GEN_1; // @[IST3.scala 451:104 IST3.scala 452:45]
  wire [32:0] _GEN_7 = _T_19 & break_5 ? $signed(33'shbf800000) : $signed(_GEN_2); // @[IST3.scala 451:104 IST3.scala 453:45]
  wire [31:0] _GEN_9 = _T_19 & break_5 ? rayid_ist3_temp_5 : _GEN_4; // @[IST3.scala 451:104 IST3.scala 455:38]
  wire  _GEN_10 = _T_19 & break_5 | _T_56; // @[IST3.scala 451:104 IST3.scala 458:41]
  wire [31:0] _GEN_11 = _T_12 & break_5 ? hitT_temp_5 : _GEN_6; // @[IST3.scala 443:104 IST3.scala 444:45]
  wire [32:0] _GEN_12 = _T_12 & break_5 ? $signed(33'shbf800000) : $signed(_GEN_7); // @[IST3.scala 443:104 IST3.scala 445:45]
  wire [31:0] _GEN_14 = _T_12 & break_5 ? rayid_ist3_temp_5 : _GEN_9; // @[IST3.scala 443:104 IST3.scala 447:38]
  wire  _GEN_15 = _T_12 & break_5 | _GEN_10; // @[IST3.scala 443:104 IST3.scala 450:41]
  wire [31:0] _GEN_16 = _T_5 & break_5 ? t_temp_5 : _GEN_11; // @[IST3.scala 435:104 IST3.scala 436:45]
  wire [32:0] _GEN_17 = _T_5 & break_5 ? $signed({{1{nodeid_ist3_temp_5[31]}},nodeid_ist3_temp_5}) : $signed(_GEN_12); // @[IST3.scala 435:104 IST3.scala 437:45]
  wire [31:0] _GEN_19 = _T_5 & break_5 ? rayid_ist3_temp_5 : _GEN_14; // @[IST3.scala 435:104 IST3.scala 439:38]
  wire  _GEN_21 = _T_5 & break_5 | _GEN_15; // @[IST3.scala 435:104 IST3.scala 442:41]
  wire [31:0] _GEN_22 = _T_3 & _T_18 & _T_6 ? hitT_temp_5 : _GEN_16; // @[IST3.scala 427:104 IST3.scala 428:45]
  wire [32:0] _GEN_23 = _T_3 & _T_18 & _T_6 ? $signed(33'shbf800000) : $signed(_GEN_17); // @[IST3.scala 427:104 IST3.scala 429:45]
  wire [31:0] _GEN_25 = _T_3 & _T_18 & _T_6 ? rayid_ist3_temp_5 : _GEN_19; // @[IST3.scala 427:104 IST3.scala 431:38]
  wire  _GEN_26 = _T_3 & _T_18 & _T_6 ? 1'h0 : _T_35; // @[IST3.scala 427:104 IST3.scala 432:45]
  wire  _GEN_27 = _T_3 & _T_18 & _T_6 ? 1'h0 : _GEN_21; // @[IST3.scala 427:104 IST3.scala 434:41]
  wire [31:0] _GEN_28 = _T_10 & ~v_cmp_0 & _T_6 ? hitT_temp_5 : _GEN_22; // @[IST3.scala 419:104 IST3.scala 420:45]
  wire [32:0] _GEN_29 = _T_10 & ~v_cmp_0 & _T_6 ? $signed(33'shbf800000) : $signed(_GEN_23); // @[IST3.scala 419:104 IST3.scala 421:45]
  wire  _GEN_30 = _T_10 & ~v_cmp_0 & _T_6 | _T_28; // @[IST3.scala 419:104 IST3.scala 422:46]
  wire [31:0] _GEN_31 = _T_10 & ~v_cmp_0 & _T_6 ? rayid_ist3_temp_5 : _GEN_25; // @[IST3.scala 419:104 IST3.scala 423:38]
  wire  _GEN_32 = _T_10 & ~v_cmp_0 & _T_6 ? 1'h0 : _GEN_26; // @[IST3.scala 419:104 IST3.scala 424:45]
  wire  _GEN_33 = _T_10 & ~v_cmp_0 & _T_6 ? 1'h0 : _GEN_27; // @[IST3.scala 419:104 IST3.scala 426:41]
  wire [31:0] _GEN_34 = ~FCMP_25_io_actual_out & enable_5 & v_cmp_0 & _T_6 ? hitT_temp_5 : _GEN_28; // @[IST3.scala 411:104 IST3.scala 412:45]
  wire [32:0] _GEN_35 = ~FCMP_25_io_actual_out & enable_5 & v_cmp_0 & _T_6 ? $signed(33'shbf800000) : $signed(_GEN_29); // @[IST3.scala 411:104 IST3.scala 413:45]
  wire  _GEN_36 = ~FCMP_25_io_actual_out & enable_5 & v_cmp_0 & _T_6 | _GEN_30; // @[IST3.scala 411:104 IST3.scala 414:46]
  wire [31:0] _GEN_37 = ~FCMP_25_io_actual_out & enable_5 & v_cmp_0 & _T_6 ? rayid_ist3_temp_5 : _GEN_31; // @[IST3.scala 411:104 IST3.scala 415:38]
  wire  _GEN_38 = ~FCMP_25_io_actual_out & enable_5 & v_cmp_0 & _T_6 ? 1'h0 : _GEN_32; // @[IST3.scala 411:104 IST3.scala 416:45]
  wire  _GEN_39 = ~FCMP_25_io_actual_out & enable_5 & v_cmp_0 & _T_6 ? 1'h0 : _GEN_33; // @[IST3.scala 411:104 IST3.scala 418:41]
  wire [32:0] _GEN_41 = FCMP_25_io_actual_out & enable_5 & v_cmp_0 & ~break_5 ? $signed({{1{nodeid_ist3_temp_5[31]}},
    nodeid_ist3_temp_5}) : $signed(_GEN_35); // @[IST3.scala 403:98 IST3.scala 405:45]
  MY_MULADD FADD_MUL_16 ( // @[IST3.scala 70:33]
    .clock(FADD_MUL_16_clock),
    .reset(FADD_MUL_16_reset),
    .io_a(FADD_MUL_16_io_a),
    .io_b(FADD_MUL_16_io_b),
    .io_c(FADD_MUL_16_io_c),
    .io_out(FADD_MUL_16_io_out)
  );
  MY_MUL FMUL_12 ( // @[IST3.scala 80:25]
    .clock(FMUL_12_clock),
    .reset(FMUL_12_reset),
    .io_a(FMUL_12_io_a),
    .io_b(FMUL_12_io_b),
    .io_out(FMUL_12_io_out)
  );
  MY_MUL FMUL_13 ( // @[IST3.scala 89:25]
    .clock(FMUL_13_clock),
    .reset(FMUL_13_reset),
    .io_a(FMUL_13_io_a),
    .io_b(FMUL_13_io_b),
    .io_out(FMUL_13_io_out)
  );
  MY_MUL FMUL_14 ( // @[IST3.scala 98:25]
    .clock(FMUL_14_clock),
    .reset(FMUL_14_reset),
    .io_a(FMUL_14_io_a),
    .io_b(FMUL_14_io_b),
    .io_out(FMUL_14_io_out)
  );
  MY_MUL FMUL_15 ( // @[IST3.scala 107:25]
    .clock(FMUL_15_clock),
    .reset(FMUL_15_reset),
    .io_a(FMUL_15_io_a),
    .io_b(FMUL_15_io_b),
    .io_out(FMUL_15_io_out)
  );
  MY_MUL FMUL_16 ( // @[IST3.scala 116:25]
    .clock(FMUL_16_clock),
    .reset(FMUL_16_reset),
    .io_a(FMUL_16_io_a),
    .io_b(FMUL_16_io_b),
    .io_out(FMUL_16_io_out)
  );
  MY_ADD FADD_9 ( // @[IST3.scala 178:24]
    .clock(FADD_9_clock),
    .reset(FADD_9_reset),
    .io_a(FADD_9_io_a),
    .io_b(FADD_9_io_b),
    .io_out(FADD_9_io_out)
  );
  MY_ADD FADD_10 ( // @[IST3.scala 187:25]
    .clock(FADD_10_clock),
    .reset(FADD_10_reset),
    .io_a(FADD_10_io_a),
    .io_b(FADD_10_io_b),
    .io_out(FADD_10_io_out)
  );
  MY_ADD FADD_11 ( // @[IST3.scala 238:25]
    .clock(FADD_11_clock),
    .reset(FADD_11_reset),
    .io_a(FADD_11_io_a),
    .io_b(FADD_11_io_b),
    .io_out(FADD_11_io_out)
  );
  MY_ADD FADD_12 ( // @[IST3.scala 247:25]
    .clock(FADD_12_clock),
    .reset(FADD_12_reset),
    .io_a(FADD_12_io_a),
    .io_b(FADD_12_io_b),
    .io_out(FADD_12_io_out)
  );
  MY_MULADD FADD_MUL_17 ( // @[IST3.scala 299:33]
    .clock(FADD_MUL_17_clock),
    .reset(FADD_MUL_17_reset),
    .io_a(FADD_MUL_17_io_a),
    .io_b(FADD_MUL_17_io_b),
    .io_c(FADD_MUL_17_io_c),
    .io_out(FADD_MUL_17_io_out)
  );
  ValExec_CompareRecF32_lt FCMP_24 ( // @[IST3.scala 350:25]
    .io_a(FCMP_24_io_a),
    .io_b(FCMP_24_io_b),
    .io_actual_out(FCMP_24_io_actual_out)
  );
  MY_ADD FADD_13 ( // @[IST3.scala 364:25]
    .clock(FADD_13_clock),
    .reset(FADD_13_reset),
    .io_a(FADD_13_io_a),
    .io_b(FADD_13_io_b),
    .io_out(FADD_13_io_out)
  );
  ValExec_CompareRecF32_le FCMP_25 ( // @[IST3.scala 398:25]
    .io_a(FCMP_25_io_a),
    .io_b(FCMP_25_io_b),
    .io_actual_out(FCMP_25_io_actual_out)
  );
  assign io_nodeid_ist3_out = nodeid_ist3_temp_5; // @[IST3.scala 397:37]
  assign io_rayid_ist3_out = FCMP_25_io_actual_out & enable_5 & v_cmp_0 & ~break_5 ? rayid_ist3_temp_5 : _GEN_37; // @[IST3.scala 403:98 IST3.scala 407:38]
  assign io_hiT_out = FCMP_25_io_actual_out & enable_5 & v_cmp_0 & ~break_5 ? t_temp_5 : _GEN_34; // @[IST3.scala 403:98 IST3.scala 404:45]
  assign io_hitT_en = FCMP_25_io_actual_out & enable_5 & v_cmp_0 & ~break_5 | _GEN_38; // @[IST3.scala 403:98 IST3.scala 408:45]
  assign io_pop_3 = FCMP_25_io_actual_out & enable_5 & v_cmp_0 & ~break_5 | _GEN_36; // @[IST3.scala 403:98 IST3.scala 406:46]
  assign io_hitIndex = _GEN_41[31:0];
  assign io_hitIndex_en = FCMP_25_io_actual_out & enable_5 & v_cmp_0 & ~break_5 | _GEN_38; // @[IST3.scala 403:98 IST3.scala 408:45]
  assign io_break_out = FCMP_25_io_actual_out & enable_5 & v_cmp_0 & ~break_5 ? 1'h0 : _GEN_39; // @[IST3.scala 403:98 IST3.scala 410:41]
  assign io_RAY_AABB_1_out = ray_aabb_1_5; // @[IST3.scala 476:37]
  assign io_RAY_AABB_2_out = ray_aabb_2_5; // @[IST3.scala 477:37]
  assign FADD_MUL_16_clock = clock;
  assign FADD_MUL_16_reset = reset;
  assign FADD_MUL_16_io_a = io_ray_o_in_x; // @[IST3.scala 71:26]
  assign FADD_MUL_16_io_b = io_v22_in_x; // @[IST3.scala 72:26]
  assign FADD_MUL_16_io_c = io_v22_in_w; // @[IST3.scala 73:26]
  assign FMUL_12_clock = clock;
  assign FMUL_12_reset = reset;
  assign FMUL_12_io_a = io_ray_o_in_y; // @[IST3.scala 81:22]
  assign FMUL_12_io_b = io_v22_in_y; // @[IST3.scala 82:22]
  assign FMUL_13_clock = clock;
  assign FMUL_13_reset = reset;
  assign FMUL_13_io_a = io_ray_o_in_z; // @[IST3.scala 90:22]
  assign FMUL_13_io_b = io_v22_in_z; // @[IST3.scala 91:22]
  assign FMUL_14_clock = clock;
  assign FMUL_14_reset = reset;
  assign FMUL_14_io_a = io_ray_d_in_x; // @[IST3.scala 99:22]
  assign FMUL_14_io_b = io_v22_in_x; // @[IST3.scala 100:22]
  assign FMUL_15_clock = clock;
  assign FMUL_15_reset = reset;
  assign FMUL_15_io_a = io_ray_d_in_y; // @[IST3.scala 108:22]
  assign FMUL_15_io_b = io_v22_in_y; // @[IST3.scala 109:22]
  assign FMUL_16_clock = clock;
  assign FMUL_16_reset = reset;
  assign FMUL_16_io_a = io_ray_d_in_z; // @[IST3.scala 117:22]
  assign FMUL_16_io_b = io_v22_in_z; // @[IST3.scala 118:22]
  assign FADD_9_clock = clock;
  assign FADD_9_reset = reset;
  assign FADD_9_io_a = temp_1; // @[IST3.scala 179:21]
  assign FADD_9_io_b = temp_2; // @[IST3.scala 180:21]
  assign FADD_10_clock = clock;
  assign FADD_10_reset = reset;
  assign FADD_10_io_a = temp_3; // @[IST3.scala 188:22]
  assign FADD_10_io_b = temp_4; // @[IST3.scala 189:22]
  assign FADD_11_clock = clock;
  assign FADD_11_reset = reset;
  assign FADD_11_io_a = temp_0_3; // @[IST3.scala 239:22]
  assign FADD_11_io_b = temp_6; // @[IST3.scala 240:22]
  assign FADD_12_clock = clock;
  assign FADD_12_reset = reset;
  assign FADD_12_io_a = temp_5_3; // @[IST3.scala 248:22]
  assign FADD_12_io_b = temp_7; // @[IST3.scala 249:22]
  assign FADD_MUL_17_clock = clock;
  assign FADD_MUL_17_reset = reset;
  assign FADD_MUL_17_io_a = t_temp_3; // @[IST3.scala 300:26]
  assign FADD_MUL_17_io_b = Dy; // @[IST3.scala 301:26]
  assign FADD_MUL_17_io_c = Oy; // @[IST3.scala 302:26]
  assign FCMP_24_io_a = 32'h0; // @[IST3.scala 351:22]
  assign FCMP_24_io_b = temp_v; // @[IST3.scala 352:22]
  assign FADD_13_clock = clock;
  assign FADD_13_reset = reset;
  assign FADD_13_io_a = temp_v; // @[IST3.scala 365:22]
  assign FADD_13_io_b = u_temp_4; // @[IST3.scala 366:22]
  assign FCMP_25_io_a = u_add_v; // @[IST3.scala 399:22]
  assign FCMP_25_io_b = 32'h3f800000; // @[IST3.scala 400:22]
  always @(posedge clock) begin
    if (reset) begin // @[IST3.scala 44:33]
      temp_0 <= 32'h0; // @[IST3.scala 44:33]
    end else begin
      temp_0 <= FADD_MUL_16_io_out; // @[IST3.scala 78:42]
    end
    if (reset) begin // @[IST3.scala 45:33]
      temp_1 <= 32'h0; // @[IST3.scala 45:33]
    end else begin
      temp_1 <= FMUL_12_io_out; // @[IST3.scala 87:42]
    end
    if (reset) begin // @[IST3.scala 46:33]
      temp_2 <= 32'h0; // @[IST3.scala 46:33]
    end else begin
      temp_2 <= FMUL_13_io_out; // @[IST3.scala 96:42]
    end
    if (reset) begin // @[IST3.scala 47:33]
      temp_3 <= 32'h0; // @[IST3.scala 47:33]
    end else begin
      temp_3 <= FMUL_14_io_out; // @[IST3.scala 105:42]
    end
    if (reset) begin // @[IST3.scala 48:33]
      temp_4 <= 32'h0; // @[IST3.scala 48:33]
    end else begin
      temp_4 <= FMUL_15_io_out; // @[IST3.scala 114:42]
    end
    if (reset) begin // @[IST3.scala 49:33]
      temp_5 <= 32'h0; // @[IST3.scala 49:33]
    end else begin
      temp_5 <= FMUL_16_io_out; // @[IST3.scala 123:42]
    end
    if (reset) begin // @[IST3.scala 51:42]
      nodeid_ist3_temp_1_temp <= 32'sh0; // @[IST3.scala 51:42]
    end else begin
      nodeid_ist3_temp_1_temp <= io_nodeid_leaf_3; // @[IST3.scala 60:34]
    end
    if (reset) begin // @[IST3.scala 52:46]
      rayid_ist3_temp_1_temp <= 32'h0; // @[IST3.scala 52:46]
    end else begin
      rayid_ist3_temp_1_temp <= io_rayid_leaf_3; // @[IST3.scala 61:37]
    end
    if (reset) begin // @[IST3.scala 53:56]
      t_temp_1_temp <= 32'h0; // @[IST3.scala 53:56]
    end else begin
      t_temp_1_temp <= io_t_in; // @[IST3.scala 62:47]
    end
    if (reset) begin // @[IST3.scala 54:54]
      u_temp_1_temp <= 32'h0; // @[IST3.scala 54:54]
    end else begin
      u_temp_1_temp <= io_u_in; // @[IST3.scala 63:46]
    end
    if (reset) begin // @[IST3.scala 55:52]
      hitT_temp_1_temp <= 32'h0; // @[IST3.scala 55:52]
    end else begin
      hitT_temp_1_temp <= io_hiT_in; // @[IST3.scala 64:43]
    end
    if (reset) begin // @[IST3.scala 56:55]
      enable_1_temp <= 1'h0; // @[IST3.scala 56:55]
    end else begin
      enable_1_temp <= io_enable_IST3; // @[IST3.scala 65:48]
    end
    if (reset) begin // @[IST3.scala 57:56]
      break_1_temp <= 1'h0; // @[IST3.scala 57:56]
    end else begin
      break_1_temp <= io_break_in; // @[IST3.scala 66:50]
    end
    if (reset) begin // @[IST3.scala 58:51]
      ray_aabb_1_temp <= 1'h0; // @[IST3.scala 58:51]
    end else begin
      ray_aabb_1_temp <= io_RAY_AABB_1; // @[IST3.scala 67:45]
    end
    if (reset) begin // @[IST3.scala 59:51]
      ray_aabb_2_temp <= 1'h0; // @[IST3.scala 59:51]
    end else begin
      ray_aabb_2_temp <= io_RAY_AABB_2; // @[IST3.scala 68:45]
    end
    if (reset) begin // @[IST3.scala 126:37]
      nodeid_ist3_temp_1 <= 32'sh0; // @[IST3.scala 126:37]
    end else begin
      nodeid_ist3_temp_1 <= nodeid_ist3_temp_1_temp; // @[IST3.scala 135:29]
    end
    if (reset) begin // @[IST3.scala 127:41]
      rayid_ist3_temp_1 <= 32'h0; // @[IST3.scala 127:41]
    end else begin
      rayid_ist3_temp_1 <= rayid_ist3_temp_1_temp; // @[IST3.scala 136:32]
    end
    if (reset) begin // @[IST3.scala 128:51]
      t_temp_1 <= 32'h0; // @[IST3.scala 128:51]
    end else begin
      t_temp_1 <= t_temp_1_temp; // @[IST3.scala 137:42]
    end
    if (reset) begin // @[IST3.scala 129:49]
      u_temp_1 <= 32'h0; // @[IST3.scala 129:49]
    end else begin
      u_temp_1 <= u_temp_1_temp; // @[IST3.scala 138:41]
    end
    if (reset) begin // @[IST3.scala 130:47]
      hitT_temp_1 <= 32'h0; // @[IST3.scala 130:47]
    end else begin
      hitT_temp_1 <= hitT_temp_1_temp; // @[IST3.scala 139:38]
    end
    if (reset) begin // @[IST3.scala 131:50]
      enable_1 <= 1'h0; // @[IST3.scala 131:50]
    end else begin
      enable_1 <= enable_1_temp; // @[IST3.scala 140:43]
    end
    if (reset) begin // @[IST3.scala 132:51]
      break_1 <= 1'h0; // @[IST3.scala 132:51]
    end else begin
      break_1 <= break_1_temp; // @[IST3.scala 141:45]
    end
    if (reset) begin // @[IST3.scala 133:46]
      ray_aabb_1 <= 1'h0; // @[IST3.scala 133:46]
    end else begin
      ray_aabb_1 <= ray_aabb_1_temp; // @[IST3.scala 142:40]
    end
    if (reset) begin // @[IST3.scala 134:46]
      ray_aabb_2 <= 1'h0; // @[IST3.scala 134:46]
    end else begin
      ray_aabb_2 <= ray_aabb_2_temp; // @[IST3.scala 143:40]
    end
    if (reset) begin // @[IST3.scala 145:43]
      nodeid_ist3_temp_2_temp <= 32'sh0; // @[IST3.scala 145:43]
    end else begin
      nodeid_ist3_temp_2_temp <= nodeid_ist3_temp_1; // @[IST3.scala 154:34]
    end
    if (reset) begin // @[IST3.scala 146:46]
      rayid_ist3_temp_2_temp <= 32'h0; // @[IST3.scala 146:46]
    end else begin
      rayid_ist3_temp_2_temp <= rayid_ist3_temp_1; // @[IST3.scala 155:37]
    end
    if (reset) begin // @[IST3.scala 147:56]
      t_temp_2_temp <= 32'h0; // @[IST3.scala 147:56]
    end else begin
      t_temp_2_temp <= t_temp_1; // @[IST3.scala 156:46]
    end
    if (reset) begin // @[IST3.scala 148:55]
      u_temp_2_temp <= 32'h0; // @[IST3.scala 148:55]
    end else begin
      u_temp_2_temp <= u_temp_1; // @[IST3.scala 157:45]
    end
    if (reset) begin // @[IST3.scala 149:52]
      hitT_temp_2_temp <= 32'h0; // @[IST3.scala 149:52]
    end else begin
      hitT_temp_2_temp <= hitT_temp_1; // @[IST3.scala 158:43]
    end
    if (reset) begin // @[IST3.scala 150:55]
      enable_2_temp <= 1'h0; // @[IST3.scala 150:55]
    end else begin
      enable_2_temp <= enable_1; // @[IST3.scala 159:47]
    end
    if (reset) begin // @[IST3.scala 151:56]
      break_2_temp <= 1'h0; // @[IST3.scala 151:56]
    end else begin
      break_2_temp <= break_1; // @[IST3.scala 160:48]
    end
    if (reset) begin // @[IST3.scala 152:48]
      ray_aabb_1_2_temp <= 1'h0; // @[IST3.scala 152:48]
    end else begin
      ray_aabb_1_2_temp <= ray_aabb_1; // @[IST3.scala 161:40]
    end
    if (reset) begin // @[IST3.scala 153:48]
      ray_aabb_2_2_temp <= 1'h0; // @[IST3.scala 153:48]
    end else begin
      ray_aabb_2_2_temp <= ray_aabb_2; // @[IST3.scala 162:40]
    end
    if (reset) begin // @[IST3.scala 164:50]
      temp_6 <= 32'h0; // @[IST3.scala 164:50]
    end else begin
      temp_6 <= FADD_9_io_out; // @[IST3.scala 185:26]
    end
    if (reset) begin // @[IST3.scala 165:50]
      temp_7 <= 32'h0; // @[IST3.scala 165:50]
    end else begin
      temp_7 <= FADD_10_io_out; // @[IST3.scala 194:26]
    end
    if (reset) begin // @[IST3.scala 166:47]
      temp_0_2 <= 32'h0; // @[IST3.scala 166:47]
    end else begin
      temp_0_2 <= temp_0; // @[IST3.scala 175:41]
    end
    if (reset) begin // @[IST3.scala 167:47]
      temp_0_3 <= 32'h0; // @[IST3.scala 167:47]
    end else begin
      temp_0_3 <= temp_0_2; // @[IST3.scala 172:41]
    end
    if (reset) begin // @[IST3.scala 168:46]
      temp_5_2 <= 32'h0; // @[IST3.scala 168:46]
    end else begin
      temp_5_2 <= temp_5; // @[IST3.scala 176:41]
    end
    if (reset) begin // @[IST3.scala 169:46]
      temp_5_3 <= 32'h0; // @[IST3.scala 169:46]
    end else begin
      temp_5_3 <= temp_5_2; // @[IST3.scala 174:41]
    end
    if (reset) begin // @[IST3.scala 196:38]
      nodeid_ist3_temp_2 <= 32'sh0; // @[IST3.scala 196:38]
    end else begin
      nodeid_ist3_temp_2 <= nodeid_ist3_temp_2_temp; // @[IST3.scala 205:29]
    end
    if (reset) begin // @[IST3.scala 197:41]
      rayid_ist3_temp_2 <= 32'h0; // @[IST3.scala 197:41]
    end else begin
      rayid_ist3_temp_2 <= rayid_ist3_temp_2_temp; // @[IST3.scala 206:32]
    end
    if (reset) begin // @[IST3.scala 198:51]
      t_temp_2 <= 32'h0; // @[IST3.scala 198:51]
    end else begin
      t_temp_2 <= t_temp_2_temp; // @[IST3.scala 207:41]
    end
    if (reset) begin // @[IST3.scala 199:50]
      u_temp_2 <= 32'h0; // @[IST3.scala 199:50]
    end else begin
      u_temp_2 <= u_temp_2_temp; // @[IST3.scala 208:40]
    end
    if (reset) begin // @[IST3.scala 200:47]
      hitT_temp_2 <= 32'h0; // @[IST3.scala 200:47]
    end else begin
      hitT_temp_2 <= hitT_temp_2_temp; // @[IST3.scala 209:38]
    end
    if (reset) begin // @[IST3.scala 201:50]
      enable_2 <= 1'h0; // @[IST3.scala 201:50]
    end else begin
      enable_2 <= enable_2_temp; // @[IST3.scala 210:42]
    end
    if (reset) begin // @[IST3.scala 202:51]
      break_2 <= 1'h0; // @[IST3.scala 202:51]
    end else begin
      break_2 <= break_2_temp; // @[IST3.scala 211:43]
    end
    if (reset) begin // @[IST3.scala 203:44]
      ray_aabb_1_2 <= 1'h0; // @[IST3.scala 203:44]
    end else begin
      ray_aabb_1_2 <= ray_aabb_1_2_temp; // @[IST3.scala 212:37]
    end
    if (reset) begin // @[IST3.scala 204:43]
      ray_aabb_2_2 <= 1'h0; // @[IST3.scala 204:43]
    end else begin
      ray_aabb_2_2 <= ray_aabb_2_2_temp; // @[IST3.scala 213:37]
    end
    if (reset) begin // @[IST3.scala 217:43]
      nodeid_ist3_temp_3_temp <= 32'sh0; // @[IST3.scala 217:43]
    end else begin
      nodeid_ist3_temp_3_temp <= nodeid_ist3_temp_2; // @[IST3.scala 226:37]
    end
    if (reset) begin // @[IST3.scala 218:46]
      rayid_ist3_temp_3_temp <= 32'h0; // @[IST3.scala 218:46]
    end else begin
      rayid_ist3_temp_3_temp <= rayid_ist3_temp_2; // @[IST3.scala 227:40]
    end
    if (reset) begin // @[IST3.scala 219:56]
      t_temp_3_temp <= 32'h0; // @[IST3.scala 219:56]
    end else begin
      t_temp_3_temp <= t_temp_2; // @[IST3.scala 228:50]
    end
    if (reset) begin // @[IST3.scala 220:55]
      u_temp_3_temp <= 32'h0; // @[IST3.scala 220:55]
    end else begin
      u_temp_3_temp <= u_temp_2; // @[IST3.scala 229:49]
    end
    if (reset) begin // @[IST3.scala 221:52]
      hitT_temp_3_temp <= 32'h0; // @[IST3.scala 221:52]
    end else begin
      hitT_temp_3_temp <= hitT_temp_2; // @[IST3.scala 230:46]
    end
    if (reset) begin // @[IST3.scala 222:55]
      enable_3_temp <= 1'h0; // @[IST3.scala 222:55]
    end else begin
      enable_3_temp <= enable_2; // @[IST3.scala 231:51]
    end
    if (reset) begin // @[IST3.scala 223:56]
      break_3_temp <= 1'h0; // @[IST3.scala 223:56]
    end else begin
      break_3_temp <= break_2; // @[IST3.scala 232:53]
    end
    if (reset) begin // @[IST3.scala 224:48]
      ray_aabb_1_3_temp <= 1'h0; // @[IST3.scala 224:48]
    end else begin
      ray_aabb_1_3_temp <= ray_aabb_1_2; // @[IST3.scala 233:45]
    end
    if (reset) begin // @[IST3.scala 225:48]
      ray_aabb_2_3_temp <= 1'h0; // @[IST3.scala 225:48]
    end else begin
      ray_aabb_2_3_temp <= ray_aabb_2_2; // @[IST3.scala 234:45]
    end
    if (reset) begin // @[IST3.scala 235:58]
      Oy <= 32'h0; // @[IST3.scala 235:58]
    end else begin
      Oy <= FADD_11_io_out; // @[IST3.scala 245:26]
    end
    if (reset) begin // @[IST3.scala 236:58]
      Dy <= 32'h0; // @[IST3.scala 236:58]
    end else begin
      Dy <= FADD_12_io_out; // @[IST3.scala 254:26]
    end
    if (reset) begin // @[IST3.scala 258:38]
      nodeid_ist3_temp_3 <= 32'sh0; // @[IST3.scala 258:38]
    end else begin
      nodeid_ist3_temp_3 <= nodeid_ist3_temp_3_temp; // @[IST3.scala 267:32]
    end
    if (reset) begin // @[IST3.scala 259:41]
      rayid_ist3_temp_3 <= 32'h0; // @[IST3.scala 259:41]
    end else begin
      rayid_ist3_temp_3 <= rayid_ist3_temp_3_temp; // @[IST3.scala 268:35]
    end
    if (reset) begin // @[IST3.scala 260:51]
      t_temp_3 <= 32'h0; // @[IST3.scala 260:51]
    end else begin
      t_temp_3 <= t_temp_3_temp; // @[IST3.scala 269:45]
    end
    if (reset) begin // @[IST3.scala 261:50]
      u_temp_3 <= 32'h0; // @[IST3.scala 261:50]
    end else begin
      u_temp_3 <= u_temp_3_temp; // @[IST3.scala 270:44]
    end
    if (reset) begin // @[IST3.scala 262:47]
      hitT_temp_3 <= 32'h0; // @[IST3.scala 262:47]
    end else begin
      hitT_temp_3 <= hitT_temp_3_temp; // @[IST3.scala 271:41]
    end
    if (reset) begin // @[IST3.scala 263:50]
      enable_3 <= 1'h0; // @[IST3.scala 263:50]
    end else begin
      enable_3 <= enable_3_temp; // @[IST3.scala 272:43]
    end
    if (reset) begin // @[IST3.scala 264:51]
      break_3 <= 1'h0; // @[IST3.scala 264:51]
    end else begin
      break_3 <= break_3_temp; // @[IST3.scala 273:45]
    end
    if (reset) begin // @[IST3.scala 265:43]
      ray_aabb_1_3 <= 1'h0; // @[IST3.scala 265:43]
    end else begin
      ray_aabb_1_3 <= ray_aabb_1_3_temp; // @[IST3.scala 274:37]
    end
    if (reset) begin // @[IST3.scala 266:43]
      ray_aabb_2_3 <= 1'h0; // @[IST3.scala 266:43]
    end else begin
      ray_aabb_2_3 <= ray_aabb_2_3_temp; // @[IST3.scala 275:37]
    end
    if (reset) begin // @[IST3.scala 279:47]
      nodeid_ist3_temp_4_temp <= 32'sh0; // @[IST3.scala 279:47]
    end else begin
      nodeid_ist3_temp_4_temp <= nodeid_ist3_temp_3; // @[IST3.scala 288:41]
    end
    if (reset) begin // @[IST3.scala 280:50]
      rayid_ist3_temp_4_temp <= 32'h0; // @[IST3.scala 280:50]
    end else begin
      rayid_ist3_temp_4_temp <= rayid_ist3_temp_3; // @[IST3.scala 289:44]
    end
    if (reset) begin // @[IST3.scala 281:60]
      t_temp_4_temp <= 32'h0; // @[IST3.scala 281:60]
    end else begin
      t_temp_4_temp <= t_temp_3; // @[IST3.scala 290:54]
    end
    if (reset) begin // @[IST3.scala 282:59]
      u_temp_4_temp <= 32'h0; // @[IST3.scala 282:59]
    end else begin
      u_temp_4_temp <= u_temp_3; // @[IST3.scala 291:53]
    end
    if (reset) begin // @[IST3.scala 283:56]
      hitT_temp_4_temp <= 32'h0; // @[IST3.scala 283:56]
    end else begin
      hitT_temp_4_temp <= hitT_temp_3; // @[IST3.scala 292:50]
    end
    if (reset) begin // @[IST3.scala 284:59]
      enable_4_temp <= 1'h0; // @[IST3.scala 284:59]
    end else begin
      enable_4_temp <= enable_3; // @[IST3.scala 293:55]
    end
    if (reset) begin // @[IST3.scala 285:60]
      break_4_temp <= 1'h0; // @[IST3.scala 285:60]
    end else begin
      break_4_temp <= break_3; // @[IST3.scala 294:56]
    end
    if (reset) begin // @[IST3.scala 286:52]
      ray_aabb_1_4_temp <= 1'h0; // @[IST3.scala 286:52]
    end else begin
      ray_aabb_1_4_temp <= ray_aabb_1_3; // @[IST3.scala 295:48]
    end
    if (reset) begin // @[IST3.scala 287:52]
      ray_aabb_2_4_temp <= 1'h0; // @[IST3.scala 287:52]
    end else begin
      ray_aabb_2_4_temp <= ray_aabb_2_3; // @[IST3.scala 296:48]
    end
    if (reset) begin // @[IST3.scala 297:67]
      temp_v <= 32'h0; // @[IST3.scala 297:67]
    end else begin
      temp_v <= FADD_MUL_17_io_out; // @[IST3.scala 307:42]
    end
    if (reset) begin // @[IST3.scala 309:42]
      nodeid_ist3_temp_4 <= 32'sh0; // @[IST3.scala 309:42]
    end else begin
      nodeid_ist3_temp_4 <= nodeid_ist3_temp_4_temp; // @[IST3.scala 318:36]
    end
    if (reset) begin // @[IST3.scala 310:45]
      rayid_ist3_temp_4 <= 32'h0; // @[IST3.scala 310:45]
    end else begin
      rayid_ist3_temp_4 <= rayid_ist3_temp_4_temp; // @[IST3.scala 319:39]
    end
    if (reset) begin // @[IST3.scala 311:55]
      t_temp_4 <= 32'h0; // @[IST3.scala 311:55]
    end else begin
      t_temp_4 <= t_temp_4_temp; // @[IST3.scala 320:49]
    end
    if (reset) begin // @[IST3.scala 312:54]
      u_temp_4 <= 32'h0; // @[IST3.scala 312:54]
    end else begin
      u_temp_4 <= u_temp_4_temp; // @[IST3.scala 321:48]
    end
    if (reset) begin // @[IST3.scala 313:51]
      hitT_temp_4 <= 32'h0; // @[IST3.scala 313:51]
    end else begin
      hitT_temp_4 <= hitT_temp_4_temp; // @[IST3.scala 322:45]
    end
    if (reset) begin // @[IST3.scala 314:54]
      enable_4 <= 1'h0; // @[IST3.scala 314:54]
    end else begin
      enable_4 <= enable_4_temp; // @[IST3.scala 323:50]
    end
    if (reset) begin // @[IST3.scala 315:55]
      break_4 <= 1'h0; // @[IST3.scala 315:55]
    end else begin
      break_4 <= break_4_temp; // @[IST3.scala 324:51]
    end
    if (reset) begin // @[IST3.scala 316:47]
      ray_aabb_1_4 <= 1'h0; // @[IST3.scala 316:47]
    end else begin
      ray_aabb_1_4 <= ray_aabb_1_4_temp; // @[IST3.scala 325:44]
    end
    if (reset) begin // @[IST3.scala 317:47]
      ray_aabb_2_4 <= 1'h0; // @[IST3.scala 317:47]
    end else begin
      ray_aabb_2_4 <= ray_aabb_2_4_temp; // @[IST3.scala 326:44]
    end
    if (reset) begin // @[IST3.scala 331:52]
      u_add_v <= 32'h0; // @[IST3.scala 331:52]
    end else begin
      u_add_v <= FADD_13_io_out; // @[IST3.scala 371:25]
    end
    if (reset) begin // @[IST3.scala 332:43]
      nodeid_ist3_temp_5_temp <= 32'sh0; // @[IST3.scala 332:43]
    end else begin
      nodeid_ist3_temp_5_temp <= nodeid_ist3_temp_4; // @[IST3.scala 342:37]
    end
    if (reset) begin // @[IST3.scala 333:46]
      rayid_ist3_temp_5_temp <= 32'h0; // @[IST3.scala 333:46]
    end else begin
      rayid_ist3_temp_5_temp <= rayid_ist3_temp_4; // @[IST3.scala 343:40]
    end
    if (reset) begin // @[IST3.scala 334:56]
      t_temp_5_temp <= 32'h0; // @[IST3.scala 334:56]
    end else begin
      t_temp_5_temp <= t_temp_4; // @[IST3.scala 344:50]
    end
    if (reset) begin // @[IST3.scala 335:61]
      v_cmp_0_0 <= 1'h0; // @[IST3.scala 335:61]
    end else begin
      v_cmp_0_0 <= _T;
    end
    if (reset) begin // @[IST3.scala 336:52]
      hitT_temp_5_temp <= 32'h0; // @[IST3.scala 336:52]
    end else begin
      hitT_temp_5_temp <= hitT_temp_4; // @[IST3.scala 345:46]
    end
    if (reset) begin // @[IST3.scala 337:55]
      enable_5_temp <= 1'h0; // @[IST3.scala 337:55]
    end else begin
      enable_5_temp <= enable_4; // @[IST3.scala 346:51]
    end
    if (reset) begin // @[IST3.scala 339:56]
      break_5_temp <= 1'h0; // @[IST3.scala 339:56]
    end else begin
      break_5_temp <= break_4; // @[IST3.scala 347:52]
    end
    if (reset) begin // @[IST3.scala 340:48]
      ray_aabb_1_5_temp <= 1'h0; // @[IST3.scala 340:48]
    end else begin
      ray_aabb_1_5_temp <= ray_aabb_1_4; // @[IST3.scala 348:42]
    end
    if (reset) begin // @[IST3.scala 341:48]
      ray_aabb_2_5_temp <= 1'h0; // @[IST3.scala 341:48]
    end else begin
      ray_aabb_2_5_temp <= ray_aabb_2_4; // @[IST3.scala 349:42]
    end
    if (reset) begin // @[IST3.scala 361:52]
      v_cmp_0 <= 1'h0; // @[IST3.scala 361:52]
    end else begin
      v_cmp_0 <= v_cmp_0_0; // @[IST3.scala 362:45]
    end
    if (reset) begin // @[IST3.scala 377:38]
      nodeid_ist3_temp_5 <= 32'sh0; // @[IST3.scala 377:38]
    end else begin
      nodeid_ist3_temp_5 <= nodeid_ist3_temp_5_temp; // @[IST3.scala 389:32]
    end
    if (reset) begin // @[IST3.scala 378:41]
      rayid_ist3_temp_5 <= 32'h0; // @[IST3.scala 378:41]
    end else begin
      rayid_ist3_temp_5 <= rayid_ist3_temp_5_temp; // @[IST3.scala 390:35]
    end
    if (reset) begin // @[IST3.scala 379:51]
      t_temp_5 <= 32'h0; // @[IST3.scala 379:51]
    end else begin
      t_temp_5 <= t_temp_5_temp; // @[IST3.scala 391:45]
    end
    if (reset) begin // @[IST3.scala 382:47]
      hitT_temp_5 <= 32'h0; // @[IST3.scala 382:47]
    end else begin
      hitT_temp_5 <= hitT_temp_5_temp; // @[IST3.scala 392:41]
    end
    if (reset) begin // @[IST3.scala 383:50]
      enable_5 <= 1'h0; // @[IST3.scala 383:50]
    end else begin
      enable_5 <= enable_5_temp; // @[IST3.scala 393:46]
    end
    if (reset) begin // @[IST3.scala 385:51]
      break_5 <= 1'h0; // @[IST3.scala 385:51]
    end else begin
      break_5 <= break_5_temp; // @[IST3.scala 394:47]
    end
    if (reset) begin // @[IST3.scala 386:43]
      ray_aabb_1_5 <= 1'h0; // @[IST3.scala 386:43]
    end else begin
      ray_aabb_1_5 <= ray_aabb_1_5_temp; // @[IST3.scala 395:40]
    end
    if (reset) begin // @[IST3.scala 387:43]
      ray_aabb_2_5 <= 1'h0; // @[IST3.scala 387:43]
    end else begin
      ray_aabb_2_5 <= ray_aabb_2_5_temp; // @[IST3.scala 396:40]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  temp_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  temp_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  temp_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  temp_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  temp_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  temp_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  nodeid_ist3_temp_1_temp = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  rayid_ist3_temp_1_temp = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  t_temp_1_temp = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  u_temp_1_temp = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  hitT_temp_1_temp = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  enable_1_temp = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  break_1_temp = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  ray_aabb_1_temp = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  ray_aabb_2_temp = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  nodeid_ist3_temp_1 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  rayid_ist3_temp_1 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  t_temp_1 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  u_temp_1 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  hitT_temp_1 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  enable_1 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  break_1 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  ray_aabb_1 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  ray_aabb_2 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  nodeid_ist3_temp_2_temp = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  rayid_ist3_temp_2_temp = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  t_temp_2_temp = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  u_temp_2_temp = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  hitT_temp_2_temp = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  enable_2_temp = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  break_2_temp = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  ray_aabb_1_2_temp = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  ray_aabb_2_2_temp = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  temp_6 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  temp_7 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  temp_0_2 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  temp_0_3 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  temp_5_2 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  temp_5_3 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  nodeid_ist3_temp_2 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  rayid_ist3_temp_2 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  t_temp_2 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  u_temp_2 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  hitT_temp_2 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  enable_2 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  break_2 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  ray_aabb_1_2 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  ray_aabb_2_2 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  nodeid_ist3_temp_3_temp = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  rayid_ist3_temp_3_temp = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  t_temp_3_temp = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  u_temp_3_temp = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  hitT_temp_3_temp = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  enable_3_temp = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  break_3_temp = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  ray_aabb_1_3_temp = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  ray_aabb_2_3_temp = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  Oy = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  Dy = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  nodeid_ist3_temp_3 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  rayid_ist3_temp_3 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  t_temp_3 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  u_temp_3 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  hitT_temp_3 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  enable_3 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  break_3 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  ray_aabb_1_3 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  ray_aabb_2_3 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  nodeid_ist3_temp_4_temp = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  rayid_ist3_temp_4_temp = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  t_temp_4_temp = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  u_temp_4_temp = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  hitT_temp_4_temp = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  enable_4_temp = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  break_4_temp = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  ray_aabb_1_4_temp = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  ray_aabb_2_4_temp = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  temp_v = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  nodeid_ist3_temp_4 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  rayid_ist3_temp_4 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  t_temp_4 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  u_temp_4 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  hitT_temp_4 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  enable_4 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  break_4 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  ray_aabb_1_4 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  ray_aabb_2_4 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  u_add_v = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  nodeid_ist3_temp_5_temp = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  rayid_ist3_temp_5_temp = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  t_temp_5_temp = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  v_cmp_0_0 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  hitT_temp_5_temp = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  enable_5_temp = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  break_5_temp = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  ray_aabb_1_5_temp = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  ray_aabb_2_5_temp = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  v_cmp_0 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  nodeid_ist3_temp_5 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  rayid_ist3_temp_5 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  t_temp_5 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  hitT_temp_5 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  enable_5 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  break_5 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  ray_aabb_1_5 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  ray_aabb_2_5 = _RAND_105[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Triangle(
  input         clock,
  input         reset,
  input         io_To_IST0_enable,
  input  [31:0] io_nodeid_leaf,
  input  [31:0] io_rayid_leaf,
  input  [31:0] io_hiT_in,
  input  [31:0] io_v00_in_x,
  input  [31:0] io_v00_in_y,
  input  [31:0] io_v00_in_z,
  input  [31:0] io_v00_in_w,
  input  [31:0] io_v11_in_x,
  input  [31:0] io_v11_in_y,
  input  [31:0] io_v11_in_z,
  input  [31:0] io_v11_in_w,
  input  [31:0] io_v22_in_x,
  input  [31:0] io_v22_in_y,
  input  [31:0] io_v22_in_z,
  input  [31:0] io_v22_in_w,
  input  [31:0] io_ray_o_in_x,
  input  [31:0] io_ray_o_in_y,
  input  [31:0] io_ray_o_in_z,
  input  [31:0] io_ray_d_in_x,
  input  [31:0] io_ray_d_in_y,
  input  [31:0] io_ray_d_in_z,
  input         io_break_in,
  input         io_RAY_AABB_1,
  input         io_RAY_AABB_2,
  output        io_pop_1,
  output        io_break_1,
  output        io_pop_2,
  output        io_break_2,
  output        io_pop_3,
  output        io_break_3,
  output [31:0] io_hiT_out_1,
  output [31:0] io_hiT_out_2,
  output [31:0] io_hiT_out_3,
  output        io_hitT_en,
  output [31:0] io_hitIndex,
  output        io_hitIndex_en,
  output [31:0] io_node_id_out_1,
  output [31:0] io_node_id_out_2,
  output [31:0] io_node_id_out_3,
  output [31:0] io_ray_id_ist1,
  output [31:0] io_ray_id_ist2,
  output [31:0] io_ray_id_ist3,
  output [63:0] io_counter_fdiv,
  output        io_RAY_AABB_1_out_IST1,
  output        io_RAY_AABB_2_out_IST1,
  output        io_RAY_AABB_1_out_IST2,
  output        io_RAY_AABB_2_out_IST2,
  output        io_RAY_AABB_1_out_IST3,
  output        io_RAY_AABB_2_out_IST3
);
  wire  IST0_clock; // @[Triangle.scala 52:49]
  wire  IST0_reset; // @[Triangle.scala 52:49]
  wire  IST0_io_enable_IST0; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_nodeid_leaf; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_rayid_leaf; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_hiT_in; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_v00_x; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_v00_y; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_v00_z; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_v00_w; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_v11_in_x; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_v11_in_y; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_v11_in_z; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_v11_in_w; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_v22_in_x; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_v22_in_y; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_v22_in_z; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_v22_in_w; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_ray_o_in_x; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_ray_o_in_y; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_ray_o_in_z; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_ray_d_in_x; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_ray_d_in_y; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_ray_d_in_z; // @[Triangle.scala 52:49]
  wire  IST0_io_RAY_AABB_1; // @[Triangle.scala 52:49]
  wire  IST0_io_RAY_AABB_2; // @[Triangle.scala 52:49]
  wire  IST0_io_break_in; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_Oz; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_invDz_div; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_nodeid_ist0_out; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_rayid_ist0_out; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_hiT_out; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_v11_out_x; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_v11_out_y; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_v11_out_z; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_v11_out_w; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_v22_out_x; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_v22_out_y; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_v22_out_z; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_v22_out_w; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_ray_o_out_x; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_ray_o_out_y; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_ray_o_out_z; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_ray_d_out_x; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_ray_d_out_y; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_ray_d_out_z; // @[Triangle.scala 52:49]
  wire  IST0_io_enable_SU_out; // @[Triangle.scala 52:49]
  wire  IST0_io_break_out; // @[Triangle.scala 52:49]
  wire  IST0_io_RAY_AABB_1_out; // @[Triangle.scala 52:49]
  wire  IST0_io_RAY_AABB_2_out; // @[Triangle.scala 52:49]
  wire  SU_clock; // @[Triangle.scala 53:50]
  wire  SU_reset; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_invDz_div; // @[Triangle.scala 53:50]
  wire  SU_io_valid_in; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_v11_x; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_v11_y; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_v11_z; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_v11_w; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_v22_x; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_v22_y; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_v22_z; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_v22_w; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_ray_in; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_Oz; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_ray_o_in_x; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_ray_o_in_y; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_ray_o_in_z; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_ray_d_in_x; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_ray_d_in_y; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_ray_d_in_z; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_node_id_in; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_hitT_in; // @[Triangle.scala 53:50]
  wire  SU_io_break_in; // @[Triangle.scala 53:50]
  wire  SU_io_RAY_AABB_1; // @[Triangle.scala 53:50]
  wire  SU_io_RAY_AABB_2; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_fdiv_out; // @[Triangle.scala 53:50]
  wire  SU_io_valid_out; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_v11_out_x; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_v11_out_y; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_v11_out_z; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_v11_out_w; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_v22_out_x; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_v22_out_y; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_v22_out_z; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_v22_out_w; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_ray_out; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_Oz_out; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_ray_o_out_x; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_ray_o_out_y; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_ray_o_out_z; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_ray_d_out_x; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_ray_d_out_y; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_ray_d_out_z; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_node_id_out; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_hitT_out; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_counter_fdiv; // @[Triangle.scala 53:50]
  wire  SU_io_break_out; // @[Triangle.scala 53:50]
  wire  SU_io_RAY_AABB_1_out; // @[Triangle.scala 53:50]
  wire  SU_io_RAY_AABB_2_out; // @[Triangle.scala 53:50]
  wire  IST1_clock; // @[Triangle.scala 54:49]
  wire  IST1_reset; // @[Triangle.scala 54:49]
  wire  IST1_io_enable_IST1; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_nodeid_leaf_1; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_rayid_leaf_1; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_hiT_in; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_Oz; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_invDz; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_v11_in_x; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_v11_in_y; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_v11_in_z; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_v11_in_w; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_v22_in_x; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_v22_in_y; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_v22_in_z; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_v22_in_w; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_ray_o_in_x; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_ray_o_in_y; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_ray_o_in_z; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_ray_d_in_x; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_ray_d_in_y; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_ray_d_in_z; // @[Triangle.scala 54:49]
  wire  IST1_io_break_in; // @[Triangle.scala 54:49]
  wire  IST1_io_RAY_AABB_1; // @[Triangle.scala 54:49]
  wire  IST1_io_RAY_AABB_2; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_nodeid_ist1_out; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_rayid_ist1_out; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_hiT_out; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_t; // @[Triangle.scala 54:49]
  wire  IST1_io_pop_1; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_v11_out_x; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_v11_out_y; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_v11_out_z; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_v11_out_w; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_v22_out_x; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_v22_out_y; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_v22_out_z; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_v22_out_w; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_ray_o_out_x; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_ray_o_out_y; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_ray_o_out_z; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_ray_d_out_x; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_ray_d_out_y; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_ray_d_out_z; // @[Triangle.scala 54:49]
  wire  IST1_io_enable_IST2; // @[Triangle.scala 54:49]
  wire  IST1_io_break_out; // @[Triangle.scala 54:49]
  wire  IST1_io_break_ist1; // @[Triangle.scala 54:49]
  wire  IST1_io_RAY_AABB_1_out; // @[Triangle.scala 54:49]
  wire  IST1_io_RAY_AABB_2_out; // @[Triangle.scala 54:49]
  wire  IST2_clock; // @[Triangle.scala 55:49]
  wire  IST2_reset; // @[Triangle.scala 55:49]
  wire  IST2_io_enable_IST2; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_nodeid_leaf_2; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_rayid_leaf_2; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_hiT_in; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_v11_in_x; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_v11_in_y; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_v11_in_z; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_v11_in_w; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_v22_in_x; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_v22_in_y; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_v22_in_z; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_v22_in_w; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_ray_o_in_x; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_ray_o_in_y; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_ray_o_in_z; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_ray_d_in_x; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_ray_d_in_y; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_ray_d_in_z; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_t; // @[Triangle.scala 55:49]
  wire  IST2_io_break_in; // @[Triangle.scala 55:49]
  wire  IST2_io_RAY_AABB_1; // @[Triangle.scala 55:49]
  wire  IST2_io_RAY_AABB_2; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_nodeid_ist2_out; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_rayid_ist2_out; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_hiT_out; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_u; // @[Triangle.scala 55:49]
  wire  IST2_io_pop_2; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_t_out; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_v22_out_x; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_v22_out_y; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_v22_out_z; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_v22_out_w; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_ray_o_out_x; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_ray_o_out_y; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_ray_o_out_z; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_ray_d_out_x; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_ray_d_out_y; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_ray_d_out_z; // @[Triangle.scala 55:49]
  wire  IST2_io_enable_IST3; // @[Triangle.scala 55:49]
  wire  IST2_io_break_ist2; // @[Triangle.scala 55:49]
  wire  IST2_io_break_out; // @[Triangle.scala 55:49]
  wire  IST2_io_RAY_AABB_1_out; // @[Triangle.scala 55:49]
  wire  IST2_io_RAY_AABB_2_out; // @[Triangle.scala 55:49]
  wire  IST3_clock; // @[Triangle.scala 56:49]
  wire  IST3_reset; // @[Triangle.scala 56:49]
  wire  IST3_io_enable_IST3; // @[Triangle.scala 56:49]
  wire [31:0] IST3_io_nodeid_leaf_3; // @[Triangle.scala 56:49]
  wire [31:0] IST3_io_rayid_leaf_3; // @[Triangle.scala 56:49]
  wire [31:0] IST3_io_hiT_in; // @[Triangle.scala 56:49]
  wire [31:0] IST3_io_t_in; // @[Triangle.scala 56:49]
  wire [31:0] IST3_io_v22_in_x; // @[Triangle.scala 56:49]
  wire [31:0] IST3_io_v22_in_y; // @[Triangle.scala 56:49]
  wire [31:0] IST3_io_v22_in_z; // @[Triangle.scala 56:49]
  wire [31:0] IST3_io_v22_in_w; // @[Triangle.scala 56:49]
  wire [31:0] IST3_io_ray_o_in_x; // @[Triangle.scala 56:49]
  wire [31:0] IST3_io_ray_o_in_y; // @[Triangle.scala 56:49]
  wire [31:0] IST3_io_ray_o_in_z; // @[Triangle.scala 56:49]
  wire [31:0] IST3_io_ray_d_in_x; // @[Triangle.scala 56:49]
  wire [31:0] IST3_io_ray_d_in_y; // @[Triangle.scala 56:49]
  wire [31:0] IST3_io_ray_d_in_z; // @[Triangle.scala 56:49]
  wire [31:0] IST3_io_u_in; // @[Triangle.scala 56:49]
  wire  IST3_io_break_in; // @[Triangle.scala 56:49]
  wire  IST3_io_RAY_AABB_1; // @[Triangle.scala 56:49]
  wire  IST3_io_RAY_AABB_2; // @[Triangle.scala 56:49]
  wire [31:0] IST3_io_nodeid_ist3_out; // @[Triangle.scala 56:49]
  wire [31:0] IST3_io_rayid_ist3_out; // @[Triangle.scala 56:49]
  wire [31:0] IST3_io_hiT_out; // @[Triangle.scala 56:49]
  wire  IST3_io_hitT_en; // @[Triangle.scala 56:49]
  wire  IST3_io_pop_3; // @[Triangle.scala 56:49]
  wire [31:0] IST3_io_hitIndex; // @[Triangle.scala 56:49]
  wire  IST3_io_hitIndex_en; // @[Triangle.scala 56:49]
  wire  IST3_io_break_out; // @[Triangle.scala 56:49]
  wire  IST3_io_RAY_AABB_1_out; // @[Triangle.scala 56:49]
  wire  IST3_io_RAY_AABB_2_out; // @[Triangle.scala 56:49]
  IST0 IST0 ( // @[Triangle.scala 52:49]
    .clock(IST0_clock),
    .reset(IST0_reset),
    .io_enable_IST0(IST0_io_enable_IST0),
    .io_nodeid_leaf(IST0_io_nodeid_leaf),
    .io_rayid_leaf(IST0_io_rayid_leaf),
    .io_hiT_in(IST0_io_hiT_in),
    .io_v00_x(IST0_io_v00_x),
    .io_v00_y(IST0_io_v00_y),
    .io_v00_z(IST0_io_v00_z),
    .io_v00_w(IST0_io_v00_w),
    .io_v11_in_x(IST0_io_v11_in_x),
    .io_v11_in_y(IST0_io_v11_in_y),
    .io_v11_in_z(IST0_io_v11_in_z),
    .io_v11_in_w(IST0_io_v11_in_w),
    .io_v22_in_x(IST0_io_v22_in_x),
    .io_v22_in_y(IST0_io_v22_in_y),
    .io_v22_in_z(IST0_io_v22_in_z),
    .io_v22_in_w(IST0_io_v22_in_w),
    .io_ray_o_in_x(IST0_io_ray_o_in_x),
    .io_ray_o_in_y(IST0_io_ray_o_in_y),
    .io_ray_o_in_z(IST0_io_ray_o_in_z),
    .io_ray_d_in_x(IST0_io_ray_d_in_x),
    .io_ray_d_in_y(IST0_io_ray_d_in_y),
    .io_ray_d_in_z(IST0_io_ray_d_in_z),
    .io_RAY_AABB_1(IST0_io_RAY_AABB_1),
    .io_RAY_AABB_2(IST0_io_RAY_AABB_2),
    .io_break_in(IST0_io_break_in),
    .io_Oz(IST0_io_Oz),
    .io_invDz_div(IST0_io_invDz_div),
    .io_nodeid_ist0_out(IST0_io_nodeid_ist0_out),
    .io_rayid_ist0_out(IST0_io_rayid_ist0_out),
    .io_hiT_out(IST0_io_hiT_out),
    .io_v11_out_x(IST0_io_v11_out_x),
    .io_v11_out_y(IST0_io_v11_out_y),
    .io_v11_out_z(IST0_io_v11_out_z),
    .io_v11_out_w(IST0_io_v11_out_w),
    .io_v22_out_x(IST0_io_v22_out_x),
    .io_v22_out_y(IST0_io_v22_out_y),
    .io_v22_out_z(IST0_io_v22_out_z),
    .io_v22_out_w(IST0_io_v22_out_w),
    .io_ray_o_out_x(IST0_io_ray_o_out_x),
    .io_ray_o_out_y(IST0_io_ray_o_out_y),
    .io_ray_o_out_z(IST0_io_ray_o_out_z),
    .io_ray_d_out_x(IST0_io_ray_d_out_x),
    .io_ray_d_out_y(IST0_io_ray_d_out_y),
    .io_ray_d_out_z(IST0_io_ray_d_out_z),
    .io_enable_SU_out(IST0_io_enable_SU_out),
    .io_break_out(IST0_io_break_out),
    .io_RAY_AABB_1_out(IST0_io_RAY_AABB_1_out),
    .io_RAY_AABB_2_out(IST0_io_RAY_AABB_2_out)
  );
  Schedule_unit SU ( // @[Triangle.scala 53:50]
    .clock(SU_clock),
    .reset(SU_reset),
    .io_invDz_div(SU_io_invDz_div),
    .io_valid_in(SU_io_valid_in),
    .io_v11_x(SU_io_v11_x),
    .io_v11_y(SU_io_v11_y),
    .io_v11_z(SU_io_v11_z),
    .io_v11_w(SU_io_v11_w),
    .io_v22_x(SU_io_v22_x),
    .io_v22_y(SU_io_v22_y),
    .io_v22_z(SU_io_v22_z),
    .io_v22_w(SU_io_v22_w),
    .io_ray_in(SU_io_ray_in),
    .io_Oz(SU_io_Oz),
    .io_ray_o_in_x(SU_io_ray_o_in_x),
    .io_ray_o_in_y(SU_io_ray_o_in_y),
    .io_ray_o_in_z(SU_io_ray_o_in_z),
    .io_ray_d_in_x(SU_io_ray_d_in_x),
    .io_ray_d_in_y(SU_io_ray_d_in_y),
    .io_ray_d_in_z(SU_io_ray_d_in_z),
    .io_node_id_in(SU_io_node_id_in),
    .io_hitT_in(SU_io_hitT_in),
    .io_break_in(SU_io_break_in),
    .io_RAY_AABB_1(SU_io_RAY_AABB_1),
    .io_RAY_AABB_2(SU_io_RAY_AABB_2),
    .io_fdiv_out(SU_io_fdiv_out),
    .io_valid_out(SU_io_valid_out),
    .io_v11_out_x(SU_io_v11_out_x),
    .io_v11_out_y(SU_io_v11_out_y),
    .io_v11_out_z(SU_io_v11_out_z),
    .io_v11_out_w(SU_io_v11_out_w),
    .io_v22_out_x(SU_io_v22_out_x),
    .io_v22_out_y(SU_io_v22_out_y),
    .io_v22_out_z(SU_io_v22_out_z),
    .io_v22_out_w(SU_io_v22_out_w),
    .io_ray_out(SU_io_ray_out),
    .io_Oz_out(SU_io_Oz_out),
    .io_ray_o_out_x(SU_io_ray_o_out_x),
    .io_ray_o_out_y(SU_io_ray_o_out_y),
    .io_ray_o_out_z(SU_io_ray_o_out_z),
    .io_ray_d_out_x(SU_io_ray_d_out_x),
    .io_ray_d_out_y(SU_io_ray_d_out_y),
    .io_ray_d_out_z(SU_io_ray_d_out_z),
    .io_node_id_out(SU_io_node_id_out),
    .io_hitT_out(SU_io_hitT_out),
    .io_counter_fdiv(SU_io_counter_fdiv),
    .io_break_out(SU_io_break_out),
    .io_RAY_AABB_1_out(SU_io_RAY_AABB_1_out),
    .io_RAY_AABB_2_out(SU_io_RAY_AABB_2_out)
  );
  IST1 IST1 ( // @[Triangle.scala 54:49]
    .clock(IST1_clock),
    .reset(IST1_reset),
    .io_enable_IST1(IST1_io_enable_IST1),
    .io_nodeid_leaf_1(IST1_io_nodeid_leaf_1),
    .io_rayid_leaf_1(IST1_io_rayid_leaf_1),
    .io_hiT_in(IST1_io_hiT_in),
    .io_Oz(IST1_io_Oz),
    .io_invDz(IST1_io_invDz),
    .io_v11_in_x(IST1_io_v11_in_x),
    .io_v11_in_y(IST1_io_v11_in_y),
    .io_v11_in_z(IST1_io_v11_in_z),
    .io_v11_in_w(IST1_io_v11_in_w),
    .io_v22_in_x(IST1_io_v22_in_x),
    .io_v22_in_y(IST1_io_v22_in_y),
    .io_v22_in_z(IST1_io_v22_in_z),
    .io_v22_in_w(IST1_io_v22_in_w),
    .io_ray_o_in_x(IST1_io_ray_o_in_x),
    .io_ray_o_in_y(IST1_io_ray_o_in_y),
    .io_ray_o_in_z(IST1_io_ray_o_in_z),
    .io_ray_d_in_x(IST1_io_ray_d_in_x),
    .io_ray_d_in_y(IST1_io_ray_d_in_y),
    .io_ray_d_in_z(IST1_io_ray_d_in_z),
    .io_break_in(IST1_io_break_in),
    .io_RAY_AABB_1(IST1_io_RAY_AABB_1),
    .io_RAY_AABB_2(IST1_io_RAY_AABB_2),
    .io_nodeid_ist1_out(IST1_io_nodeid_ist1_out),
    .io_rayid_ist1_out(IST1_io_rayid_ist1_out),
    .io_hiT_out(IST1_io_hiT_out),
    .io_t(IST1_io_t),
    .io_pop_1(IST1_io_pop_1),
    .io_v11_out_x(IST1_io_v11_out_x),
    .io_v11_out_y(IST1_io_v11_out_y),
    .io_v11_out_z(IST1_io_v11_out_z),
    .io_v11_out_w(IST1_io_v11_out_w),
    .io_v22_out_x(IST1_io_v22_out_x),
    .io_v22_out_y(IST1_io_v22_out_y),
    .io_v22_out_z(IST1_io_v22_out_z),
    .io_v22_out_w(IST1_io_v22_out_w),
    .io_ray_o_out_x(IST1_io_ray_o_out_x),
    .io_ray_o_out_y(IST1_io_ray_o_out_y),
    .io_ray_o_out_z(IST1_io_ray_o_out_z),
    .io_ray_d_out_x(IST1_io_ray_d_out_x),
    .io_ray_d_out_y(IST1_io_ray_d_out_y),
    .io_ray_d_out_z(IST1_io_ray_d_out_z),
    .io_enable_IST2(IST1_io_enable_IST2),
    .io_break_out(IST1_io_break_out),
    .io_break_ist1(IST1_io_break_ist1),
    .io_RAY_AABB_1_out(IST1_io_RAY_AABB_1_out),
    .io_RAY_AABB_2_out(IST1_io_RAY_AABB_2_out)
  );
  IST2 IST2 ( // @[Triangle.scala 55:49]
    .clock(IST2_clock),
    .reset(IST2_reset),
    .io_enable_IST2(IST2_io_enable_IST2),
    .io_nodeid_leaf_2(IST2_io_nodeid_leaf_2),
    .io_rayid_leaf_2(IST2_io_rayid_leaf_2),
    .io_hiT_in(IST2_io_hiT_in),
    .io_v11_in_x(IST2_io_v11_in_x),
    .io_v11_in_y(IST2_io_v11_in_y),
    .io_v11_in_z(IST2_io_v11_in_z),
    .io_v11_in_w(IST2_io_v11_in_w),
    .io_v22_in_x(IST2_io_v22_in_x),
    .io_v22_in_y(IST2_io_v22_in_y),
    .io_v22_in_z(IST2_io_v22_in_z),
    .io_v22_in_w(IST2_io_v22_in_w),
    .io_ray_o_in_x(IST2_io_ray_o_in_x),
    .io_ray_o_in_y(IST2_io_ray_o_in_y),
    .io_ray_o_in_z(IST2_io_ray_o_in_z),
    .io_ray_d_in_x(IST2_io_ray_d_in_x),
    .io_ray_d_in_y(IST2_io_ray_d_in_y),
    .io_ray_d_in_z(IST2_io_ray_d_in_z),
    .io_t(IST2_io_t),
    .io_break_in(IST2_io_break_in),
    .io_RAY_AABB_1(IST2_io_RAY_AABB_1),
    .io_RAY_AABB_2(IST2_io_RAY_AABB_2),
    .io_nodeid_ist2_out(IST2_io_nodeid_ist2_out),
    .io_rayid_ist2_out(IST2_io_rayid_ist2_out),
    .io_hiT_out(IST2_io_hiT_out),
    .io_u(IST2_io_u),
    .io_pop_2(IST2_io_pop_2),
    .io_t_out(IST2_io_t_out),
    .io_v22_out_x(IST2_io_v22_out_x),
    .io_v22_out_y(IST2_io_v22_out_y),
    .io_v22_out_z(IST2_io_v22_out_z),
    .io_v22_out_w(IST2_io_v22_out_w),
    .io_ray_o_out_x(IST2_io_ray_o_out_x),
    .io_ray_o_out_y(IST2_io_ray_o_out_y),
    .io_ray_o_out_z(IST2_io_ray_o_out_z),
    .io_ray_d_out_x(IST2_io_ray_d_out_x),
    .io_ray_d_out_y(IST2_io_ray_d_out_y),
    .io_ray_d_out_z(IST2_io_ray_d_out_z),
    .io_enable_IST3(IST2_io_enable_IST3),
    .io_break_ist2(IST2_io_break_ist2),
    .io_break_out(IST2_io_break_out),
    .io_RAY_AABB_1_out(IST2_io_RAY_AABB_1_out),
    .io_RAY_AABB_2_out(IST2_io_RAY_AABB_2_out)
  );
  IST3 IST3 ( // @[Triangle.scala 56:49]
    .clock(IST3_clock),
    .reset(IST3_reset),
    .io_enable_IST3(IST3_io_enable_IST3),
    .io_nodeid_leaf_3(IST3_io_nodeid_leaf_3),
    .io_rayid_leaf_3(IST3_io_rayid_leaf_3),
    .io_hiT_in(IST3_io_hiT_in),
    .io_t_in(IST3_io_t_in),
    .io_v22_in_x(IST3_io_v22_in_x),
    .io_v22_in_y(IST3_io_v22_in_y),
    .io_v22_in_z(IST3_io_v22_in_z),
    .io_v22_in_w(IST3_io_v22_in_w),
    .io_ray_o_in_x(IST3_io_ray_o_in_x),
    .io_ray_o_in_y(IST3_io_ray_o_in_y),
    .io_ray_o_in_z(IST3_io_ray_o_in_z),
    .io_ray_d_in_x(IST3_io_ray_d_in_x),
    .io_ray_d_in_y(IST3_io_ray_d_in_y),
    .io_ray_d_in_z(IST3_io_ray_d_in_z),
    .io_u_in(IST3_io_u_in),
    .io_break_in(IST3_io_break_in),
    .io_RAY_AABB_1(IST3_io_RAY_AABB_1),
    .io_RAY_AABB_2(IST3_io_RAY_AABB_2),
    .io_nodeid_ist3_out(IST3_io_nodeid_ist3_out),
    .io_rayid_ist3_out(IST3_io_rayid_ist3_out),
    .io_hiT_out(IST3_io_hiT_out),
    .io_hitT_en(IST3_io_hitT_en),
    .io_pop_3(IST3_io_pop_3),
    .io_hitIndex(IST3_io_hitIndex),
    .io_hitIndex_en(IST3_io_hitIndex_en),
    .io_break_out(IST3_io_break_out),
    .io_RAY_AABB_1_out(IST3_io_RAY_AABB_1_out),
    .io_RAY_AABB_2_out(IST3_io_RAY_AABB_2_out)
  );
  assign io_pop_1 = IST1_io_pop_1; // @[Triangle.scala 129:41]
  assign io_break_1 = IST1_io_break_out; // @[Triangle.scala 132:39]
  assign io_pop_2 = IST2_io_pop_2; // @[Triangle.scala 133:41]
  assign io_break_2 = IST2_io_break_out; // @[Triangle.scala 136:39]
  assign io_pop_3 = IST3_io_pop_3; // @[Triangle.scala 137:41]
  assign io_break_3 = IST3_io_break_out; // @[Triangle.scala 140:39]
  assign io_hiT_out_1 = IST1_io_hiT_out; // @[Triangle.scala 141:37]
  assign io_hiT_out_2 = IST2_io_hiT_out; // @[Triangle.scala 142:37]
  assign io_hiT_out_3 = IST3_io_hiT_out; // @[Triangle.scala 143:37]
  assign io_hitT_en = IST3_io_hitT_en; // @[Triangle.scala 144:40]
  assign io_hitIndex = IST3_io_hitIndex; // @[Triangle.scala 146:40]
  assign io_hitIndex_en = IST3_io_hitIndex_en; // @[Triangle.scala 145:35]
  assign io_node_id_out_1 = IST1_io_nodeid_ist1_out; // @[Triangle.scala 131:30]
  assign io_node_id_out_2 = IST2_io_nodeid_ist2_out; // @[Triangle.scala 135:30]
  assign io_node_id_out_3 = IST3_io_nodeid_ist3_out; // @[Triangle.scala 139:30]
  assign io_ray_id_ist1 = IST1_io_rayid_ist1_out; // @[Triangle.scala 130:37]
  assign io_ray_id_ist2 = IST2_io_rayid_ist2_out; // @[Triangle.scala 134:37]
  assign io_ray_id_ist3 = IST3_io_rayid_ist3_out; // @[Triangle.scala 138:37]
  assign io_counter_fdiv = {{32'd0}, SU_io_counter_fdiv}; // @[Triangle.scala 85:37]
  assign io_RAY_AABB_1_out_IST1 = IST1_io_RAY_AABB_1_out; // @[Triangle.scala 148:33]
  assign io_RAY_AABB_2_out_IST1 = IST1_io_RAY_AABB_2_out; // @[Triangle.scala 149:33]
  assign io_RAY_AABB_1_out_IST2 = IST2_io_RAY_AABB_1_out; // @[Triangle.scala 150:33]
  assign io_RAY_AABB_2_out_IST2 = IST2_io_RAY_AABB_2_out; // @[Triangle.scala 151:33]
  assign io_RAY_AABB_1_out_IST3 = IST3_io_RAY_AABB_1_out; // @[Triangle.scala 152:33]
  assign io_RAY_AABB_2_out_IST3 = IST3_io_RAY_AABB_2_out; // @[Triangle.scala 153:33]
  assign IST0_clock = clock;
  assign IST0_reset = reset;
  assign IST0_io_enable_IST0 = io_To_IST0_enable; // @[Triangle.scala 61:32]
  assign IST0_io_nodeid_leaf = io_nodeid_leaf; // @[Triangle.scala 62:33]
  assign IST0_io_rayid_leaf = io_rayid_leaf; // @[Triangle.scala 63:36]
  assign IST0_io_hiT_in = io_hiT_in; // @[Triangle.scala 64:40]
  assign IST0_io_v00_x = io_v00_in_x; // @[Triangle.scala 65:43]
  assign IST0_io_v00_y = io_v00_in_y; // @[Triangle.scala 65:43]
  assign IST0_io_v00_z = io_v00_in_z; // @[Triangle.scala 65:43]
  assign IST0_io_v00_w = io_v00_in_w; // @[Triangle.scala 65:43]
  assign IST0_io_v11_in_x = io_v11_in_x; // @[Triangle.scala 66:40]
  assign IST0_io_v11_in_y = io_v11_in_y; // @[Triangle.scala 66:40]
  assign IST0_io_v11_in_z = io_v11_in_z; // @[Triangle.scala 66:40]
  assign IST0_io_v11_in_w = io_v11_in_w; // @[Triangle.scala 66:40]
  assign IST0_io_v22_in_x = io_v22_in_x; // @[Triangle.scala 67:40]
  assign IST0_io_v22_in_y = io_v22_in_y; // @[Triangle.scala 67:40]
  assign IST0_io_v22_in_z = io_v22_in_z; // @[Triangle.scala 67:40]
  assign IST0_io_v22_in_w = io_v22_in_w; // @[Triangle.scala 67:40]
  assign IST0_io_ray_o_in_x = io_ray_o_in_x; // @[Triangle.scala 68:37]
  assign IST0_io_ray_o_in_y = io_ray_o_in_y; // @[Triangle.scala 68:37]
  assign IST0_io_ray_o_in_z = io_ray_o_in_z; // @[Triangle.scala 68:37]
  assign IST0_io_ray_d_in_x = io_ray_d_in_x; // @[Triangle.scala 69:37]
  assign IST0_io_ray_d_in_y = io_ray_d_in_y; // @[Triangle.scala 69:37]
  assign IST0_io_ray_d_in_z = io_ray_d_in_z; // @[Triangle.scala 69:37]
  assign IST0_io_RAY_AABB_1 = io_RAY_AABB_1; // @[Triangle.scala 59:31]
  assign IST0_io_RAY_AABB_2 = io_RAY_AABB_2; // @[Triangle.scala 60:31]
  assign IST0_io_break_in = io_break_in; // @[Triangle.scala 70:37]
  assign SU_clock = clock;
  assign SU_reset = reset;
  assign SU_io_invDz_div = IST0_io_invDz_div; // @[Triangle.scala 77:36]
  assign SU_io_valid_in = IST0_io_enable_SU_out; // @[Triangle.scala 75:39]
  assign SU_io_v11_x = IST0_io_v11_out_x; // @[Triangle.scala 81:43]
  assign SU_io_v11_y = IST0_io_v11_out_y; // @[Triangle.scala 81:43]
  assign SU_io_v11_z = IST0_io_v11_out_z; // @[Triangle.scala 81:43]
  assign SU_io_v11_w = IST0_io_v11_out_w; // @[Triangle.scala 81:43]
  assign SU_io_v22_x = IST0_io_v22_out_x; // @[Triangle.scala 82:43]
  assign SU_io_v22_y = IST0_io_v22_out_y; // @[Triangle.scala 82:43]
  assign SU_io_v22_z = IST0_io_v22_out_z; // @[Triangle.scala 82:43]
  assign SU_io_v22_w = IST0_io_v22_out_w; // @[Triangle.scala 82:43]
  assign SU_io_ray_in = IST0_io_rayid_ist0_out; // @[Triangle.scala 79:40]
  assign SU_io_Oz = IST0_io_Oz; // @[Triangle.scala 76:44]
  assign SU_io_ray_o_in_x = IST0_io_ray_o_out_x; // @[Triangle.scala 83:37]
  assign SU_io_ray_o_in_y = IST0_io_ray_o_out_y; // @[Triangle.scala 83:37]
  assign SU_io_ray_o_in_z = IST0_io_ray_o_out_z; // @[Triangle.scala 83:37]
  assign SU_io_ray_d_in_x = IST0_io_ray_d_out_x; // @[Triangle.scala 84:37]
  assign SU_io_ray_d_in_y = IST0_io_ray_d_out_y; // @[Triangle.scala 84:37]
  assign SU_io_ray_d_in_z = IST0_io_ray_d_out_z; // @[Triangle.scala 84:37]
  assign SU_io_node_id_in = IST0_io_nodeid_ist0_out; // @[Triangle.scala 78:33]
  assign SU_io_hitT_in = IST0_io_hiT_out; // @[Triangle.scala 80:39]
  assign SU_io_break_in = IST0_io_break_out; // @[Triangle.scala 74:37]
  assign SU_io_RAY_AABB_1 = IST0_io_RAY_AABB_1_out; // @[Triangle.scala 72:31]
  assign SU_io_RAY_AABB_2 = IST0_io_RAY_AABB_2_out; // @[Triangle.scala 73:31]
  assign IST1_clock = clock;
  assign IST1_reset = reset;
  assign IST1_io_enable_IST1 = SU_io_valid_out; // @[Triangle.scala 90:32]
  assign IST1_io_nodeid_leaf_1 = SU_io_node_id_out; // @[Triangle.scala 91:30]
  assign IST1_io_rayid_leaf_1 = SU_io_ray_out; // @[Triangle.scala 92:33]
  assign IST1_io_hiT_in = SU_io_hitT_out; // @[Triangle.scala 93:40]
  assign IST1_io_Oz = SU_io_Oz_out; // @[Triangle.scala 94:44]
  assign IST1_io_invDz = SU_io_fdiv_out; // @[Triangle.scala 95:41]
  assign IST1_io_v11_in_x = SU_io_v11_out_x; // @[Triangle.scala 96:40]
  assign IST1_io_v11_in_y = SU_io_v11_out_y; // @[Triangle.scala 96:40]
  assign IST1_io_v11_in_z = SU_io_v11_out_z; // @[Triangle.scala 96:40]
  assign IST1_io_v11_in_w = SU_io_v11_out_w; // @[Triangle.scala 96:40]
  assign IST1_io_v22_in_x = SU_io_v22_out_x; // @[Triangle.scala 97:40]
  assign IST1_io_v22_in_y = SU_io_v22_out_y; // @[Triangle.scala 97:40]
  assign IST1_io_v22_in_z = SU_io_v22_out_z; // @[Triangle.scala 97:40]
  assign IST1_io_v22_in_w = SU_io_v22_out_w; // @[Triangle.scala 97:40]
  assign IST1_io_ray_o_in_x = SU_io_ray_o_out_x; // @[Triangle.scala 98:37]
  assign IST1_io_ray_o_in_y = SU_io_ray_o_out_y; // @[Triangle.scala 98:37]
  assign IST1_io_ray_o_in_z = SU_io_ray_o_out_z; // @[Triangle.scala 98:37]
  assign IST1_io_ray_d_in_x = SU_io_ray_d_out_x; // @[Triangle.scala 99:37]
  assign IST1_io_ray_d_in_y = SU_io_ray_d_out_y; // @[Triangle.scala 99:37]
  assign IST1_io_ray_d_in_z = SU_io_ray_d_out_z; // @[Triangle.scala 99:37]
  assign IST1_io_break_in = SU_io_break_out; // @[Triangle.scala 89:36]
  assign IST1_io_RAY_AABB_1 = SU_io_RAY_AABB_1_out; // @[Triangle.scala 87:30]
  assign IST1_io_RAY_AABB_2 = SU_io_RAY_AABB_2_out; // @[Triangle.scala 88:30]
  assign IST2_clock = clock;
  assign IST2_reset = reset;
  assign IST2_io_enable_IST2 = IST1_io_enable_IST2; // @[Triangle.scala 105:35]
  assign IST2_io_nodeid_leaf_2 = IST1_io_nodeid_ist1_out; // @[Triangle.scala 106:33]
  assign IST2_io_rayid_leaf_2 = IST1_io_rayid_ist1_out; // @[Triangle.scala 107:36]
  assign IST2_io_hiT_in = IST1_io_hiT_out; // @[Triangle.scala 108:42]
  assign IST2_io_v11_in_x = IST1_io_v11_out_x; // @[Triangle.scala 109:42]
  assign IST2_io_v11_in_y = IST1_io_v11_out_y; // @[Triangle.scala 109:42]
  assign IST2_io_v11_in_z = IST1_io_v11_out_z; // @[Triangle.scala 109:42]
  assign IST2_io_v11_in_w = IST1_io_v11_out_w; // @[Triangle.scala 109:42]
  assign IST2_io_v22_in_x = IST1_io_v22_out_x; // @[Triangle.scala 110:42]
  assign IST2_io_v22_in_y = IST1_io_v22_out_y; // @[Triangle.scala 110:42]
  assign IST2_io_v22_in_z = IST1_io_v22_out_z; // @[Triangle.scala 110:42]
  assign IST2_io_v22_in_w = IST1_io_v22_out_w; // @[Triangle.scala 110:42]
  assign IST2_io_ray_o_in_x = IST1_io_ray_o_out_x; // @[Triangle.scala 111:40]
  assign IST2_io_ray_o_in_y = IST1_io_ray_o_out_y; // @[Triangle.scala 111:40]
  assign IST2_io_ray_o_in_z = IST1_io_ray_o_out_z; // @[Triangle.scala 111:40]
  assign IST2_io_ray_d_in_x = IST1_io_ray_d_out_x; // @[Triangle.scala 112:40]
  assign IST2_io_ray_d_in_y = IST1_io_ray_d_out_y; // @[Triangle.scala 112:40]
  assign IST2_io_ray_d_in_z = IST1_io_ray_d_out_z; // @[Triangle.scala 112:40]
  assign IST2_io_t = IST1_io_t; // @[Triangle.scala 113:49]
  assign IST2_io_break_in = IST1_io_break_ist1; // @[Triangle.scala 103:39]
  assign IST2_io_RAY_AABB_1 = IST1_io_RAY_AABB_1_out; // @[Triangle.scala 101:33]
  assign IST2_io_RAY_AABB_2 = IST1_io_RAY_AABB_2_out; // @[Triangle.scala 102:33]
  assign IST3_clock = clock;
  assign IST3_reset = reset;
  assign IST3_io_enable_IST3 = IST2_io_enable_IST3; // @[Triangle.scala 118:38]
  assign IST3_io_nodeid_leaf_3 = IST2_io_nodeid_ist2_out; // @[Triangle.scala 119:36]
  assign IST3_io_rayid_leaf_3 = IST2_io_rayid_ist2_out; // @[Triangle.scala 120:39]
  assign IST3_io_hiT_in = IST2_io_hiT_out; // @[Triangle.scala 121:45]
  assign IST3_io_t_in = IST2_io_t_out; // @[Triangle.scala 122:48]
  assign IST3_io_v22_in_x = IST2_io_v22_out_x; // @[Triangle.scala 123:45]
  assign IST3_io_v22_in_y = IST2_io_v22_out_y; // @[Triangle.scala 123:45]
  assign IST3_io_v22_in_z = IST2_io_v22_out_z; // @[Triangle.scala 123:45]
  assign IST3_io_v22_in_w = IST2_io_v22_out_w; // @[Triangle.scala 123:45]
  assign IST3_io_ray_o_in_x = IST2_io_ray_o_out_x; // @[Triangle.scala 124:41]
  assign IST3_io_ray_o_in_y = IST2_io_ray_o_out_y; // @[Triangle.scala 124:41]
  assign IST3_io_ray_o_in_z = IST2_io_ray_o_out_z; // @[Triangle.scala 124:41]
  assign IST3_io_ray_d_in_x = IST2_io_ray_d_out_x; // @[Triangle.scala 125:41]
  assign IST3_io_ray_d_in_y = IST2_io_ray_d_out_y; // @[Triangle.scala 125:41]
  assign IST3_io_ray_d_in_z = IST2_io_ray_d_out_z; // @[Triangle.scala 125:41]
  assign IST3_io_u_in = IST2_io_u; // @[Triangle.scala 126:47]
  assign IST3_io_break_in = IST2_io_break_ist2; // @[Triangle.scala 117:42]
  assign IST3_io_RAY_AABB_1 = IST2_io_RAY_AABB_1_out; // @[Triangle.scala 115:35]
  assign IST3_io_RAY_AABB_2 = IST2_io_RAY_AABB_2_out; // @[Triangle.scala 116:35]
endmodule
module TOP_AO(
  input         clock,
  input         reset,
  output [31:0] io_hitT,
  output [31:0] io_hitIndex,
  output        io_rtp_finish,
  output [31:0] io_ray_id_triangle,
  output [63:0] io_counter_fdiv,
  output [63:0] io_TRV_1_valid,
  output [63:0] io_TRV_2_valid,
  output [63:0] io_IST_1_valid,
  output [63:0] io_clock_count
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [63:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  wire  Ray_Dispatch_clock; // @[Top_AO.scala 24:44]
  wire  Ray_Dispatch_reset; // @[Top_AO.scala 24:44]
  wire  Ray_Dispatch_io_dispatch; // @[Top_AO.scala 24:44]
  wire  Ray_Dispatch_io_dispatch_2; // @[Top_AO.scala 24:44]
  wire [31:0] Ray_Dispatch_io_rayid_id; // @[Top_AO.scala 24:44]
  wire [31:0] Ray_Dispatch_io_rayid_id_2; // @[Top_AO.scala 24:44]
  wire  Ray_Dispatch_io_ray_out; // @[Top_AO.scala 24:44]
  wire  Ray_Dispatch_io_ray_out_2; // @[Top_AO.scala 24:44]
  wire  Ray_Dispatch_io_ray_finish; // @[Top_AO.scala 24:44]
  wire  Ray_origx_clock; // @[Top_AO.scala 25:48]
  wire [31:0] Ray_origx_io_Ray_id; // @[Top_AO.scala 25:48]
  wire [31:0] Ray_origx_io_Ray_id_2; // @[Top_AO.scala 25:48]
  wire [31:0] Ray_origx_io_Ray_out; // @[Top_AO.scala 25:48]
  wire [31:0] Ray_origx_io_Ray_out_2; // @[Top_AO.scala 25:48]
  wire  Ray_origy_clock; // @[Top_AO.scala 26:48]
  wire [31:0] Ray_origy_io_Ray_id; // @[Top_AO.scala 26:48]
  wire [31:0] Ray_origy_io_Ray_id_2; // @[Top_AO.scala 26:48]
  wire [31:0] Ray_origy_io_Ray_out; // @[Top_AO.scala 26:48]
  wire [31:0] Ray_origy_io_Ray_out_2; // @[Top_AO.scala 26:48]
  wire  Ray_origz_clock; // @[Top_AO.scala 27:48]
  wire [31:0] Ray_origz_io_Ray_id; // @[Top_AO.scala 27:48]
  wire [31:0] Ray_origz_io_Ray_id_2; // @[Top_AO.scala 27:48]
  wire [31:0] Ray_origz_io_Ray_out; // @[Top_AO.scala 27:48]
  wire [31:0] Ray_origz_io_Ray_out_2; // @[Top_AO.scala 27:48]
  wire  Ray_dirx_clock; // @[Top_AO.scala 30:50]
  wire [31:0] Ray_dirx_io_Ray_id; // @[Top_AO.scala 30:50]
  wire [31:0] Ray_dirx_io_Ray_id_2; // @[Top_AO.scala 30:50]
  wire [31:0] Ray_dirx_io_Ray_out; // @[Top_AO.scala 30:50]
  wire [31:0] Ray_dirx_io_Ray_out_2; // @[Top_AO.scala 30:50]
  wire  Ray_diry_clock; // @[Top_AO.scala 31:49]
  wire [31:0] Ray_diry_io_Ray_id; // @[Top_AO.scala 31:49]
  wire [31:0] Ray_diry_io_Ray_id_2; // @[Top_AO.scala 31:49]
  wire [31:0] Ray_diry_io_Ray_out; // @[Top_AO.scala 31:49]
  wire [31:0] Ray_diry_io_Ray_out_2; // @[Top_AO.scala 31:49]
  wire  Ray_dirz_clock; // @[Top_AO.scala 32:49]
  wire [31:0] Ray_dirz_io_Ray_id; // @[Top_AO.scala 32:49]
  wire [31:0] Ray_dirz_io_Ray_id_2; // @[Top_AO.scala 32:49]
  wire [31:0] Ray_dirz_io_Ray_out; // @[Top_AO.scala 32:49]
  wire [31:0] Ray_dirz_io_Ray_out_2; // @[Top_AO.scala 32:49]
  wire  Ray_hitT_clock; // @[Top_AO.scala 33:49]
  wire [31:0] Ray_hitT_io_Ray_id; // @[Top_AO.scala 33:49]
  wire [31:0] Ray_hitT_io_Ray_id_2; // @[Top_AO.scala 33:49]
  wire [31:0] Ray_hitT_io_Ray_out; // @[Top_AO.scala 33:49]
  wire [31:0] Ray_hitT_io_Ray_out_2; // @[Top_AO.scala 33:49]
  wire  Ray_idirx_clock; // @[Top_AO.scala 35:49]
  wire [31:0] Ray_idirx_io_Ray_id; // @[Top_AO.scala 35:49]
  wire [31:0] Ray_idirx_io_Ray_id_2; // @[Top_AO.scala 35:49]
  wire [31:0] Ray_idirx_io_Ray_out; // @[Top_AO.scala 35:49]
  wire [31:0] Ray_idirx_io_Ray_out_2; // @[Top_AO.scala 35:49]
  wire  Ray_idiry_clock; // @[Top_AO.scala 36:49]
  wire [31:0] Ray_idiry_io_Ray_id; // @[Top_AO.scala 36:49]
  wire [31:0] Ray_idiry_io_Ray_id_2; // @[Top_AO.scala 36:49]
  wire [31:0] Ray_idiry_io_Ray_out; // @[Top_AO.scala 36:49]
  wire [31:0] Ray_idiry_io_Ray_out_2; // @[Top_AO.scala 36:49]
  wire  Ray_idirz_clock; // @[Top_AO.scala 37:49]
  wire [31:0] Ray_idirz_io_Ray_id; // @[Top_AO.scala 37:49]
  wire [31:0] Ray_idirz_io_Ray_id_2; // @[Top_AO.scala 37:49]
  wire [31:0] Ray_idirz_io_Ray_out; // @[Top_AO.scala 37:49]
  wire [31:0] Ray_idirz_io_Ray_out_2; // @[Top_AO.scala 37:49]
  wire  Ray_oodx_clock; // @[Top_AO.scala 39:48]
  wire [31:0] Ray_oodx_io_Ray_id; // @[Top_AO.scala 39:48]
  wire [31:0] Ray_oodx_io_Ray_id_2; // @[Top_AO.scala 39:48]
  wire [31:0] Ray_oodx_io_Ray_out; // @[Top_AO.scala 39:48]
  wire [31:0] Ray_oodx_io_Ray_out_2; // @[Top_AO.scala 39:48]
  wire  Ray_oody_clock; // @[Top_AO.scala 40:48]
  wire [31:0] Ray_oody_io_Ray_id; // @[Top_AO.scala 40:48]
  wire [31:0] Ray_oody_io_Ray_id_2; // @[Top_AO.scala 40:48]
  wire [31:0] Ray_oody_io_Ray_out; // @[Top_AO.scala 40:48]
  wire [31:0] Ray_oody_io_Ray_out_2; // @[Top_AO.scala 40:48]
  wire  Ray_oodz_clock; // @[Top_AO.scala 41:48]
  wire [31:0] Ray_oodz_io_Ray_id; // @[Top_AO.scala 41:48]
  wire [31:0] Ray_oodz_io_Ray_id_2; // @[Top_AO.scala 41:48]
  wire [31:0] Ray_oodz_io_Ray_out; // @[Top_AO.scala 41:48]
  wire [31:0] Ray_oodz_io_Ray_out_2; // @[Top_AO.scala 41:48]
  wire  BVH_RAM_0_x_clock; // @[Top_AO.scala 43:41]
  wire [31:0] BVH_RAM_0_x_io_BVH_id; // @[Top_AO.scala 43:41]
  wire [31:0] BVH_RAM_0_x_io_BVH_id_2; // @[Top_AO.scala 43:41]
  wire [31:0] BVH_RAM_0_x_io_BVH_out; // @[Top_AO.scala 43:41]
  wire [31:0] BVH_RAM_0_x_io_BVH_out_2; // @[Top_AO.scala 43:41]
  wire  BVH_RAM_0_y_clock; // @[Top_AO.scala 44:41]
  wire [31:0] BVH_RAM_0_y_io_BVH_id; // @[Top_AO.scala 44:41]
  wire [31:0] BVH_RAM_0_y_io_BVH_id_2; // @[Top_AO.scala 44:41]
  wire [31:0] BVH_RAM_0_y_io_BVH_out; // @[Top_AO.scala 44:41]
  wire [31:0] BVH_RAM_0_y_io_BVH_out_2; // @[Top_AO.scala 44:41]
  wire  BVH_RAM_0_z_clock; // @[Top_AO.scala 45:41]
  wire [31:0] BVH_RAM_0_z_io_BVH_id; // @[Top_AO.scala 45:41]
  wire [31:0] BVH_RAM_0_z_io_BVH_id_2; // @[Top_AO.scala 45:41]
  wire [31:0] BVH_RAM_0_z_io_BVH_out; // @[Top_AO.scala 45:41]
  wire [31:0] BVH_RAM_0_z_io_BVH_out_2; // @[Top_AO.scala 45:41]
  wire  BVH_RAM_0_w_clock; // @[Top_AO.scala 46:40]
  wire [31:0] BVH_RAM_0_w_io_BVH_id; // @[Top_AO.scala 46:40]
  wire [31:0] BVH_RAM_0_w_io_BVH_id_2; // @[Top_AO.scala 46:40]
  wire [31:0] BVH_RAM_0_w_io_BVH_out; // @[Top_AO.scala 46:40]
  wire [31:0] BVH_RAM_0_w_io_BVH_out_2; // @[Top_AO.scala 46:40]
  wire  BVH_RAM_1_x_clock; // @[Top_AO.scala 48:41]
  wire [31:0] BVH_RAM_1_x_io_BVH_id; // @[Top_AO.scala 48:41]
  wire [31:0] BVH_RAM_1_x_io_BVH_id_2; // @[Top_AO.scala 48:41]
  wire [31:0] BVH_RAM_1_x_io_BVH_out; // @[Top_AO.scala 48:41]
  wire [31:0] BVH_RAM_1_x_io_BVH_out_2; // @[Top_AO.scala 48:41]
  wire  BVH_RAM_1_y_clock; // @[Top_AO.scala 49:41]
  wire [31:0] BVH_RAM_1_y_io_BVH_id; // @[Top_AO.scala 49:41]
  wire [31:0] BVH_RAM_1_y_io_BVH_id_2; // @[Top_AO.scala 49:41]
  wire [31:0] BVH_RAM_1_y_io_BVH_out; // @[Top_AO.scala 49:41]
  wire [31:0] BVH_RAM_1_y_io_BVH_out_2; // @[Top_AO.scala 49:41]
  wire  BVH_RAM_1_z_clock; // @[Top_AO.scala 50:41]
  wire [31:0] BVH_RAM_1_z_io_BVH_id; // @[Top_AO.scala 50:41]
  wire [31:0] BVH_RAM_1_z_io_BVH_id_2; // @[Top_AO.scala 50:41]
  wire [31:0] BVH_RAM_1_z_io_BVH_out; // @[Top_AO.scala 50:41]
  wire [31:0] BVH_RAM_1_z_io_BVH_out_2; // @[Top_AO.scala 50:41]
  wire  BVH_RAM_1_w_clock; // @[Top_AO.scala 51:40]
  wire [31:0] BVH_RAM_1_w_io_BVH_id; // @[Top_AO.scala 51:40]
  wire [31:0] BVH_RAM_1_w_io_BVH_id_2; // @[Top_AO.scala 51:40]
  wire [31:0] BVH_RAM_1_w_io_BVH_out; // @[Top_AO.scala 51:40]
  wire [31:0] BVH_RAM_1_w_io_BVH_out_2; // @[Top_AO.scala 51:40]
  wire  BVH_RAM_z_x_clock; // @[Top_AO.scala 53:41]
  wire [31:0] BVH_RAM_z_x_io_BVH_id; // @[Top_AO.scala 53:41]
  wire [31:0] BVH_RAM_z_x_io_BVH_id_2; // @[Top_AO.scala 53:41]
  wire [31:0] BVH_RAM_z_x_io_BVH_out; // @[Top_AO.scala 53:41]
  wire [31:0] BVH_RAM_z_x_io_BVH_out_2; // @[Top_AO.scala 53:41]
  wire  BVH_RAM_z_y_clock; // @[Top_AO.scala 54:41]
  wire [31:0] BVH_RAM_z_y_io_BVH_id; // @[Top_AO.scala 54:41]
  wire [31:0] BVH_RAM_z_y_io_BVH_id_2; // @[Top_AO.scala 54:41]
  wire [31:0] BVH_RAM_z_y_io_BVH_out; // @[Top_AO.scala 54:41]
  wire [31:0] BVH_RAM_z_y_io_BVH_out_2; // @[Top_AO.scala 54:41]
  wire  BVH_RAM_z_z_clock; // @[Top_AO.scala 55:41]
  wire [31:0] BVH_RAM_z_z_io_BVH_id; // @[Top_AO.scala 55:41]
  wire [31:0] BVH_RAM_z_z_io_BVH_id_2; // @[Top_AO.scala 55:41]
  wire [31:0] BVH_RAM_z_z_io_BVH_out; // @[Top_AO.scala 55:41]
  wire [31:0] BVH_RAM_z_z_io_BVH_out_2; // @[Top_AO.scala 55:41]
  wire  BVH_RAM_z_w_clock; // @[Top_AO.scala 56:40]
  wire [31:0] BVH_RAM_z_w_io_BVH_id; // @[Top_AO.scala 56:40]
  wire [31:0] BVH_RAM_z_w_io_BVH_id_2; // @[Top_AO.scala 56:40]
  wire [31:0] BVH_RAM_z_w_io_BVH_out; // @[Top_AO.scala 56:40]
  wire [31:0] BVH_RAM_z_w_io_BVH_out_2; // @[Top_AO.scala 56:40]
  wire  BVH_RAM_tmp_x_clock; // @[Top_AO.scala 58:37]
  wire [31:0] BVH_RAM_tmp_x_io_BVH_id; // @[Top_AO.scala 58:37]
  wire [31:0] BVH_RAM_tmp_x_io_BVH_id_2; // @[Top_AO.scala 58:37]
  wire [31:0] BVH_RAM_tmp_x_io_BVH_out; // @[Top_AO.scala 58:37]
  wire [31:0] BVH_RAM_tmp_x_io_BVH_out_2; // @[Top_AO.scala 58:37]
  wire  BVH_RAM_tmp_y_clock; // @[Top_AO.scala 59:37]
  wire [31:0] BVH_RAM_tmp_y_io_BVH_id; // @[Top_AO.scala 59:37]
  wire [31:0] BVH_RAM_tmp_y_io_BVH_id_2; // @[Top_AO.scala 59:37]
  wire [31:0] BVH_RAM_tmp_y_io_BVH_out; // @[Top_AO.scala 59:37]
  wire [31:0] BVH_RAM_tmp_y_io_BVH_out_2; // @[Top_AO.scala 59:37]
  wire  TRI_RAM_x_clock; // @[Top_AO.scala 61:50]
  wire [31:0] TRI_RAM_x_io_Triangle_id; // @[Top_AO.scala 61:50]
  wire [31:0] TRI_RAM_x_io_v00_out; // @[Top_AO.scala 61:50]
  wire [31:0] TRI_RAM_x_io_v11_out; // @[Top_AO.scala 61:50]
  wire [31:0] TRI_RAM_x_io_v22_out; // @[Top_AO.scala 61:50]
  wire [31:0] TRI_RAM_x_io_valid; // @[Top_AO.scala 61:50]
  wire  TRI_RAM_y_clock; // @[Top_AO.scala 62:50]
  wire [31:0] TRI_RAM_y_io_Triangle_id; // @[Top_AO.scala 62:50]
  wire [31:0] TRI_RAM_y_io_v00_out; // @[Top_AO.scala 62:50]
  wire [31:0] TRI_RAM_y_io_v11_out; // @[Top_AO.scala 62:50]
  wire [31:0] TRI_RAM_y_io_v22_out; // @[Top_AO.scala 62:50]
  wire  TRI_RAM_z_clock; // @[Top_AO.scala 63:50]
  wire [31:0] TRI_RAM_z_io_Triangle_id; // @[Top_AO.scala 63:50]
  wire [31:0] TRI_RAM_z_io_v00_out; // @[Top_AO.scala 63:50]
  wire [31:0] TRI_RAM_z_io_v11_out; // @[Top_AO.scala 63:50]
  wire [31:0] TRI_RAM_z_io_v22_out; // @[Top_AO.scala 63:50]
  wire  TRI_RAM_w_clock; // @[Top_AO.scala 64:49]
  wire [31:0] TRI_RAM_w_io_Triangle_id; // @[Top_AO.scala 64:49]
  wire [31:0] TRI_RAM_w_io_v00_out; // @[Top_AO.scala 64:49]
  wire [31:0] TRI_RAM_w_io_v11_out; // @[Top_AO.scala 64:49]
  wire [31:0] TRI_RAM_w_io_v22_out; // @[Top_AO.scala 64:49]
  wire  RAY_AABB_clock; // @[Top_AO.scala 65:46]
  wire  RAY_AABB_reset; // @[Top_AO.scala 65:46]
  wire [31:0] RAY_AABB_io_ray_idir_x; // @[Top_AO.scala 65:46]
  wire [31:0] RAY_AABB_io_ray_idir_y; // @[Top_AO.scala 65:46]
  wire [31:0] RAY_AABB_io_ray_idir_z; // @[Top_AO.scala 65:46]
  wire [31:0] RAY_AABB_io_ray_ood_x; // @[Top_AO.scala 65:46]
  wire [31:0] RAY_AABB_io_ray_ood_y; // @[Top_AO.scala 65:46]
  wire [31:0] RAY_AABB_io_ray_ood_z; // @[Top_AO.scala 65:46]
  wire [31:0] RAY_AABB_io_ray_hitT; // @[Top_AO.scala 65:46]
  wire [31:0] RAY_AABB_io_bvh_n0xy_x; // @[Top_AO.scala 65:46]
  wire [31:0] RAY_AABB_io_bvh_n0xy_y; // @[Top_AO.scala 65:46]
  wire [31:0] RAY_AABB_io_bvh_n0xy_z; // @[Top_AO.scala 65:46]
  wire [31:0] RAY_AABB_io_bvh_n0xy_w; // @[Top_AO.scala 65:46]
  wire [31:0] RAY_AABB_io_bvh_n1xy_x; // @[Top_AO.scala 65:46]
  wire [31:0] RAY_AABB_io_bvh_n1xy_y; // @[Top_AO.scala 65:46]
  wire [31:0] RAY_AABB_io_bvh_n1xy_z; // @[Top_AO.scala 65:46]
  wire [31:0] RAY_AABB_io_bvh_n1xy_w; // @[Top_AO.scala 65:46]
  wire [31:0] RAY_AABB_io_bvh_nz_x; // @[Top_AO.scala 65:46]
  wire [31:0] RAY_AABB_io_bvh_nz_y; // @[Top_AO.scala 65:46]
  wire [31:0] RAY_AABB_io_bvh_nz_z; // @[Top_AO.scala 65:46]
  wire [31:0] RAY_AABB_io_bvh_nz_w; // @[Top_AO.scala 65:46]
  wire [31:0] RAY_AABB_io_bvh_temp_x; // @[Top_AO.scala 65:46]
  wire [31:0] RAY_AABB_io_bvh_temp_y; // @[Top_AO.scala 65:46]
  wire [31:0] RAY_AABB_io_rayid; // @[Top_AO.scala 65:46]
  wire  RAY_AABB_io_valid_en; // @[Top_AO.scala 65:46]
  wire [31:0] RAY_AABB_io_rayid_out; // @[Top_AO.scala 65:46]
  wire [31:0] RAY_AABB_io_nodeIdx_0; // @[Top_AO.scala 65:46]
  wire [31:0] RAY_AABB_io_nodeIdx_1; // @[Top_AO.scala 65:46]
  wire [31:0] RAY_AABB_io_nodeIdx_2; // @[Top_AO.scala 65:46]
  wire  RAY_AABB_io_push; // @[Top_AO.scala 65:46]
  wire  RAY_AABB_io_pop; // @[Top_AO.scala 65:46]
  wire  RAY_AABB_io_leaf; // @[Top_AO.scala 65:46]
  wire  RAY_AABB_io_back; // @[Top_AO.scala 65:46]
  wire [31:0] RAY_AABB_io_hitT_out; // @[Top_AO.scala 65:46]
  wire  RAY_AABB_io_valid_out; // @[Top_AO.scala 65:46]
  wire  RAY_AABB_2_clock; // @[Top_AO.scala 66:48]
  wire  RAY_AABB_2_reset; // @[Top_AO.scala 66:48]
  wire [31:0] RAY_AABB_2_io_ray_idir_x; // @[Top_AO.scala 66:48]
  wire [31:0] RAY_AABB_2_io_ray_idir_y; // @[Top_AO.scala 66:48]
  wire [31:0] RAY_AABB_2_io_ray_idir_z; // @[Top_AO.scala 66:48]
  wire [31:0] RAY_AABB_2_io_ray_ood_x; // @[Top_AO.scala 66:48]
  wire [31:0] RAY_AABB_2_io_ray_ood_y; // @[Top_AO.scala 66:48]
  wire [31:0] RAY_AABB_2_io_ray_ood_z; // @[Top_AO.scala 66:48]
  wire [31:0] RAY_AABB_2_io_ray_hitT; // @[Top_AO.scala 66:48]
  wire [31:0] RAY_AABB_2_io_bvh_n0xy_x; // @[Top_AO.scala 66:48]
  wire [31:0] RAY_AABB_2_io_bvh_n0xy_y; // @[Top_AO.scala 66:48]
  wire [31:0] RAY_AABB_2_io_bvh_n0xy_z; // @[Top_AO.scala 66:48]
  wire [31:0] RAY_AABB_2_io_bvh_n0xy_w; // @[Top_AO.scala 66:48]
  wire [31:0] RAY_AABB_2_io_bvh_n1xy_x; // @[Top_AO.scala 66:48]
  wire [31:0] RAY_AABB_2_io_bvh_n1xy_y; // @[Top_AO.scala 66:48]
  wire [31:0] RAY_AABB_2_io_bvh_n1xy_z; // @[Top_AO.scala 66:48]
  wire [31:0] RAY_AABB_2_io_bvh_n1xy_w; // @[Top_AO.scala 66:48]
  wire [31:0] RAY_AABB_2_io_bvh_nz_x; // @[Top_AO.scala 66:48]
  wire [31:0] RAY_AABB_2_io_bvh_nz_y; // @[Top_AO.scala 66:48]
  wire [31:0] RAY_AABB_2_io_bvh_nz_z; // @[Top_AO.scala 66:48]
  wire [31:0] RAY_AABB_2_io_bvh_nz_w; // @[Top_AO.scala 66:48]
  wire [31:0] RAY_AABB_2_io_bvh_temp_x; // @[Top_AO.scala 66:48]
  wire [31:0] RAY_AABB_2_io_bvh_temp_y; // @[Top_AO.scala 66:48]
  wire [31:0] RAY_AABB_2_io_rayid; // @[Top_AO.scala 66:48]
  wire  RAY_AABB_2_io_valid_en; // @[Top_AO.scala 66:48]
  wire [31:0] RAY_AABB_2_io_rayid_out; // @[Top_AO.scala 66:48]
  wire [31:0] RAY_AABB_2_io_nodeIdx_0; // @[Top_AO.scala 66:48]
  wire [31:0] RAY_AABB_2_io_nodeIdx_1; // @[Top_AO.scala 66:48]
  wire [31:0] RAY_AABB_2_io_nodeIdx_2; // @[Top_AO.scala 66:48]
  wire  RAY_AABB_2_io_push; // @[Top_AO.scala 66:48]
  wire  RAY_AABB_2_io_pop; // @[Top_AO.scala 66:48]
  wire  RAY_AABB_2_io_leaf; // @[Top_AO.scala 66:48]
  wire  RAY_AABB_2_io_back; // @[Top_AO.scala 66:48]
  wire [31:0] RAY_AABB_2_io_hitT_out; // @[Top_AO.scala 66:48]
  wire  RAY_AABB_2_io_valid_out; // @[Top_AO.scala 66:48]
  wire  Arbitration_1_clock; // @[Top_AO.scala 67:50]
  wire  Arbitration_1_reset; // @[Top_AO.scala 67:50]
  wire [31:0] Arbitration_1_io_node_id_0; // @[Top_AO.scala 67:50]
  wire [63:0] Arbitration_1_io_ray_id_0; // @[Top_AO.scala 67:50]
  wire [31:0] Arbitration_1_io_hit_0; // @[Top_AO.scala 67:50]
  wire  Arbitration_1_io_valid_0; // @[Top_AO.scala 67:50]
  wire [31:0] Arbitration_1_io_node_id_1; // @[Top_AO.scala 67:50]
  wire [31:0] Arbitration_1_io_ray_id_1; // @[Top_AO.scala 67:50]
  wire  Arbitration_1_io_valid_1; // @[Top_AO.scala 67:50]
  wire [31:0] Arbitration_1_io_ray_id_2; // @[Top_AO.scala 67:50]
  wire  Arbitration_1_io_valid_2; // @[Top_AO.scala 67:50]
  wire [31:0] Arbitration_1_io_node_id_out; // @[Top_AO.scala 67:50]
  wire [31:0] Arbitration_1_io_ray_id_out; // @[Top_AO.scala 67:50]
  wire [31:0] Arbitration_1_io_hit_out; // @[Top_AO.scala 67:50]
  wire  Arbitration_1_io_valid_out; // @[Top_AO.scala 67:50]
  wire  Arbitration_1_2_clock; // @[Top_AO.scala 68:47]
  wire  Arbitration_1_2_reset; // @[Top_AO.scala 68:47]
  wire [31:0] Arbitration_1_2_io_node_id_0; // @[Top_AO.scala 68:47]
  wire [63:0] Arbitration_1_2_io_ray_id_0; // @[Top_AO.scala 68:47]
  wire [31:0] Arbitration_1_2_io_hit_0; // @[Top_AO.scala 68:47]
  wire  Arbitration_1_2_io_valid_0; // @[Top_AO.scala 68:47]
  wire [31:0] Arbitration_1_2_io_node_id_1; // @[Top_AO.scala 68:47]
  wire [31:0] Arbitration_1_2_io_ray_id_1; // @[Top_AO.scala 68:47]
  wire  Arbitration_1_2_io_valid_1; // @[Top_AO.scala 68:47]
  wire [31:0] Arbitration_1_2_io_ray_id_2; // @[Top_AO.scala 68:47]
  wire  Arbitration_1_2_io_valid_2; // @[Top_AO.scala 68:47]
  wire [31:0] Arbitration_1_2_io_node_id_out; // @[Top_AO.scala 68:47]
  wire [31:0] Arbitration_1_2_io_ray_id_out; // @[Top_AO.scala 68:47]
  wire [31:0] Arbitration_1_2_io_hit_out; // @[Top_AO.scala 68:47]
  wire  Arbitration_1_2_io_valid_out; // @[Top_AO.scala 68:47]
  wire  Arbitration_2_clock; // @[Top_AO.scala 70:45]
  wire  Arbitration_2_reset; // @[Top_AO.scala 70:45]
  wire [31:0] Arbitration_2_io_ray_id_2_0; // @[Top_AO.scala 70:45]
  wire [31:0] Arbitration_2_io_hit_2_0; // @[Top_AO.scala 70:45]
  wire  Arbitration_2_io_valid_2_0; // @[Top_AO.scala 70:45]
  wire [31:0] Arbitration_2_io_ray_id_2_1; // @[Top_AO.scala 70:45]
  wire [31:0] Arbitration_2_io_hit_2_1; // @[Top_AO.scala 70:45]
  wire  Arbitration_2_io_valid_2_1; // @[Top_AO.scala 70:45]
  wire [31:0] Arbitration_2_io_ray_id_2_2; // @[Top_AO.scala 70:45]
  wire [31:0] Arbitration_2_io_hit_2_2; // @[Top_AO.scala 70:45]
  wire  Arbitration_2_io_valid_2_2; // @[Top_AO.scala 70:45]
  wire [31:0] Arbitration_2_io_ray_id_2_3; // @[Top_AO.scala 70:45]
  wire [31:0] Arbitration_2_io_hit_2_3; // @[Top_AO.scala 70:45]
  wire  Arbitration_2_io_valid_2_3; // @[Top_AO.scala 70:45]
  wire [31:0] Arbitration_2_io_ray_id_out; // @[Top_AO.scala 70:45]
  wire [31:0] Arbitration_2_io_hit_out; // @[Top_AO.scala 70:45]
  wire  Arbitration_2_io_valid_out; // @[Top_AO.scala 70:45]
  wire  Arbitration_2_2_clock; // @[Top_AO.scala 71:42]
  wire  Arbitration_2_2_reset; // @[Top_AO.scala 71:42]
  wire [31:0] Arbitration_2_2_io_ray_id_2_0; // @[Top_AO.scala 71:42]
  wire [31:0] Arbitration_2_2_io_hit_2_0; // @[Top_AO.scala 71:42]
  wire  Arbitration_2_2_io_valid_2_0; // @[Top_AO.scala 71:42]
  wire [31:0] Arbitration_2_2_io_ray_id_2_1; // @[Top_AO.scala 71:42]
  wire [31:0] Arbitration_2_2_io_hit_2_1; // @[Top_AO.scala 71:42]
  wire  Arbitration_2_2_io_valid_2_1; // @[Top_AO.scala 71:42]
  wire [31:0] Arbitration_2_2_io_ray_id_2_2; // @[Top_AO.scala 71:42]
  wire [31:0] Arbitration_2_2_io_hit_2_2; // @[Top_AO.scala 71:42]
  wire  Arbitration_2_2_io_valid_2_2; // @[Top_AO.scala 71:42]
  wire [31:0] Arbitration_2_2_io_ray_id_2_3; // @[Top_AO.scala 71:42]
  wire [31:0] Arbitration_2_2_io_hit_2_3; // @[Top_AO.scala 71:42]
  wire  Arbitration_2_2_io_valid_2_3; // @[Top_AO.scala 71:42]
  wire [31:0] Arbitration_2_2_io_ray_id_out; // @[Top_AO.scala 71:42]
  wire [31:0] Arbitration_2_2_io_hit_out; // @[Top_AO.scala 71:42]
  wire  Arbitration_2_2_io_valid_out; // @[Top_AO.scala 71:42]
  wire  Arbitration_3_clock; // @[Top_AO.scala 72:45]
  wire  Arbitration_3_reset; // @[Top_AO.scala 72:45]
  wire [31:0] Arbitration_3_io_node_id_3_0; // @[Top_AO.scala 72:45]
  wire [31:0] Arbitration_3_io_ray_id_3_0; // @[Top_AO.scala 72:45]
  wire [31:0] Arbitration_3_io_hit_3_0; // @[Top_AO.scala 72:45]
  wire  Arbitration_3_io_valid_3_0; // @[Top_AO.scala 72:45]
  wire [31:0] Arbitration_3_io_node_id_3_1; // @[Top_AO.scala 72:45]
  wire [31:0] Arbitration_3_io_ray_id_3_1; // @[Top_AO.scala 72:45]
  wire [31:0] Arbitration_3_io_hit_3_1; // @[Top_AO.scala 72:45]
  wire  Arbitration_3_io_valid_3_1; // @[Top_AO.scala 72:45]
  wire [31:0] Arbitration_3_io_node_id_3_2; // @[Top_AO.scala 72:45]
  wire [31:0] Arbitration_3_io_ray_id_3_2; // @[Top_AO.scala 72:45]
  wire [31:0] Arbitration_3_io_hit_3_2; // @[Top_AO.scala 72:45]
  wire  Arbitration_3_io_valid_3_2; // @[Top_AO.scala 72:45]
  wire [31:0] Arbitration_3_io_node_id_3_3; // @[Top_AO.scala 72:45]
  wire [31:0] Arbitration_3_io_ray_id_3_3; // @[Top_AO.scala 72:45]
  wire [31:0] Arbitration_3_io_hit_3_3; // @[Top_AO.scala 72:45]
  wire  Arbitration_3_io_valid_3_3; // @[Top_AO.scala 72:45]
  wire [31:0] Arbitration_3_io_node_id_3_4; // @[Top_AO.scala 72:45]
  wire [31:0] Arbitration_3_io_ray_id_3_4; // @[Top_AO.scala 72:45]
  wire [31:0] Arbitration_3_io_hit_3_4; // @[Top_AO.scala 72:45]
  wire  Arbitration_3_io_valid_3_4; // @[Top_AO.scala 72:45]
  wire [31:0] Arbitration_3_io_node_id_out; // @[Top_AO.scala 72:45]
  wire [31:0] Arbitration_3_io_ray_id_out; // @[Top_AO.scala 72:45]
  wire [31:0] Arbitration_3_io_hit_out; // @[Top_AO.scala 72:45]
  wire  Arbitration_3_io_valid_out; // @[Top_AO.scala 72:45]
  wire  Arbitration_3_2_clock; // @[Top_AO.scala 73:42]
  wire  Arbitration_3_2_reset; // @[Top_AO.scala 73:42]
  wire [31:0] Arbitration_3_2_io_node_id_3_0; // @[Top_AO.scala 73:42]
  wire [31:0] Arbitration_3_2_io_ray_id_3_0; // @[Top_AO.scala 73:42]
  wire [31:0] Arbitration_3_2_io_hit_3_0; // @[Top_AO.scala 73:42]
  wire  Arbitration_3_2_io_valid_3_0; // @[Top_AO.scala 73:42]
  wire [31:0] Arbitration_3_2_io_node_id_3_1; // @[Top_AO.scala 73:42]
  wire [31:0] Arbitration_3_2_io_ray_id_3_1; // @[Top_AO.scala 73:42]
  wire [31:0] Arbitration_3_2_io_hit_3_1; // @[Top_AO.scala 73:42]
  wire  Arbitration_3_2_io_valid_3_1; // @[Top_AO.scala 73:42]
  wire [31:0] Arbitration_3_2_io_node_id_3_2; // @[Top_AO.scala 73:42]
  wire [31:0] Arbitration_3_2_io_ray_id_3_2; // @[Top_AO.scala 73:42]
  wire [31:0] Arbitration_3_2_io_hit_3_2; // @[Top_AO.scala 73:42]
  wire  Arbitration_3_2_io_valid_3_2; // @[Top_AO.scala 73:42]
  wire [31:0] Arbitration_3_2_io_node_id_3_3; // @[Top_AO.scala 73:42]
  wire [31:0] Arbitration_3_2_io_ray_id_3_3; // @[Top_AO.scala 73:42]
  wire [31:0] Arbitration_3_2_io_hit_3_3; // @[Top_AO.scala 73:42]
  wire  Arbitration_3_2_io_valid_3_3; // @[Top_AO.scala 73:42]
  wire [31:0] Arbitration_3_2_io_node_id_3_4; // @[Top_AO.scala 73:42]
  wire [31:0] Arbitration_3_2_io_ray_id_3_4; // @[Top_AO.scala 73:42]
  wire [31:0] Arbitration_3_2_io_hit_3_4; // @[Top_AO.scala 73:42]
  wire  Arbitration_3_2_io_valid_3_4; // @[Top_AO.scala 73:42]
  wire [31:0] Arbitration_3_2_io_node_id_out; // @[Top_AO.scala 73:42]
  wire [31:0] Arbitration_3_2_io_ray_id_out; // @[Top_AO.scala 73:42]
  wire [31:0] Arbitration_3_2_io_hit_out; // @[Top_AO.scala 73:42]
  wire  Arbitration_3_2_io_valid_out; // @[Top_AO.scala 73:42]
  wire  Arbitration_4_clock; // @[Top_AO.scala 74:45]
  wire  Arbitration_4_reset; // @[Top_AO.scala 74:45]
  wire [31:0] Arbitration_4_io_node_id_4_0; // @[Top_AO.scala 74:45]
  wire [31:0] Arbitration_4_io_ray_id_4_0; // @[Top_AO.scala 74:45]
  wire [31:0] Arbitration_4_io_hit_4_0; // @[Top_AO.scala 74:45]
  wire  Arbitration_4_io_valid_4_0; // @[Top_AO.scala 74:45]
  wire [31:0] Arbitration_4_io_node_id_4_1; // @[Top_AO.scala 74:45]
  wire [31:0] Arbitration_4_io_ray_id_4_1; // @[Top_AO.scala 74:45]
  wire [31:0] Arbitration_4_io_hit_4_1; // @[Top_AO.scala 74:45]
  wire  Arbitration_4_io_valid_4_1; // @[Top_AO.scala 74:45]
  wire [31:0] Arbitration_4_io_node_id_out; // @[Top_AO.scala 74:45]
  wire [31:0] Arbitration_4_io_ray_id_out; // @[Top_AO.scala 74:45]
  wire [31:0] Arbitration_4_io_hit_out; // @[Top_AO.scala 74:45]
  wire  Arbitration_4_io_RAY_AABB_out; // @[Top_AO.scala 74:45]
  wire  Arbitration_4_io_RAY_AABB_2_out; // @[Top_AO.scala 74:45]
  wire  Arbitration_4_io_valid_out; // @[Top_AO.scala 74:45]
  wire  Stack_manage_clock; // @[Top_AO.scala 76:41]
  wire  Stack_manage_reset; // @[Top_AO.scala 76:41]
  wire  Stack_manage_io_push; // @[Top_AO.scala 76:41]
  wire  Stack_manage_io_push_en; // @[Top_AO.scala 76:41]
  wire  Stack_manage_io_pop; // @[Top_AO.scala 76:41]
  wire  Stack_manage_io_pop_en; // @[Top_AO.scala 76:41]
  wire [31:0] Stack_manage_io_ray_id_push; // @[Top_AO.scala 76:41]
  wire [31:0] Stack_manage_io_ray_id_pop; // @[Top_AO.scala 76:41]
  wire [31:0] Stack_manage_io_node_id_push_in; // @[Top_AO.scala 76:41]
  wire [31:0] Stack_manage_io_hitT_in; // @[Top_AO.scala 76:41]
  wire  Stack_manage_io_clear; // @[Top_AO.scala 76:41]
  wire [31:0] Stack_manage_io_hitT_out; // @[Top_AO.scala 76:41]
  wire [31:0] Stack_manage_io_node_id_out; // @[Top_AO.scala 76:41]
  wire [31:0] Stack_manage_io_ray_id_out; // @[Top_AO.scala 76:41]
  wire  Stack_manage_io_pop_valid; // @[Top_AO.scala 76:41]
  wire  Stack_manage_io_Dis_en; // @[Top_AO.scala 76:41]
  wire  Stack_manage_io_Finish; // @[Top_AO.scala 76:41]
  wire  Stack_manage_2_clock; // @[Top_AO.scala 77:38]
  wire  Stack_manage_2_reset; // @[Top_AO.scala 77:38]
  wire  Stack_manage_2_io_push; // @[Top_AO.scala 77:38]
  wire  Stack_manage_2_io_push_en; // @[Top_AO.scala 77:38]
  wire  Stack_manage_2_io_pop; // @[Top_AO.scala 77:38]
  wire  Stack_manage_2_io_pop_en; // @[Top_AO.scala 77:38]
  wire [31:0] Stack_manage_2_io_ray_id_push; // @[Top_AO.scala 77:38]
  wire [31:0] Stack_manage_2_io_ray_id_pop; // @[Top_AO.scala 77:38]
  wire [31:0] Stack_manage_2_io_node_id_push_in; // @[Top_AO.scala 77:38]
  wire [31:0] Stack_manage_2_io_hitT_in; // @[Top_AO.scala 77:38]
  wire  Stack_manage_2_io_clear; // @[Top_AO.scala 77:38]
  wire [31:0] Stack_manage_2_io_hitT_out; // @[Top_AO.scala 77:38]
  wire [31:0] Stack_manage_2_io_node_id_out; // @[Top_AO.scala 77:38]
  wire [31:0] Stack_manage_2_io_ray_id_out; // @[Top_AO.scala 77:38]
  wire  Stack_manage_2_io_pop_valid; // @[Top_AO.scala 77:38]
  wire  Stack_manage_2_io_Dis_en; // @[Top_AO.scala 77:38]
  wire  Stack_manage_2_io_Finish; // @[Top_AO.scala 77:38]
  wire  Triangle_clock; // @[Top_AO.scala 78:51]
  wire  Triangle_reset; // @[Top_AO.scala 78:51]
  wire  Triangle_io_To_IST0_enable; // @[Top_AO.scala 78:51]
  wire [31:0] Triangle_io_nodeid_leaf; // @[Top_AO.scala 78:51]
  wire [31:0] Triangle_io_rayid_leaf; // @[Top_AO.scala 78:51]
  wire [31:0] Triangle_io_hiT_in; // @[Top_AO.scala 78:51]
  wire [31:0] Triangle_io_v00_in_x; // @[Top_AO.scala 78:51]
  wire [31:0] Triangle_io_v00_in_y; // @[Top_AO.scala 78:51]
  wire [31:0] Triangle_io_v00_in_z; // @[Top_AO.scala 78:51]
  wire [31:0] Triangle_io_v00_in_w; // @[Top_AO.scala 78:51]
  wire [31:0] Triangle_io_v11_in_x; // @[Top_AO.scala 78:51]
  wire [31:0] Triangle_io_v11_in_y; // @[Top_AO.scala 78:51]
  wire [31:0] Triangle_io_v11_in_z; // @[Top_AO.scala 78:51]
  wire [31:0] Triangle_io_v11_in_w; // @[Top_AO.scala 78:51]
  wire [31:0] Triangle_io_v22_in_x; // @[Top_AO.scala 78:51]
  wire [31:0] Triangle_io_v22_in_y; // @[Top_AO.scala 78:51]
  wire [31:0] Triangle_io_v22_in_z; // @[Top_AO.scala 78:51]
  wire [31:0] Triangle_io_v22_in_w; // @[Top_AO.scala 78:51]
  wire [31:0] Triangle_io_ray_o_in_x; // @[Top_AO.scala 78:51]
  wire [31:0] Triangle_io_ray_o_in_y; // @[Top_AO.scala 78:51]
  wire [31:0] Triangle_io_ray_o_in_z; // @[Top_AO.scala 78:51]
  wire [31:0] Triangle_io_ray_d_in_x; // @[Top_AO.scala 78:51]
  wire [31:0] Triangle_io_ray_d_in_y; // @[Top_AO.scala 78:51]
  wire [31:0] Triangle_io_ray_d_in_z; // @[Top_AO.scala 78:51]
  wire  Triangle_io_break_in; // @[Top_AO.scala 78:51]
  wire  Triangle_io_RAY_AABB_1; // @[Top_AO.scala 78:51]
  wire  Triangle_io_RAY_AABB_2; // @[Top_AO.scala 78:51]
  wire  Triangle_io_pop_1; // @[Top_AO.scala 78:51]
  wire  Triangle_io_break_1; // @[Top_AO.scala 78:51]
  wire  Triangle_io_pop_2; // @[Top_AO.scala 78:51]
  wire  Triangle_io_break_2; // @[Top_AO.scala 78:51]
  wire  Triangle_io_pop_3; // @[Top_AO.scala 78:51]
  wire  Triangle_io_break_3; // @[Top_AO.scala 78:51]
  wire [31:0] Triangle_io_hiT_out_1; // @[Top_AO.scala 78:51]
  wire [31:0] Triangle_io_hiT_out_2; // @[Top_AO.scala 78:51]
  wire [31:0] Triangle_io_hiT_out_3; // @[Top_AO.scala 78:51]
  wire  Triangle_io_hitT_en; // @[Top_AO.scala 78:51]
  wire [31:0] Triangle_io_hitIndex; // @[Top_AO.scala 78:51]
  wire  Triangle_io_hitIndex_en; // @[Top_AO.scala 78:51]
  wire [31:0] Triangle_io_node_id_out_1; // @[Top_AO.scala 78:51]
  wire [31:0] Triangle_io_node_id_out_2; // @[Top_AO.scala 78:51]
  wire [31:0] Triangle_io_node_id_out_3; // @[Top_AO.scala 78:51]
  wire [31:0] Triangle_io_ray_id_ist1; // @[Top_AO.scala 78:51]
  wire [31:0] Triangle_io_ray_id_ist2; // @[Top_AO.scala 78:51]
  wire [31:0] Triangle_io_ray_id_ist3; // @[Top_AO.scala 78:51]
  wire [63:0] Triangle_io_counter_fdiv; // @[Top_AO.scala 78:51]
  wire  Triangle_io_RAY_AABB_1_out_IST1; // @[Top_AO.scala 78:51]
  wire  Triangle_io_RAY_AABB_2_out_IST1; // @[Top_AO.scala 78:51]
  wire  Triangle_io_RAY_AABB_1_out_IST2; // @[Top_AO.scala 78:51]
  wire  Triangle_io_RAY_AABB_2_out_IST2; // @[Top_AO.scala 78:51]
  wire  Triangle_io_RAY_AABB_1_out_IST3; // @[Top_AO.scala 78:51]
  wire  Triangle_io_RAY_AABB_2_out_IST3; // @[Top_AO.scala 78:51]
  reg [63:0] clock_counter; // @[Top_AO.scala 80:42]
  wire [63:0] _T_1 = clock_counter + 64'h1; // @[Top_AO.scala 81:53]
  reg  memory_valid; // @[Top_AO.scala 135:54]
  reg [31:0] hit_temp; // @[Top_AO.scala 136:61]
  reg [31:0] ray_id_temp; // @[Top_AO.scala 137:57]
  reg  hit_from_arb; // @[Top_AO.scala 138:57]
  reg [63:0] TRV_1; // @[Top_AO.scala 139:64]
  wire  _T_14 = Arbitration_1_io_valid_out & Arbitration_1_io_hit_out != 32'h0; // @[Top_AO.scala 140:36]
  wire [32:0] _T_15 = $signed(Arbitration_1_io_node_id_out) / 32'sh4; // @[Top_AO.scala 149:75]
  wire  _T_30 = Arbitration_1_io_valid_out & Arbitration_1_io_hit_out == 32'h0; // @[Top_AO.scala 165:42]
  wire [31:0] _GEN_13 = Arbitration_1_io_ray_id_out; // @[Top_AO.scala 165:76 Top_AO.scala 167:53]
  wire  _GEN_31 = Arbitration_1_io_valid_out & Arbitration_1_io_hit_out != 32'h0 | _T_30; // @[Top_AO.scala 140:70 Top_AO.scala 141:51]
  wire [32:0] _GEN_34 = Arbitration_1_io_valid_out & Arbitration_1_io_hit_out != 32'h0 ? $signed(_T_15) : $signed(_T_15)
    ; // @[Top_AO.scala 140:70 Top_AO.scala 149:44]
  wire [31:0] _GEN_51 = hit_from_arb ? hit_temp : Ray_hitT_io_Ray_out; // @[Top_AO.scala 204:33 Top_AO.scala 205:53 Top_AO.scala 207:53]
  wire [63:0] _T_48 = TRV_1 + 64'h1; // @[Top_AO.scala 228:79]
  reg  memory_valid_2; // @[Top_AO.scala 270:56]
  reg [31:0] hit_temp_2; // @[Top_AO.scala 271:63]
  reg [31:0] ray_id_temp_2; // @[Top_AO.scala 272:59]
  reg  hit_from_arb_2; // @[Top_AO.scala 273:59]
  reg [63:0] TRV_2; // @[Top_AO.scala 274:70]
  wire  _T_51 = Arbitration_1_2_io_valid_out & Arbitration_1_2_io_hit_out != 32'h0; // @[Top_AO.scala 275:38]
  wire [32:0] _T_52 = $signed(Arbitration_1_2_io_node_id_out) / 32'sh4; // @[Top_AO.scala 286:79]
  wire  _T_67 = Arbitration_1_2_io_valid_out & Arbitration_1_2_io_hit_out == 32'h0; // @[Top_AO.scala 302:44]
  wire [31:0] _GEN_81 = Arbitration_1_2_io_ray_id_out; // @[Top_AO.scala 302:80 Top_AO.scala 306:54]
  wire  _GEN_98 = Arbitration_1_2_io_valid_out & Arbitration_1_2_io_hit_out != 32'h0 | _T_67; // @[Top_AO.scala 275:74 Top_AO.scala 276:58]
  wire [32:0] _GEN_101 = Arbitration_1_2_io_valid_out & Arbitration_1_2_io_hit_out != 32'h0 ? $signed(_T_52) : $signed(
    _T_52); // @[Top_AO.scala 275:74 Top_AO.scala 286:46]
  wire [31:0] _GEN_118 = hit_from_arb_2 ? hit_temp_2 : Ray_hitT_io_Ray_out_2; // @[Top_AO.scala 343:35 Top_AO.scala 344:55 Top_AO.scala 346:55]
  wire [63:0] _T_85 = TRV_2 + 64'h1; // @[Top_AO.scala 364:85]
  wire  hi = ~RAY_AABB_io_nodeIdx_2[31]; // @[common.scala 128:29]
  wire [30:0] lo = ~RAY_AABB_io_nodeIdx_2[30:0]; // @[common.scala 128:45]
  wire [31:0] _T_94 = {hi,lo}; // @[common.scala 128:56]
  wire  hi_1 = ~RAY_AABB_2_io_nodeIdx_2[31]; // @[common.scala 128:29]
  wire [30:0] lo_1 = ~RAY_AABB_2_io_nodeIdx_2[30:0]; // @[common.scala 128:45]
  wire [31:0] _T_100 = {hi_1,lo_1}; // @[common.scala 128:56]
  wire  _T_102 = ~Stack_manage_io_node_id_out[31]; // @[common.scala 100:25]
  wire [30:0] lo_2 = ~Stack_manage_io_node_id_out[30:0]; // @[common.scala 128:45]
  wire [31:0] _T_115 = {_T_102,lo_2}; // @[common.scala 128:56]
  wire [31:0] _GEN_168 = _T_102 & Stack_manage_io_pop_valid ? Stack_manage_io_ray_id_out : 32'h0; // @[Top_AO.scala 457:81 Top_AO.scala 459:50]
  wire  _T_117 = ~Stack_manage_2_io_node_id_out[31]; // @[common.scala 100:25]
  wire [30:0] lo_3 = ~Stack_manage_2_io_node_id_out[30:0]; // @[common.scala 128:45]
  wire [31:0] _T_130 = {_T_117,lo_3}; // @[common.scala 128:56]
  wire [31:0] _GEN_182 = _T_117 & Stack_manage_2_io_pop_valid ? Stack_manage_2_io_ray_id_out : 32'h0; // @[Top_AO.scala 477:85 Top_AO.scala 479:52]
  wire [31:0] _T_134 = $signed(Triangle_io_node_id_out_1) + 32'sh3; // @[Top_AO.scala 523:71]
  wire [31:0] _T_142 = $signed(Triangle_io_node_id_out_2) + 32'sh3; // @[Top_AO.scala 548:71]
  wire [31:0] _T_150 = $signed(Triangle_io_node_id_out_3) + 32'sh3; // @[Top_AO.scala 572:71]
  reg  leaf_memory_valid; // @[Top_AO.scala 672:58]
  reg [31:0] hitT_temp; // @[Top_AO.scala 673:68]
  reg [31:0] ray_leaf_temp; // @[Top_AO.scala 674:64]
  reg [31:0] leaf_node_id_temp; // @[Top_AO.scala 675:57]
  reg  ray_aabb; // @[Top_AO.scala 676:69]
  reg  ray_aabb_2; // @[Top_AO.scala 677:71]
  reg [63:0] IST_1; // @[Top_AO.scala 678:75]
  wire  _GEN_239 = Arbitration_4_io_valid_out; // @[Top_AO.scala 679:37 Top_AO.scala 680:50 Top_AO.scala 697:50]
  wire  _GEN_245 = Arbitration_4_io_valid_out & Arbitration_4_io_RAY_AABB_out; // @[Top_AO.scala 679:37 Top_AO.scala 694:64 Top_AO.scala 701:64]
  wire  _GEN_246 = Arbitration_4_io_valid_out & Arbitration_4_io_RAY_AABB_2_out; // @[Top_AO.scala 679:37 Top_AO.scala 695:61 Top_AO.scala 702:61]
  wire [63:0] _T_165 = IST_1 + 64'h1; // @[Top_AO.scala 730:76]
  ray_dispatch Ray_Dispatch ( // @[Top_AO.scala 24:44]
    .clock(Ray_Dispatch_clock),
    .reset(Ray_Dispatch_reset),
    .io_dispatch(Ray_Dispatch_io_dispatch),
    .io_dispatch_2(Ray_Dispatch_io_dispatch_2),
    .io_rayid_id(Ray_Dispatch_io_rayid_id),
    .io_rayid_id_2(Ray_Dispatch_io_rayid_id_2),
    .io_ray_out(Ray_Dispatch_io_ray_out),
    .io_ray_out_2(Ray_Dispatch_io_ray_out_2),
    .io_ray_finish(Ray_Dispatch_io_ray_finish)
  );
  ray_memory Ray_origx ( // @[Top_AO.scala 25:48]
    .clock(Ray_origx_clock),
    .io_Ray_id(Ray_origx_io_Ray_id),
    .io_Ray_id_2(Ray_origx_io_Ray_id_2),
    .io_Ray_out(Ray_origx_io_Ray_out),
    .io_Ray_out_2(Ray_origx_io_Ray_out_2)
  );
  ray_memory Ray_origy ( // @[Top_AO.scala 26:48]
    .clock(Ray_origy_clock),
    .io_Ray_id(Ray_origy_io_Ray_id),
    .io_Ray_id_2(Ray_origy_io_Ray_id_2),
    .io_Ray_out(Ray_origy_io_Ray_out),
    .io_Ray_out_2(Ray_origy_io_Ray_out_2)
  );
  ray_memory Ray_origz ( // @[Top_AO.scala 27:48]
    .clock(Ray_origz_clock),
    .io_Ray_id(Ray_origz_io_Ray_id),
    .io_Ray_id_2(Ray_origz_io_Ray_id_2),
    .io_Ray_out(Ray_origz_io_Ray_out),
    .io_Ray_out_2(Ray_origz_io_Ray_out_2)
  );
  ray_memory Ray_dirx ( // @[Top_AO.scala 30:50]
    .clock(Ray_dirx_clock),
    .io_Ray_id(Ray_dirx_io_Ray_id),
    .io_Ray_id_2(Ray_dirx_io_Ray_id_2),
    .io_Ray_out(Ray_dirx_io_Ray_out),
    .io_Ray_out_2(Ray_dirx_io_Ray_out_2)
  );
  ray_memory Ray_diry ( // @[Top_AO.scala 31:49]
    .clock(Ray_diry_clock),
    .io_Ray_id(Ray_diry_io_Ray_id),
    .io_Ray_id_2(Ray_diry_io_Ray_id_2),
    .io_Ray_out(Ray_diry_io_Ray_out),
    .io_Ray_out_2(Ray_diry_io_Ray_out_2)
  );
  ray_memory Ray_dirz ( // @[Top_AO.scala 32:49]
    .clock(Ray_dirz_clock),
    .io_Ray_id(Ray_dirz_io_Ray_id),
    .io_Ray_id_2(Ray_dirz_io_Ray_id_2),
    .io_Ray_out(Ray_dirz_io_Ray_out),
    .io_Ray_out_2(Ray_dirz_io_Ray_out_2)
  );
  ray_memory Ray_hitT ( // @[Top_AO.scala 33:49]
    .clock(Ray_hitT_clock),
    .io_Ray_id(Ray_hitT_io_Ray_id),
    .io_Ray_id_2(Ray_hitT_io_Ray_id_2),
    .io_Ray_out(Ray_hitT_io_Ray_out),
    .io_Ray_out_2(Ray_hitT_io_Ray_out_2)
  );
  ray_memory Ray_idirx ( // @[Top_AO.scala 35:49]
    .clock(Ray_idirx_clock),
    .io_Ray_id(Ray_idirx_io_Ray_id),
    .io_Ray_id_2(Ray_idirx_io_Ray_id_2),
    .io_Ray_out(Ray_idirx_io_Ray_out),
    .io_Ray_out_2(Ray_idirx_io_Ray_out_2)
  );
  ray_memory Ray_idiry ( // @[Top_AO.scala 36:49]
    .clock(Ray_idiry_clock),
    .io_Ray_id(Ray_idiry_io_Ray_id),
    .io_Ray_id_2(Ray_idiry_io_Ray_id_2),
    .io_Ray_out(Ray_idiry_io_Ray_out),
    .io_Ray_out_2(Ray_idiry_io_Ray_out_2)
  );
  ray_memory Ray_idirz ( // @[Top_AO.scala 37:49]
    .clock(Ray_idirz_clock),
    .io_Ray_id(Ray_idirz_io_Ray_id),
    .io_Ray_id_2(Ray_idirz_io_Ray_id_2),
    .io_Ray_out(Ray_idirz_io_Ray_out),
    .io_Ray_out_2(Ray_idirz_io_Ray_out_2)
  );
  ray_memory Ray_oodx ( // @[Top_AO.scala 39:48]
    .clock(Ray_oodx_clock),
    .io_Ray_id(Ray_oodx_io_Ray_id),
    .io_Ray_id_2(Ray_oodx_io_Ray_id_2),
    .io_Ray_out(Ray_oodx_io_Ray_out),
    .io_Ray_out_2(Ray_oodx_io_Ray_out_2)
  );
  ray_memory Ray_oody ( // @[Top_AO.scala 40:48]
    .clock(Ray_oody_clock),
    .io_Ray_id(Ray_oody_io_Ray_id),
    .io_Ray_id_2(Ray_oody_io_Ray_id_2),
    .io_Ray_out(Ray_oody_io_Ray_out),
    .io_Ray_out_2(Ray_oody_io_Ray_out_2)
  );
  ray_memory Ray_oodz ( // @[Top_AO.scala 41:48]
    .clock(Ray_oodz_clock),
    .io_Ray_id(Ray_oodz_io_Ray_id),
    .io_Ray_id_2(Ray_oodz_io_Ray_id_2),
    .io_Ray_out(Ray_oodz_io_Ray_out),
    .io_Ray_out_2(Ray_oodz_io_Ray_out_2)
  );
  BVH_memory BVH_RAM_0_x ( // @[Top_AO.scala 43:41]
    .clock(BVH_RAM_0_x_clock),
    .io_BVH_id(BVH_RAM_0_x_io_BVH_id),
    .io_BVH_id_2(BVH_RAM_0_x_io_BVH_id_2),
    .io_BVH_out(BVH_RAM_0_x_io_BVH_out),
    .io_BVH_out_2(BVH_RAM_0_x_io_BVH_out_2)
  );
  BVH_memory BVH_RAM_0_y ( // @[Top_AO.scala 44:41]
    .clock(BVH_RAM_0_y_clock),
    .io_BVH_id(BVH_RAM_0_y_io_BVH_id),
    .io_BVH_id_2(BVH_RAM_0_y_io_BVH_id_2),
    .io_BVH_out(BVH_RAM_0_y_io_BVH_out),
    .io_BVH_out_2(BVH_RAM_0_y_io_BVH_out_2)
  );
  BVH_memory BVH_RAM_0_z ( // @[Top_AO.scala 45:41]
    .clock(BVH_RAM_0_z_clock),
    .io_BVH_id(BVH_RAM_0_z_io_BVH_id),
    .io_BVH_id_2(BVH_RAM_0_z_io_BVH_id_2),
    .io_BVH_out(BVH_RAM_0_z_io_BVH_out),
    .io_BVH_out_2(BVH_RAM_0_z_io_BVH_out_2)
  );
  BVH_memory BVH_RAM_0_w ( // @[Top_AO.scala 46:40]
    .clock(BVH_RAM_0_w_clock),
    .io_BVH_id(BVH_RAM_0_w_io_BVH_id),
    .io_BVH_id_2(BVH_RAM_0_w_io_BVH_id_2),
    .io_BVH_out(BVH_RAM_0_w_io_BVH_out),
    .io_BVH_out_2(BVH_RAM_0_w_io_BVH_out_2)
  );
  BVH_memory BVH_RAM_1_x ( // @[Top_AO.scala 48:41]
    .clock(BVH_RAM_1_x_clock),
    .io_BVH_id(BVH_RAM_1_x_io_BVH_id),
    .io_BVH_id_2(BVH_RAM_1_x_io_BVH_id_2),
    .io_BVH_out(BVH_RAM_1_x_io_BVH_out),
    .io_BVH_out_2(BVH_RAM_1_x_io_BVH_out_2)
  );
  BVH_memory BVH_RAM_1_y ( // @[Top_AO.scala 49:41]
    .clock(BVH_RAM_1_y_clock),
    .io_BVH_id(BVH_RAM_1_y_io_BVH_id),
    .io_BVH_id_2(BVH_RAM_1_y_io_BVH_id_2),
    .io_BVH_out(BVH_RAM_1_y_io_BVH_out),
    .io_BVH_out_2(BVH_RAM_1_y_io_BVH_out_2)
  );
  BVH_memory BVH_RAM_1_z ( // @[Top_AO.scala 50:41]
    .clock(BVH_RAM_1_z_clock),
    .io_BVH_id(BVH_RAM_1_z_io_BVH_id),
    .io_BVH_id_2(BVH_RAM_1_z_io_BVH_id_2),
    .io_BVH_out(BVH_RAM_1_z_io_BVH_out),
    .io_BVH_out_2(BVH_RAM_1_z_io_BVH_out_2)
  );
  BVH_memory BVH_RAM_1_w ( // @[Top_AO.scala 51:40]
    .clock(BVH_RAM_1_w_clock),
    .io_BVH_id(BVH_RAM_1_w_io_BVH_id),
    .io_BVH_id_2(BVH_RAM_1_w_io_BVH_id_2),
    .io_BVH_out(BVH_RAM_1_w_io_BVH_out),
    .io_BVH_out_2(BVH_RAM_1_w_io_BVH_out_2)
  );
  BVH_memory BVH_RAM_z_x ( // @[Top_AO.scala 53:41]
    .clock(BVH_RAM_z_x_clock),
    .io_BVH_id(BVH_RAM_z_x_io_BVH_id),
    .io_BVH_id_2(BVH_RAM_z_x_io_BVH_id_2),
    .io_BVH_out(BVH_RAM_z_x_io_BVH_out),
    .io_BVH_out_2(BVH_RAM_z_x_io_BVH_out_2)
  );
  BVH_memory BVH_RAM_z_y ( // @[Top_AO.scala 54:41]
    .clock(BVH_RAM_z_y_clock),
    .io_BVH_id(BVH_RAM_z_y_io_BVH_id),
    .io_BVH_id_2(BVH_RAM_z_y_io_BVH_id_2),
    .io_BVH_out(BVH_RAM_z_y_io_BVH_out),
    .io_BVH_out_2(BVH_RAM_z_y_io_BVH_out_2)
  );
  BVH_memory BVH_RAM_z_z ( // @[Top_AO.scala 55:41]
    .clock(BVH_RAM_z_z_clock),
    .io_BVH_id(BVH_RAM_z_z_io_BVH_id),
    .io_BVH_id_2(BVH_RAM_z_z_io_BVH_id_2),
    .io_BVH_out(BVH_RAM_z_z_io_BVH_out),
    .io_BVH_out_2(BVH_RAM_z_z_io_BVH_out_2)
  );
  BVH_memory BVH_RAM_z_w ( // @[Top_AO.scala 56:40]
    .clock(BVH_RAM_z_w_clock),
    .io_BVH_id(BVH_RAM_z_w_io_BVH_id),
    .io_BVH_id_2(BVH_RAM_z_w_io_BVH_id_2),
    .io_BVH_out(BVH_RAM_z_w_io_BVH_out),
    .io_BVH_out_2(BVH_RAM_z_w_io_BVH_out_2)
  );
  BVH_memory_0 BVH_RAM_tmp_x ( // @[Top_AO.scala 58:37]
    .clock(BVH_RAM_tmp_x_clock),
    .io_BVH_id(BVH_RAM_tmp_x_io_BVH_id),
    .io_BVH_id_2(BVH_RAM_tmp_x_io_BVH_id_2),
    .io_BVH_out(BVH_RAM_tmp_x_io_BVH_out),
    .io_BVH_out_2(BVH_RAM_tmp_x_io_BVH_out_2)
  );
  BVH_memory_0 BVH_RAM_tmp_y ( // @[Top_AO.scala 59:37]
    .clock(BVH_RAM_tmp_y_clock),
    .io_BVH_id(BVH_RAM_tmp_y_io_BVH_id),
    .io_BVH_id_2(BVH_RAM_tmp_y_io_BVH_id_2),
    .io_BVH_out(BVH_RAM_tmp_y_io_BVH_out),
    .io_BVH_out_2(BVH_RAM_tmp_y_io_BVH_out_2)
  );
  Triangle_memory_valid TRI_RAM_x ( // @[Top_AO.scala 61:50]
    .clock(TRI_RAM_x_clock),
    .io_Triangle_id(TRI_RAM_x_io_Triangle_id),
    .io_v00_out(TRI_RAM_x_io_v00_out),
    .io_v11_out(TRI_RAM_x_io_v11_out),
    .io_v22_out(TRI_RAM_x_io_v22_out),
    .io_valid(TRI_RAM_x_io_valid)
  );
  Triangle_memory TRI_RAM_y ( // @[Top_AO.scala 62:50]
    .clock(TRI_RAM_y_clock),
    .io_Triangle_id(TRI_RAM_y_io_Triangle_id),
    .io_v00_out(TRI_RAM_y_io_v00_out),
    .io_v11_out(TRI_RAM_y_io_v11_out),
    .io_v22_out(TRI_RAM_y_io_v22_out)
  );
  Triangle_memory TRI_RAM_z ( // @[Top_AO.scala 63:50]
    .clock(TRI_RAM_z_clock),
    .io_Triangle_id(TRI_RAM_z_io_Triangle_id),
    .io_v00_out(TRI_RAM_z_io_v00_out),
    .io_v11_out(TRI_RAM_z_io_v11_out),
    .io_v22_out(TRI_RAM_z_io_v22_out)
  );
  Triangle_memory TRI_RAM_w ( // @[Top_AO.scala 64:49]
    .clock(TRI_RAM_w_clock),
    .io_Triangle_id(TRI_RAM_w_io_Triangle_id),
    .io_v00_out(TRI_RAM_w_io_v00_out),
    .io_v11_out(TRI_RAM_w_io_v11_out),
    .io_v22_out(TRI_RAM_w_io_v22_out)
  );
  ray_AABB_1 RAY_AABB ( // @[Top_AO.scala 65:46]
    .clock(RAY_AABB_clock),
    .reset(RAY_AABB_reset),
    .io_ray_idir_x(RAY_AABB_io_ray_idir_x),
    .io_ray_idir_y(RAY_AABB_io_ray_idir_y),
    .io_ray_idir_z(RAY_AABB_io_ray_idir_z),
    .io_ray_ood_x(RAY_AABB_io_ray_ood_x),
    .io_ray_ood_y(RAY_AABB_io_ray_ood_y),
    .io_ray_ood_z(RAY_AABB_io_ray_ood_z),
    .io_ray_hitT(RAY_AABB_io_ray_hitT),
    .io_bvh_n0xy_x(RAY_AABB_io_bvh_n0xy_x),
    .io_bvh_n0xy_y(RAY_AABB_io_bvh_n0xy_y),
    .io_bvh_n0xy_z(RAY_AABB_io_bvh_n0xy_z),
    .io_bvh_n0xy_w(RAY_AABB_io_bvh_n0xy_w),
    .io_bvh_n1xy_x(RAY_AABB_io_bvh_n1xy_x),
    .io_bvh_n1xy_y(RAY_AABB_io_bvh_n1xy_y),
    .io_bvh_n1xy_z(RAY_AABB_io_bvh_n1xy_z),
    .io_bvh_n1xy_w(RAY_AABB_io_bvh_n1xy_w),
    .io_bvh_nz_x(RAY_AABB_io_bvh_nz_x),
    .io_bvh_nz_y(RAY_AABB_io_bvh_nz_y),
    .io_bvh_nz_z(RAY_AABB_io_bvh_nz_z),
    .io_bvh_nz_w(RAY_AABB_io_bvh_nz_w),
    .io_bvh_temp_x(RAY_AABB_io_bvh_temp_x),
    .io_bvh_temp_y(RAY_AABB_io_bvh_temp_y),
    .io_rayid(RAY_AABB_io_rayid),
    .io_valid_en(RAY_AABB_io_valid_en),
    .io_rayid_out(RAY_AABB_io_rayid_out),
    .io_nodeIdx_0(RAY_AABB_io_nodeIdx_0),
    .io_nodeIdx_1(RAY_AABB_io_nodeIdx_1),
    .io_nodeIdx_2(RAY_AABB_io_nodeIdx_2),
    .io_push(RAY_AABB_io_push),
    .io_pop(RAY_AABB_io_pop),
    .io_leaf(RAY_AABB_io_leaf),
    .io_back(RAY_AABB_io_back),
    .io_hitT_out(RAY_AABB_io_hitT_out),
    .io_valid_out(RAY_AABB_io_valid_out)
  );
  ray_AABB_1 RAY_AABB_2 ( // @[Top_AO.scala 66:48]
    .clock(RAY_AABB_2_clock),
    .reset(RAY_AABB_2_reset),
    .io_ray_idir_x(RAY_AABB_2_io_ray_idir_x),
    .io_ray_idir_y(RAY_AABB_2_io_ray_idir_y),
    .io_ray_idir_z(RAY_AABB_2_io_ray_idir_z),
    .io_ray_ood_x(RAY_AABB_2_io_ray_ood_x),
    .io_ray_ood_y(RAY_AABB_2_io_ray_ood_y),
    .io_ray_ood_z(RAY_AABB_2_io_ray_ood_z),
    .io_ray_hitT(RAY_AABB_2_io_ray_hitT),
    .io_bvh_n0xy_x(RAY_AABB_2_io_bvh_n0xy_x),
    .io_bvh_n0xy_y(RAY_AABB_2_io_bvh_n0xy_y),
    .io_bvh_n0xy_z(RAY_AABB_2_io_bvh_n0xy_z),
    .io_bvh_n0xy_w(RAY_AABB_2_io_bvh_n0xy_w),
    .io_bvh_n1xy_x(RAY_AABB_2_io_bvh_n1xy_x),
    .io_bvh_n1xy_y(RAY_AABB_2_io_bvh_n1xy_y),
    .io_bvh_n1xy_z(RAY_AABB_2_io_bvh_n1xy_z),
    .io_bvh_n1xy_w(RAY_AABB_2_io_bvh_n1xy_w),
    .io_bvh_nz_x(RAY_AABB_2_io_bvh_nz_x),
    .io_bvh_nz_y(RAY_AABB_2_io_bvh_nz_y),
    .io_bvh_nz_z(RAY_AABB_2_io_bvh_nz_z),
    .io_bvh_nz_w(RAY_AABB_2_io_bvh_nz_w),
    .io_bvh_temp_x(RAY_AABB_2_io_bvh_temp_x),
    .io_bvh_temp_y(RAY_AABB_2_io_bvh_temp_y),
    .io_rayid(RAY_AABB_2_io_rayid),
    .io_valid_en(RAY_AABB_2_io_valid_en),
    .io_rayid_out(RAY_AABB_2_io_rayid_out),
    .io_nodeIdx_0(RAY_AABB_2_io_nodeIdx_0),
    .io_nodeIdx_1(RAY_AABB_2_io_nodeIdx_1),
    .io_nodeIdx_2(RAY_AABB_2_io_nodeIdx_2),
    .io_push(RAY_AABB_2_io_push),
    .io_pop(RAY_AABB_2_io_pop),
    .io_leaf(RAY_AABB_2_io_leaf),
    .io_back(RAY_AABB_2_io_back),
    .io_hitT_out(RAY_AABB_2_io_hitT_out),
    .io_valid_out(RAY_AABB_2_io_valid_out)
  );
  Arbitration_1 Arbitration_1 ( // @[Top_AO.scala 67:50]
    .clock(Arbitration_1_clock),
    .reset(Arbitration_1_reset),
    .io_node_id_0(Arbitration_1_io_node_id_0),
    .io_ray_id_0(Arbitration_1_io_ray_id_0),
    .io_hit_0(Arbitration_1_io_hit_0),
    .io_valid_0(Arbitration_1_io_valid_0),
    .io_node_id_1(Arbitration_1_io_node_id_1),
    .io_ray_id_1(Arbitration_1_io_ray_id_1),
    .io_valid_1(Arbitration_1_io_valid_1),
    .io_ray_id_2(Arbitration_1_io_ray_id_2),
    .io_valid_2(Arbitration_1_io_valid_2),
    .io_node_id_out(Arbitration_1_io_node_id_out),
    .io_ray_id_out(Arbitration_1_io_ray_id_out),
    .io_hit_out(Arbitration_1_io_hit_out),
    .io_valid_out(Arbitration_1_io_valid_out)
  );
  Arbitration_1 Arbitration_1_2 ( // @[Top_AO.scala 68:47]
    .clock(Arbitration_1_2_clock),
    .reset(Arbitration_1_2_reset),
    .io_node_id_0(Arbitration_1_2_io_node_id_0),
    .io_ray_id_0(Arbitration_1_2_io_ray_id_0),
    .io_hit_0(Arbitration_1_2_io_hit_0),
    .io_valid_0(Arbitration_1_2_io_valid_0),
    .io_node_id_1(Arbitration_1_2_io_node_id_1),
    .io_ray_id_1(Arbitration_1_2_io_ray_id_1),
    .io_valid_1(Arbitration_1_2_io_valid_1),
    .io_ray_id_2(Arbitration_1_2_io_ray_id_2),
    .io_valid_2(Arbitration_1_2_io_valid_2),
    .io_node_id_out(Arbitration_1_2_io_node_id_out),
    .io_ray_id_out(Arbitration_1_2_io_ray_id_out),
    .io_hit_out(Arbitration_1_2_io_hit_out),
    .io_valid_out(Arbitration_1_2_io_valid_out)
  );
  Arbitration_2_1 Arbitration_2 ( // @[Top_AO.scala 70:45]
    .clock(Arbitration_2_clock),
    .reset(Arbitration_2_reset),
    .io_ray_id_2_0(Arbitration_2_io_ray_id_2_0),
    .io_hit_2_0(Arbitration_2_io_hit_2_0),
    .io_valid_2_0(Arbitration_2_io_valid_2_0),
    .io_ray_id_2_1(Arbitration_2_io_ray_id_2_1),
    .io_hit_2_1(Arbitration_2_io_hit_2_1),
    .io_valid_2_1(Arbitration_2_io_valid_2_1),
    .io_ray_id_2_2(Arbitration_2_io_ray_id_2_2),
    .io_hit_2_2(Arbitration_2_io_hit_2_2),
    .io_valid_2_2(Arbitration_2_io_valid_2_2),
    .io_ray_id_2_3(Arbitration_2_io_ray_id_2_3),
    .io_hit_2_3(Arbitration_2_io_hit_2_3),
    .io_valid_2_3(Arbitration_2_io_valid_2_3),
    .io_ray_id_out(Arbitration_2_io_ray_id_out),
    .io_hit_out(Arbitration_2_io_hit_out),
    .io_valid_out(Arbitration_2_io_valid_out)
  );
  Arbitration_2_1 Arbitration_2_2 ( // @[Top_AO.scala 71:42]
    .clock(Arbitration_2_2_clock),
    .reset(Arbitration_2_2_reset),
    .io_ray_id_2_0(Arbitration_2_2_io_ray_id_2_0),
    .io_hit_2_0(Arbitration_2_2_io_hit_2_0),
    .io_valid_2_0(Arbitration_2_2_io_valid_2_0),
    .io_ray_id_2_1(Arbitration_2_2_io_ray_id_2_1),
    .io_hit_2_1(Arbitration_2_2_io_hit_2_1),
    .io_valid_2_1(Arbitration_2_2_io_valid_2_1),
    .io_ray_id_2_2(Arbitration_2_2_io_ray_id_2_2),
    .io_hit_2_2(Arbitration_2_2_io_hit_2_2),
    .io_valid_2_2(Arbitration_2_2_io_valid_2_2),
    .io_ray_id_2_3(Arbitration_2_2_io_ray_id_2_3),
    .io_hit_2_3(Arbitration_2_2_io_hit_2_3),
    .io_valid_2_3(Arbitration_2_2_io_valid_2_3),
    .io_ray_id_out(Arbitration_2_2_io_ray_id_out),
    .io_hit_out(Arbitration_2_2_io_hit_out),
    .io_valid_out(Arbitration_2_2_io_valid_out)
  );
  Arbitration_3 Arbitration_3 ( // @[Top_AO.scala 72:45]
    .clock(Arbitration_3_clock),
    .reset(Arbitration_3_reset),
    .io_node_id_3_0(Arbitration_3_io_node_id_3_0),
    .io_ray_id_3_0(Arbitration_3_io_ray_id_3_0),
    .io_hit_3_0(Arbitration_3_io_hit_3_0),
    .io_valid_3_0(Arbitration_3_io_valid_3_0),
    .io_node_id_3_1(Arbitration_3_io_node_id_3_1),
    .io_ray_id_3_1(Arbitration_3_io_ray_id_3_1),
    .io_hit_3_1(Arbitration_3_io_hit_3_1),
    .io_valid_3_1(Arbitration_3_io_valid_3_1),
    .io_node_id_3_2(Arbitration_3_io_node_id_3_2),
    .io_ray_id_3_2(Arbitration_3_io_ray_id_3_2),
    .io_hit_3_2(Arbitration_3_io_hit_3_2),
    .io_valid_3_2(Arbitration_3_io_valid_3_2),
    .io_node_id_3_3(Arbitration_3_io_node_id_3_3),
    .io_ray_id_3_3(Arbitration_3_io_ray_id_3_3),
    .io_hit_3_3(Arbitration_3_io_hit_3_3),
    .io_valid_3_3(Arbitration_3_io_valid_3_3),
    .io_node_id_3_4(Arbitration_3_io_node_id_3_4),
    .io_ray_id_3_4(Arbitration_3_io_ray_id_3_4),
    .io_hit_3_4(Arbitration_3_io_hit_3_4),
    .io_valid_3_4(Arbitration_3_io_valid_3_4),
    .io_node_id_out(Arbitration_3_io_node_id_out),
    .io_ray_id_out(Arbitration_3_io_ray_id_out),
    .io_hit_out(Arbitration_3_io_hit_out),
    .io_valid_out(Arbitration_3_io_valid_out)
  );
  Arbitration_3 Arbitration_3_2 ( // @[Top_AO.scala 73:42]
    .clock(Arbitration_3_2_clock),
    .reset(Arbitration_3_2_reset),
    .io_node_id_3_0(Arbitration_3_2_io_node_id_3_0),
    .io_ray_id_3_0(Arbitration_3_2_io_ray_id_3_0),
    .io_hit_3_0(Arbitration_3_2_io_hit_3_0),
    .io_valid_3_0(Arbitration_3_2_io_valid_3_0),
    .io_node_id_3_1(Arbitration_3_2_io_node_id_3_1),
    .io_ray_id_3_1(Arbitration_3_2_io_ray_id_3_1),
    .io_hit_3_1(Arbitration_3_2_io_hit_3_1),
    .io_valid_3_1(Arbitration_3_2_io_valid_3_1),
    .io_node_id_3_2(Arbitration_3_2_io_node_id_3_2),
    .io_ray_id_3_2(Arbitration_3_2_io_ray_id_3_2),
    .io_hit_3_2(Arbitration_3_2_io_hit_3_2),
    .io_valid_3_2(Arbitration_3_2_io_valid_3_2),
    .io_node_id_3_3(Arbitration_3_2_io_node_id_3_3),
    .io_ray_id_3_3(Arbitration_3_2_io_ray_id_3_3),
    .io_hit_3_3(Arbitration_3_2_io_hit_3_3),
    .io_valid_3_3(Arbitration_3_2_io_valid_3_3),
    .io_node_id_3_4(Arbitration_3_2_io_node_id_3_4),
    .io_ray_id_3_4(Arbitration_3_2_io_ray_id_3_4),
    .io_hit_3_4(Arbitration_3_2_io_hit_3_4),
    .io_valid_3_4(Arbitration_3_2_io_valid_3_4),
    .io_node_id_out(Arbitration_3_2_io_node_id_out),
    .io_ray_id_out(Arbitration_3_2_io_ray_id_out),
    .io_hit_out(Arbitration_3_2_io_hit_out),
    .io_valid_out(Arbitration_3_2_io_valid_out)
  );
  Arbitration_4 Arbitration_4 ( // @[Top_AO.scala 74:45]
    .clock(Arbitration_4_clock),
    .reset(Arbitration_4_reset),
    .io_node_id_4_0(Arbitration_4_io_node_id_4_0),
    .io_ray_id_4_0(Arbitration_4_io_ray_id_4_0),
    .io_hit_4_0(Arbitration_4_io_hit_4_0),
    .io_valid_4_0(Arbitration_4_io_valid_4_0),
    .io_node_id_4_1(Arbitration_4_io_node_id_4_1),
    .io_ray_id_4_1(Arbitration_4_io_ray_id_4_1),
    .io_hit_4_1(Arbitration_4_io_hit_4_1),
    .io_valid_4_1(Arbitration_4_io_valid_4_1),
    .io_node_id_out(Arbitration_4_io_node_id_out),
    .io_ray_id_out(Arbitration_4_io_ray_id_out),
    .io_hit_out(Arbitration_4_io_hit_out),
    .io_RAY_AABB_out(Arbitration_4_io_RAY_AABB_out),
    .io_RAY_AABB_2_out(Arbitration_4_io_RAY_AABB_2_out),
    .io_valid_out(Arbitration_4_io_valid_out)
  );
  Stackmanage Stack_manage ( // @[Top_AO.scala 76:41]
    .clock(Stack_manage_clock),
    .reset(Stack_manage_reset),
    .io_push(Stack_manage_io_push),
    .io_push_en(Stack_manage_io_push_en),
    .io_pop(Stack_manage_io_pop),
    .io_pop_en(Stack_manage_io_pop_en),
    .io_ray_id_push(Stack_manage_io_ray_id_push),
    .io_ray_id_pop(Stack_manage_io_ray_id_pop),
    .io_node_id_push_in(Stack_manage_io_node_id_push_in),
    .io_hitT_in(Stack_manage_io_hitT_in),
    .io_clear(Stack_manage_io_clear),
    .io_hitT_out(Stack_manage_io_hitT_out),
    .io_node_id_out(Stack_manage_io_node_id_out),
    .io_ray_id_out(Stack_manage_io_ray_id_out),
    .io_pop_valid(Stack_manage_io_pop_valid),
    .io_Dis_en(Stack_manage_io_Dis_en),
    .io_Finish(Stack_manage_io_Finish)
  );
  Stackmanage Stack_manage_2 ( // @[Top_AO.scala 77:38]
    .clock(Stack_manage_2_clock),
    .reset(Stack_manage_2_reset),
    .io_push(Stack_manage_2_io_push),
    .io_push_en(Stack_manage_2_io_push_en),
    .io_pop(Stack_manage_2_io_pop),
    .io_pop_en(Stack_manage_2_io_pop_en),
    .io_ray_id_push(Stack_manage_2_io_ray_id_push),
    .io_ray_id_pop(Stack_manage_2_io_ray_id_pop),
    .io_node_id_push_in(Stack_manage_2_io_node_id_push_in),
    .io_hitT_in(Stack_manage_2_io_hitT_in),
    .io_clear(Stack_manage_2_io_clear),
    .io_hitT_out(Stack_manage_2_io_hitT_out),
    .io_node_id_out(Stack_manage_2_io_node_id_out),
    .io_ray_id_out(Stack_manage_2_io_ray_id_out),
    .io_pop_valid(Stack_manage_2_io_pop_valid),
    .io_Dis_en(Stack_manage_2_io_Dis_en),
    .io_Finish(Stack_manage_2_io_Finish)
  );
  Triangle Triangle ( // @[Top_AO.scala 78:51]
    .clock(Triangle_clock),
    .reset(Triangle_reset),
    .io_To_IST0_enable(Triangle_io_To_IST0_enable),
    .io_nodeid_leaf(Triangle_io_nodeid_leaf),
    .io_rayid_leaf(Triangle_io_rayid_leaf),
    .io_hiT_in(Triangle_io_hiT_in),
    .io_v00_in_x(Triangle_io_v00_in_x),
    .io_v00_in_y(Triangle_io_v00_in_y),
    .io_v00_in_z(Triangle_io_v00_in_z),
    .io_v00_in_w(Triangle_io_v00_in_w),
    .io_v11_in_x(Triangle_io_v11_in_x),
    .io_v11_in_y(Triangle_io_v11_in_y),
    .io_v11_in_z(Triangle_io_v11_in_z),
    .io_v11_in_w(Triangle_io_v11_in_w),
    .io_v22_in_x(Triangle_io_v22_in_x),
    .io_v22_in_y(Triangle_io_v22_in_y),
    .io_v22_in_z(Triangle_io_v22_in_z),
    .io_v22_in_w(Triangle_io_v22_in_w),
    .io_ray_o_in_x(Triangle_io_ray_o_in_x),
    .io_ray_o_in_y(Triangle_io_ray_o_in_y),
    .io_ray_o_in_z(Triangle_io_ray_o_in_z),
    .io_ray_d_in_x(Triangle_io_ray_d_in_x),
    .io_ray_d_in_y(Triangle_io_ray_d_in_y),
    .io_ray_d_in_z(Triangle_io_ray_d_in_z),
    .io_break_in(Triangle_io_break_in),
    .io_RAY_AABB_1(Triangle_io_RAY_AABB_1),
    .io_RAY_AABB_2(Triangle_io_RAY_AABB_2),
    .io_pop_1(Triangle_io_pop_1),
    .io_break_1(Triangle_io_break_1),
    .io_pop_2(Triangle_io_pop_2),
    .io_break_2(Triangle_io_break_2),
    .io_pop_3(Triangle_io_pop_3),
    .io_break_3(Triangle_io_break_3),
    .io_hiT_out_1(Triangle_io_hiT_out_1),
    .io_hiT_out_2(Triangle_io_hiT_out_2),
    .io_hiT_out_3(Triangle_io_hiT_out_3),
    .io_hitT_en(Triangle_io_hitT_en),
    .io_hitIndex(Triangle_io_hitIndex),
    .io_hitIndex_en(Triangle_io_hitIndex_en),
    .io_node_id_out_1(Triangle_io_node_id_out_1),
    .io_node_id_out_2(Triangle_io_node_id_out_2),
    .io_node_id_out_3(Triangle_io_node_id_out_3),
    .io_ray_id_ist1(Triangle_io_ray_id_ist1),
    .io_ray_id_ist2(Triangle_io_ray_id_ist2),
    .io_ray_id_ist3(Triangle_io_ray_id_ist3),
    .io_counter_fdiv(Triangle_io_counter_fdiv),
    .io_RAY_AABB_1_out_IST1(Triangle_io_RAY_AABB_1_out_IST1),
    .io_RAY_AABB_2_out_IST1(Triangle_io_RAY_AABB_2_out_IST1),
    .io_RAY_AABB_1_out_IST2(Triangle_io_RAY_AABB_1_out_IST2),
    .io_RAY_AABB_2_out_IST2(Triangle_io_RAY_AABB_2_out_IST2),
    .io_RAY_AABB_1_out_IST3(Triangle_io_RAY_AABB_1_out_IST3),
    .io_RAY_AABB_2_out_IST3(Triangle_io_RAY_AABB_2_out_IST3)
  );
  assign io_hitT = Triangle_io_hitT_en ? Triangle_io_hiT_out_3 : 32'h0; // @[Top_AO.scala 770:30 Top_AO.scala 771:65 Top_AO.scala 775:65]
  assign io_hitIndex = Triangle_io_hitT_en ? $signed(Triangle_io_hitIndex) : $signed(32'sh0); // @[Top_AO.scala 770:30 Top_AO.scala 772:65 Top_AO.scala 776:65]
  assign io_rtp_finish = Ray_Dispatch_io_ray_finish & Stack_manage_io_Finish; // @[Top_AO.scala 113:87]
  assign io_ray_id_triangle = Triangle_io_hitT_en ? Triangle_io_ray_id_ist3 : 32'h0; // @[Top_AO.scala 770:30 Top_AO.scala 773:65 Top_AO.scala 777:65]
  assign io_counter_fdiv = Triangle_io_counter_fdiv; // @[Top_AO.scala 765:57]
  assign io_TRV_1_valid = TRV_1; // @[Top_AO.scala 256:61]
  assign io_TRV_2_valid = TRV_2; // @[Top_AO.scala 402:66]
  assign io_IST_1_valid = IST_1; // @[Top_AO.scala 759:59]
  assign io_clock_count = clock_counter; // @[Top_AO.scala 82:37]
  assign Ray_Dispatch_clock = clock;
  assign Ray_Dispatch_reset = reset;
  assign Ray_Dispatch_io_dispatch = Stack_manage_io_Dis_en | Triangle_io_hitIndex_en & Triangle_io_RAY_AABB_1_out_IST3; // @[Top_AO.scala 85:79]
  assign Ray_Dispatch_io_dispatch_2 = Stack_manage_2_io_Dis_en | Triangle_io_hitIndex_en &
    Triangle_io_RAY_AABB_2_out_IST3; // @[Top_AO.scala 86:81]
  assign Ray_origx_clock = clock;
  assign Ray_origx_io_Ray_id = Arbitration_4_io_ray_id_out; // @[Top_AO.scala 679:37 Top_AO.scala 685:54]
  assign Ray_origx_io_Ray_id_2 = 32'h0;
  assign Ray_origy_clock = clock;
  assign Ray_origy_io_Ray_id = Arbitration_4_io_ray_id_out; // @[Top_AO.scala 679:37 Top_AO.scala 685:54]
  assign Ray_origy_io_Ray_id_2 = 32'h0;
  assign Ray_origz_clock = clock;
  assign Ray_origz_io_Ray_id = Arbitration_4_io_ray_id_out; // @[Top_AO.scala 679:37 Top_AO.scala 685:54]
  assign Ray_origz_io_Ray_id_2 = 32'h0;
  assign Ray_dirx_clock = clock;
  assign Ray_dirx_io_Ray_id = Arbitration_4_io_ray_id_out; // @[Top_AO.scala 679:37 Top_AO.scala 685:54]
  assign Ray_dirx_io_Ray_id_2 = 32'h0;
  assign Ray_diry_clock = clock;
  assign Ray_diry_io_Ray_id = Arbitration_4_io_ray_id_out; // @[Top_AO.scala 679:37 Top_AO.scala 685:54]
  assign Ray_diry_io_Ray_id_2 = 32'h0;
  assign Ray_dirz_clock = clock;
  assign Ray_dirz_io_Ray_id = Arbitration_4_io_ray_id_out; // @[Top_AO.scala 679:37 Top_AO.scala 685:54]
  assign Ray_dirz_io_Ray_id_2 = 32'h0;
  assign Ray_hitT_clock = clock;
  assign Ray_hitT_io_Ray_id = Arbitration_1_io_hit_out; // @[Top_AO.scala 165:76 Top_AO.scala 188:53]
  assign Ray_hitT_io_Ray_id_2 = Arbitration_1_2_io_ray_id_out; // @[Top_AO.scala 302:80 Top_AO.scala 306:54]
  assign Ray_idirx_clock = clock;
  assign Ray_idirx_io_Ray_id = Arbitration_1_io_valid_out & Arbitration_1_io_hit_out != 32'h0 ?
    Arbitration_1_io_ray_id_out : _GEN_13; // @[Top_AO.scala 140:70 Top_AO.scala 142:51]
  assign Ray_idirx_io_Ray_id_2 = Arbitration_1_2_io_valid_out & Arbitration_1_2_io_hit_out != 32'h0 ?
    Arbitration_1_2_io_ray_id_out : _GEN_81; // @[Top_AO.scala 275:74 Top_AO.scala 279:55]
  assign Ray_idiry_clock = clock;
  assign Ray_idiry_io_Ray_id = Arbitration_1_io_valid_out & Arbitration_1_io_hit_out != 32'h0 ?
    Arbitration_1_io_ray_id_out : _GEN_13; // @[Top_AO.scala 140:70 Top_AO.scala 142:51]
  assign Ray_idiry_io_Ray_id_2 = Arbitration_1_2_io_valid_out & Arbitration_1_2_io_hit_out != 32'h0 ?
    Arbitration_1_2_io_ray_id_out : _GEN_81; // @[Top_AO.scala 275:74 Top_AO.scala 279:55]
  assign Ray_idirz_clock = clock;
  assign Ray_idirz_io_Ray_id = Arbitration_1_io_valid_out & Arbitration_1_io_hit_out != 32'h0 ?
    Arbitration_1_io_ray_id_out : _GEN_13; // @[Top_AO.scala 140:70 Top_AO.scala 142:51]
  assign Ray_idirz_io_Ray_id_2 = Arbitration_1_2_io_valid_out & Arbitration_1_2_io_hit_out != 32'h0 ?
    Arbitration_1_2_io_ray_id_out : _GEN_81; // @[Top_AO.scala 275:74 Top_AO.scala 279:55]
  assign Ray_oodx_clock = clock;
  assign Ray_oodx_io_Ray_id = Arbitration_1_io_valid_out & Arbitration_1_io_hit_out != 32'h0 ?
    Arbitration_1_io_ray_id_out : _GEN_13; // @[Top_AO.scala 140:70 Top_AO.scala 142:51]
  assign Ray_oodx_io_Ray_id_2 = Arbitration_1_2_io_valid_out & Arbitration_1_2_io_hit_out != 32'h0 ?
    Arbitration_1_2_io_ray_id_out : _GEN_81; // @[Top_AO.scala 275:74 Top_AO.scala 279:55]
  assign Ray_oody_clock = clock;
  assign Ray_oody_io_Ray_id = Arbitration_1_io_valid_out & Arbitration_1_io_hit_out != 32'h0 ?
    Arbitration_1_io_ray_id_out : _GEN_13; // @[Top_AO.scala 140:70 Top_AO.scala 142:51]
  assign Ray_oody_io_Ray_id_2 = Arbitration_1_2_io_valid_out & Arbitration_1_2_io_hit_out != 32'h0 ?
    Arbitration_1_2_io_ray_id_out : _GEN_81; // @[Top_AO.scala 275:74 Top_AO.scala 279:55]
  assign Ray_oodz_clock = clock;
  assign Ray_oodz_io_Ray_id = Arbitration_1_io_valid_out & Arbitration_1_io_hit_out != 32'h0 ?
    Arbitration_1_io_ray_id_out : _GEN_13; // @[Top_AO.scala 140:70 Top_AO.scala 142:51]
  assign Ray_oodz_io_Ray_id_2 = Arbitration_1_2_io_valid_out & Arbitration_1_2_io_hit_out != 32'h0 ?
    Arbitration_1_2_io_ray_id_out : _GEN_81; // @[Top_AO.scala 275:74 Top_AO.scala 279:55]
  assign BVH_RAM_0_x_clock = clock;
  assign BVH_RAM_0_x_io_BVH_id = _GEN_34[31:0];
  assign BVH_RAM_0_x_io_BVH_id_2 = _GEN_101[31:0];
  assign BVH_RAM_0_y_clock = clock;
  assign BVH_RAM_0_y_io_BVH_id = _GEN_34[31:0];
  assign BVH_RAM_0_y_io_BVH_id_2 = _GEN_101[31:0];
  assign BVH_RAM_0_z_clock = clock;
  assign BVH_RAM_0_z_io_BVH_id = _GEN_34[31:0];
  assign BVH_RAM_0_z_io_BVH_id_2 = _GEN_101[31:0];
  assign BVH_RAM_0_w_clock = clock;
  assign BVH_RAM_0_w_io_BVH_id = _GEN_34[31:0];
  assign BVH_RAM_0_w_io_BVH_id_2 = _GEN_101[31:0];
  assign BVH_RAM_1_x_clock = clock;
  assign BVH_RAM_1_x_io_BVH_id = _GEN_34[31:0];
  assign BVH_RAM_1_x_io_BVH_id_2 = _GEN_101[31:0];
  assign BVH_RAM_1_y_clock = clock;
  assign BVH_RAM_1_y_io_BVH_id = _GEN_34[31:0];
  assign BVH_RAM_1_y_io_BVH_id_2 = _GEN_101[31:0];
  assign BVH_RAM_1_z_clock = clock;
  assign BVH_RAM_1_z_io_BVH_id = _GEN_34[31:0];
  assign BVH_RAM_1_z_io_BVH_id_2 = _GEN_101[31:0];
  assign BVH_RAM_1_w_clock = clock;
  assign BVH_RAM_1_w_io_BVH_id = _GEN_34[31:0];
  assign BVH_RAM_1_w_io_BVH_id_2 = _GEN_101[31:0];
  assign BVH_RAM_z_x_clock = clock;
  assign BVH_RAM_z_x_io_BVH_id = _GEN_34[31:0];
  assign BVH_RAM_z_x_io_BVH_id_2 = _GEN_101[31:0];
  assign BVH_RAM_z_y_clock = clock;
  assign BVH_RAM_z_y_io_BVH_id = _GEN_34[31:0];
  assign BVH_RAM_z_y_io_BVH_id_2 = _GEN_101[31:0];
  assign BVH_RAM_z_z_clock = clock;
  assign BVH_RAM_z_z_io_BVH_id = _GEN_34[31:0];
  assign BVH_RAM_z_z_io_BVH_id_2 = _GEN_101[31:0];
  assign BVH_RAM_z_w_clock = clock;
  assign BVH_RAM_z_w_io_BVH_id = _GEN_34[31:0];
  assign BVH_RAM_z_w_io_BVH_id_2 = _GEN_101[31:0];
  assign BVH_RAM_tmp_x_clock = clock;
  assign BVH_RAM_tmp_x_io_BVH_id = _GEN_34[31:0];
  assign BVH_RAM_tmp_x_io_BVH_id_2 = _GEN_101[31:0];
  assign BVH_RAM_tmp_y_clock = clock;
  assign BVH_RAM_tmp_y_io_BVH_id = _GEN_34[31:0];
  assign BVH_RAM_tmp_y_io_BVH_id_2 = _GEN_101[31:0];
  assign TRI_RAM_x_clock = clock;
  assign TRI_RAM_x_io_Triangle_id = Arbitration_4_io_node_id_out; // @[Top_AO.scala 679:37 Top_AO.scala 681:47]
  assign TRI_RAM_y_clock = clock;
  assign TRI_RAM_y_io_Triangle_id = Arbitration_4_io_node_id_out; // @[Top_AO.scala 679:37 Top_AO.scala 681:47]
  assign TRI_RAM_z_clock = clock;
  assign TRI_RAM_z_io_Triangle_id = Arbitration_4_io_node_id_out; // @[Top_AO.scala 679:37 Top_AO.scala 681:47]
  assign TRI_RAM_w_clock = clock;
  assign TRI_RAM_w_io_Triangle_id = Arbitration_4_io_node_id_out; // @[Top_AO.scala 679:37 Top_AO.scala 681:47]
  assign RAY_AABB_clock = clock;
  assign RAY_AABB_reset = reset;
  assign RAY_AABB_io_ray_idir_x = memory_valid ? Ray_idirx_io_Ray_out : 32'h0; // @[Top_AO.scala 196:29 Top_AO.scala 197:53 Top_AO.scala 230:53]
  assign RAY_AABB_io_ray_idir_y = memory_valid ? Ray_idiry_io_Ray_out : 32'h0; // @[Top_AO.scala 196:29 Top_AO.scala 198:53 Top_AO.scala 231:53]
  assign RAY_AABB_io_ray_idir_z = memory_valid ? Ray_idirz_io_Ray_out : 32'h0; // @[Top_AO.scala 196:29 Top_AO.scala 199:53 Top_AO.scala 232:53]
  assign RAY_AABB_io_ray_ood_x = memory_valid ? Ray_oodx_io_Ray_out : 32'h0; // @[Top_AO.scala 196:29 Top_AO.scala 200:51 Top_AO.scala 233:51]
  assign RAY_AABB_io_ray_ood_y = memory_valid ? Ray_oody_io_Ray_out : 32'h0; // @[Top_AO.scala 196:29 Top_AO.scala 201:51 Top_AO.scala 234:51]
  assign RAY_AABB_io_ray_ood_z = memory_valid ? Ray_oodz_io_Ray_out : 32'h0; // @[Top_AO.scala 196:29 Top_AO.scala 202:51 Top_AO.scala 235:51]
  assign RAY_AABB_io_ray_hitT = memory_valid ? _GEN_51 : 32'h0; // @[Top_AO.scala 196:29 Top_AO.scala 236:53]
  assign RAY_AABB_io_bvh_n0xy_x = memory_valid ? BVH_RAM_0_x_io_BVH_out : 32'h0; // @[Top_AO.scala 196:29 Top_AO.scala 209:49 Top_AO.scala 238:49]
  assign RAY_AABB_io_bvh_n0xy_y = memory_valid ? BVH_RAM_0_y_io_BVH_out : 32'h0; // @[Top_AO.scala 196:29 Top_AO.scala 210:49 Top_AO.scala 239:49]
  assign RAY_AABB_io_bvh_n0xy_z = memory_valid ? BVH_RAM_0_z_io_BVH_out : 32'h0; // @[Top_AO.scala 196:29 Top_AO.scala 211:49 Top_AO.scala 240:49]
  assign RAY_AABB_io_bvh_n0xy_w = memory_valid ? BVH_RAM_0_w_io_BVH_out : 32'h0; // @[Top_AO.scala 196:29 Top_AO.scala 212:48 Top_AO.scala 241:48]
  assign RAY_AABB_io_bvh_n1xy_x = memory_valid ? BVH_RAM_1_x_io_BVH_out : 32'h0; // @[Top_AO.scala 196:29 Top_AO.scala 214:49 Top_AO.scala 242:49]
  assign RAY_AABB_io_bvh_n1xy_y = memory_valid ? BVH_RAM_1_y_io_BVH_out : 32'h0; // @[Top_AO.scala 196:29 Top_AO.scala 215:49 Top_AO.scala 243:49]
  assign RAY_AABB_io_bvh_n1xy_z = memory_valid ? BVH_RAM_1_z_io_BVH_out : 32'h0; // @[Top_AO.scala 196:29 Top_AO.scala 216:49 Top_AO.scala 244:49]
  assign RAY_AABB_io_bvh_n1xy_w = memory_valid ? BVH_RAM_1_w_io_BVH_out : 32'h0; // @[Top_AO.scala 196:29 Top_AO.scala 217:48 Top_AO.scala 245:48]
  assign RAY_AABB_io_bvh_nz_x = memory_valid ? BVH_RAM_z_x_io_BVH_out : 32'h0; // @[Top_AO.scala 196:29 Top_AO.scala 219:51 Top_AO.scala 246:51]
  assign RAY_AABB_io_bvh_nz_y = memory_valid ? BVH_RAM_z_y_io_BVH_out : 32'h0; // @[Top_AO.scala 196:29 Top_AO.scala 220:51 Top_AO.scala 247:51]
  assign RAY_AABB_io_bvh_nz_z = memory_valid ? BVH_RAM_z_z_io_BVH_out : 32'h0; // @[Top_AO.scala 196:29 Top_AO.scala 221:51 Top_AO.scala 248:51]
  assign RAY_AABB_io_bvh_nz_w = memory_valid ? BVH_RAM_z_w_io_BVH_out : 32'h0; // @[Top_AO.scala 196:29 Top_AO.scala 222:50 Top_AO.scala 249:49]
  assign RAY_AABB_io_bvh_temp_x = memory_valid ? $signed(BVH_RAM_tmp_x_io_BVH_out) : $signed(32'sh0); // @[Top_AO.scala 196:29 Top_AO.scala 224:48 Top_AO.scala 250:48]
  assign RAY_AABB_io_bvh_temp_y = memory_valid ? $signed(BVH_RAM_tmp_y_io_BVH_out) : $signed(32'sh0); // @[Top_AO.scala 196:29 Top_AO.scala 225:48 Top_AO.scala 251:48]
  assign RAY_AABB_io_rayid = memory_valid ? ray_id_temp : 32'h0; // @[Top_AO.scala 196:29 Top_AO.scala 226:57 Top_AO.scala 252:57]
  assign RAY_AABB_io_valid_en = memory_valid; // @[Top_AO.scala 196:29 Top_AO.scala 227:53 Top_AO.scala 253:53]
  assign RAY_AABB_2_clock = clock;
  assign RAY_AABB_2_reset = reset;
  assign RAY_AABB_2_io_ray_idir_x = memory_valid_2 ? Ray_idirx_io_Ray_out_2 : 32'h0; // @[Top_AO.scala 335:31 Top_AO.scala 336:55 Top_AO.scala 366:55]
  assign RAY_AABB_2_io_ray_idir_y = memory_valid_2 ? Ray_idiry_io_Ray_out_2 : 32'h0; // @[Top_AO.scala 335:31 Top_AO.scala 337:55 Top_AO.scala 367:55]
  assign RAY_AABB_2_io_ray_idir_z = memory_valid_2 ? Ray_idirz_io_Ray_out_2 : 32'h0; // @[Top_AO.scala 335:31 Top_AO.scala 338:55 Top_AO.scala 368:55]
  assign RAY_AABB_2_io_ray_ood_x = memory_valid_2 ? Ray_oodx_io_Ray_out_2 : 32'h0; // @[Top_AO.scala 335:31 Top_AO.scala 339:53 Top_AO.scala 369:53]
  assign RAY_AABB_2_io_ray_ood_y = memory_valid_2 ? Ray_oody_io_Ray_out_2 : 32'h0; // @[Top_AO.scala 335:31 Top_AO.scala 340:53 Top_AO.scala 370:53]
  assign RAY_AABB_2_io_ray_ood_z = memory_valid_2 ? Ray_oodz_io_Ray_out_2 : 32'h0; // @[Top_AO.scala 335:31 Top_AO.scala 341:53 Top_AO.scala 371:53]
  assign RAY_AABB_2_io_ray_hitT = memory_valid_2 ? _GEN_118 : 32'h0; // @[Top_AO.scala 335:31 Top_AO.scala 372:55]
  assign RAY_AABB_2_io_bvh_n0xy_x = memory_valid_2 ? BVH_RAM_0_x_io_BVH_out_2 : 32'h0; // @[Top_AO.scala 335:31 Top_AO.scala 348:51 Top_AO.scala 374:51]
  assign RAY_AABB_2_io_bvh_n0xy_y = memory_valid_2 ? BVH_RAM_0_y_io_BVH_out_2 : 32'h0; // @[Top_AO.scala 335:31 Top_AO.scala 349:51 Top_AO.scala 375:51]
  assign RAY_AABB_2_io_bvh_n0xy_z = memory_valid_2 ? BVH_RAM_0_z_io_BVH_out_2 : 32'h0; // @[Top_AO.scala 335:31 Top_AO.scala 350:51 Top_AO.scala 376:51]
  assign RAY_AABB_2_io_bvh_n0xy_w = memory_valid_2 ? BVH_RAM_0_w_io_BVH_out_2 : 32'h0; // @[Top_AO.scala 335:31 Top_AO.scala 351:50 Top_AO.scala 377:50]
  assign RAY_AABB_2_io_bvh_n1xy_x = memory_valid_2 ? BVH_RAM_1_x_io_BVH_out_2 : 32'h0; // @[Top_AO.scala 335:31 Top_AO.scala 352:51 Top_AO.scala 378:51]
  assign RAY_AABB_2_io_bvh_n1xy_y = memory_valid_2 ? BVH_RAM_1_y_io_BVH_out_2 : 32'h0; // @[Top_AO.scala 335:31 Top_AO.scala 353:51 Top_AO.scala 379:51]
  assign RAY_AABB_2_io_bvh_n1xy_z = memory_valid_2 ? BVH_RAM_1_z_io_BVH_out_2 : 32'h0; // @[Top_AO.scala 335:31 Top_AO.scala 354:51 Top_AO.scala 380:51]
  assign RAY_AABB_2_io_bvh_n1xy_w = memory_valid_2 ? BVH_RAM_1_w_io_BVH_out_2 : 32'h0; // @[Top_AO.scala 335:31 Top_AO.scala 355:50 Top_AO.scala 381:50]
  assign RAY_AABB_2_io_bvh_nz_x = memory_valid_2 ? BVH_RAM_z_x_io_BVH_out_2 : 32'h0; // @[Top_AO.scala 335:31 Top_AO.scala 356:53 Top_AO.scala 382:53]
  assign RAY_AABB_2_io_bvh_nz_y = memory_valid_2 ? BVH_RAM_z_y_io_BVH_out_2 : 32'h0; // @[Top_AO.scala 335:31 Top_AO.scala 357:53 Top_AO.scala 383:53]
  assign RAY_AABB_2_io_bvh_nz_z = memory_valid_2 ? BVH_RAM_z_z_io_BVH_out_2 : 32'h0; // @[Top_AO.scala 335:31 Top_AO.scala 358:53 Top_AO.scala 384:53]
  assign RAY_AABB_2_io_bvh_nz_w = memory_valid_2 ? BVH_RAM_z_w_io_BVH_out_2 : 32'h0; // @[Top_AO.scala 335:31 Top_AO.scala 359:52 Top_AO.scala 385:51]
  assign RAY_AABB_2_io_bvh_temp_x = memory_valid_2 ? $signed(BVH_RAM_tmp_x_io_BVH_out_2) : $signed(32'sh0); // @[Top_AO.scala 335:31 Top_AO.scala 360:50 Top_AO.scala 387:50]
  assign RAY_AABB_2_io_bvh_temp_y = memory_valid_2 ? $signed(BVH_RAM_tmp_y_io_BVH_out_2) : $signed(32'sh0); // @[Top_AO.scala 335:31 Top_AO.scala 361:50 Top_AO.scala 388:50]
  assign RAY_AABB_2_io_rayid = memory_valid_2 ? ray_id_temp_2 : 32'h0; // @[Top_AO.scala 335:31 Top_AO.scala 362:59 Top_AO.scala 389:59]
  assign RAY_AABB_2_io_valid_en = memory_valid_2; // @[Top_AO.scala 335:31 Top_AO.scala 363:55 Top_AO.scala 390:55]
  assign Arbitration_1_clock = clock;
  assign Arbitration_1_reset = reset;
  assign Arbitration_1_io_node_id_0 = _T_102 & Stack_manage_io_pop_valid ? $signed(Stack_manage_io_node_id_out) :
    $signed(32'sh0); // @[Top_AO.scala 457:81 Top_AO.scala 458:47]
  assign Arbitration_1_io_ray_id_0 = {{32'd0}, _GEN_168}; // @[Top_AO.scala 457:81 Top_AO.scala 459:50]
  assign Arbitration_1_io_hit_0 = _T_102 & Stack_manage_io_pop_valid ? Stack_manage_io_hitT_out : 32'h0; // @[Top_AO.scala 457:81 Top_AO.scala 460:54]
  assign Arbitration_1_io_valid_0 = _T_102 & Stack_manage_io_pop_valid; // @[Top_AO.scala 457:53]
  assign Arbitration_1_io_node_id_1 = RAY_AABB_io_back & RAY_AABB_io_valid_out ? $signed(RAY_AABB_io_nodeIdx_1) :
    $signed(32'sh0); // @[Top_AO.scala 116:50 Top_AO.scala 117:37 Top_AO.scala 121:37]
  assign Arbitration_1_io_ray_id_1 = RAY_AABB_io_back & RAY_AABB_io_valid_out ? RAY_AABB_io_rayid_out : 32'h0; // @[Top_AO.scala 116:50 Top_AO.scala 118:40 Top_AO.scala 122:40]
  assign Arbitration_1_io_valid_1 = RAY_AABB_io_back & RAY_AABB_io_valid_out & RAY_AABB_io_back; // @[Top_AO.scala 116:50 Top_AO.scala 119:42 Top_AO.scala 123:42]
  assign Arbitration_1_io_ray_id_2 = Ray_Dispatch_io_ray_out ? Ray_Dispatch_io_rayid_id : 32'h0; // @[Top_AO.scala 93:43 Top_AO.scala 95:56 Top_AO.scala 99:56]
  assign Arbitration_1_io_valid_2 = Ray_Dispatch_io_ray_out; // @[Top_AO.scala 93:33]
  assign Arbitration_1_2_clock = clock;
  assign Arbitration_1_2_reset = reset;
  assign Arbitration_1_2_io_node_id_0 = _T_117 & Stack_manage_2_io_pop_valid ? $signed(Stack_manage_2_io_node_id_out) :
    $signed(32'sh0); // @[Top_AO.scala 477:85 Top_AO.scala 478:49]
  assign Arbitration_1_2_io_ray_id_0 = {{32'd0}, _GEN_182}; // @[Top_AO.scala 477:85 Top_AO.scala 479:52]
  assign Arbitration_1_2_io_hit_0 = _T_117 & Stack_manage_2_io_pop_valid ? Stack_manage_2_io_hitT_out : 32'h0; // @[Top_AO.scala 477:85 Top_AO.scala 480:56]
  assign Arbitration_1_2_io_valid_0 = _T_117 & Stack_manage_2_io_pop_valid; // @[Top_AO.scala 477:55]
  assign Arbitration_1_2_io_node_id_1 = RAY_AABB_2_io_back & RAY_AABB_2_io_valid_out ? $signed(RAY_AABB_2_io_nodeIdx_1)
     : $signed(32'sh0); // @[Top_AO.scala 125:54 Top_AO.scala 126:39 Top_AO.scala 130:39]
  assign Arbitration_1_2_io_ray_id_1 = RAY_AABB_2_io_back & RAY_AABB_2_io_valid_out ? RAY_AABB_2_io_rayid_out : 32'h0; // @[Top_AO.scala 125:54 Top_AO.scala 127:42 Top_AO.scala 131:42]
  assign Arbitration_1_2_io_valid_1 = RAY_AABB_2_io_back & RAY_AABB_2_io_valid_out & RAY_AABB_2_io_back; // @[Top_AO.scala 125:54 Top_AO.scala 128:44 Top_AO.scala 132:44]
  assign Arbitration_1_2_io_ray_id_2 = Ray_Dispatch_io_ray_out_2 ? Ray_Dispatch_io_rayid_id_2 : 32'h0; // @[Top_AO.scala 103:45 Top_AO.scala 105:58 Top_AO.scala 109:58]
  assign Arbitration_1_2_io_valid_2 = Ray_Dispatch_io_ray_out_2; // @[Top_AO.scala 103:35]
  assign Arbitration_2_clock = clock;
  assign Arbitration_2_reset = reset;
  assign Arbitration_2_io_ray_id_2_0 = Triangle_io_break_3 & Triangle_io_RAY_AABB_1_out_IST3 ? Triangle_io_ray_id_ist3
     : 32'h0; // @[Top_AO.scala 645:63 Top_AO.scala 647:46 Top_AO.scala 652:46]
  assign Arbitration_2_io_hit_2_0 = Triangle_io_break_3 & Triangle_io_RAY_AABB_1_out_IST3 ? Triangle_io_hiT_out_3 : 32'h0
    ; // @[Top_AO.scala 645:63 Top_AO.scala 648:50 Top_AO.scala 653:50]
  assign Arbitration_2_io_valid_2_0 = Triangle_io_break_3 & Triangle_io_RAY_AABB_1_out_IST3; // @[Top_AO.scala 645:29]
  assign Arbitration_2_io_ray_id_2_1 = Triangle_io_break_2 & Triangle_io_RAY_AABB_1_out_IST2 ? Triangle_io_ray_id_ist2
     : 32'h0; // @[Top_AO.scala 621:63 Top_AO.scala 623:46 Top_AO.scala 628:46]
  assign Arbitration_2_io_hit_2_1 = Triangle_io_break_2 & Triangle_io_RAY_AABB_1_out_IST2 ? Triangle_io_hiT_out_2 : 32'h0
    ; // @[Top_AO.scala 621:63 Top_AO.scala 624:50 Top_AO.scala 629:50]
  assign Arbitration_2_io_valid_2_1 = Triangle_io_break_2 & Triangle_io_RAY_AABB_1_out_IST2; // @[Top_AO.scala 621:29]
  assign Arbitration_2_io_ray_id_2_2 = Triangle_io_break_1 & Triangle_io_RAY_AABB_1_out_IST1 ? Triangle_io_ray_id_ist1
     : 32'h0; // @[Top_AO.scala 596:63 Top_AO.scala 598:46 Top_AO.scala 603:46]
  assign Arbitration_2_io_hit_2_2 = Triangle_io_break_1 & Triangle_io_RAY_AABB_1_out_IST1 ? Triangle_io_hiT_out_1 : 32'h0
    ; // @[Top_AO.scala 596:63 Top_AO.scala 599:50 Top_AO.scala 604:50]
  assign Arbitration_2_io_valid_2_2 = Triangle_io_break_1 & Triangle_io_RAY_AABB_1_out_IST1; // @[Top_AO.scala 596:29]
  assign Arbitration_2_io_ray_id_2_3 = RAY_AABB_io_pop & RAY_AABB_io_valid_out ? RAY_AABB_io_rayid_out : 32'h0; // @[Top_AO.scala 257:49 Top_AO.scala 259:48 Top_AO.scala 264:48]
  assign Arbitration_2_io_hit_2_3 = RAY_AABB_io_pop & RAY_AABB_io_valid_out ? RAY_AABB_io_hitT_out : 32'h0; // @[Top_AO.scala 257:49 Top_AO.scala 260:52 Top_AO.scala 265:52]
  assign Arbitration_2_io_valid_2_3 = RAY_AABB_io_pop & RAY_AABB_io_valid_out; // @[Top_AO.scala 257:25]
  assign Arbitration_2_2_clock = clock;
  assign Arbitration_2_2_reset = reset;
  assign Arbitration_2_2_io_ray_id_2_0 = Triangle_io_break_3 & Triangle_io_RAY_AABB_2_out_IST3 ? Triangle_io_ray_id_ist3
     : 32'h0; // @[Top_AO.scala 657:60 Top_AO.scala 659:48 Top_AO.scala 664:48]
  assign Arbitration_2_2_io_hit_2_0 = Triangle_io_break_3 & Triangle_io_RAY_AABB_2_out_IST3 ? Triangle_io_hiT_out_3 : 32'h0
    ; // @[Top_AO.scala 657:60 Top_AO.scala 660:52 Top_AO.scala 665:52]
  assign Arbitration_2_2_io_valid_2_0 = Triangle_io_break_3 & Triangle_io_RAY_AABB_2_out_IST3; // @[Top_AO.scala 657:26]
  assign Arbitration_2_2_io_ray_id_2_1 = Triangle_io_break_2 & Triangle_io_RAY_AABB_2_out_IST2 ? Triangle_io_ray_id_ist2
     : 32'h0; // @[Top_AO.scala 632:63 Top_AO.scala 634:48 Top_AO.scala 639:48]
  assign Arbitration_2_2_io_hit_2_1 = Triangle_io_break_2 & Triangle_io_RAY_AABB_2_out_IST2 ? Triangle_io_hiT_out_2 : 32'h0
    ; // @[Top_AO.scala 632:63 Top_AO.scala 635:52 Top_AO.scala 640:52]
  assign Arbitration_2_2_io_valid_2_1 = Triangle_io_break_2 & Triangle_io_RAY_AABB_2_out_IST2; // @[Top_AO.scala 632:29]
  assign Arbitration_2_2_io_ray_id_2_2 = Triangle_io_break_1 & Triangle_io_RAY_AABB_2_out_IST1 ? Triangle_io_ray_id_ist1
     : 32'h0; // @[Top_AO.scala 608:63 Top_AO.scala 610:48 Top_AO.scala 615:48]
  assign Arbitration_2_2_io_hit_2_2 = Triangle_io_break_1 & Triangle_io_RAY_AABB_2_out_IST1 ? Triangle_io_hiT_out_1 : 32'h0
    ; // @[Top_AO.scala 608:63 Top_AO.scala 611:52 Top_AO.scala 616:52]
  assign Arbitration_2_2_io_valid_2_2 = Triangle_io_break_1 & Triangle_io_RAY_AABB_2_out_IST1; // @[Top_AO.scala 608:29]
  assign Arbitration_2_2_io_ray_id_2_3 = RAY_AABB_2_io_pop & RAY_AABB_2_io_valid_out ? RAY_AABB_2_io_rayid_out : 32'h0; // @[Top_AO.scala 393:53 Top_AO.scala 394:50 Top_AO.scala 398:50]
  assign Arbitration_2_2_io_hit_2_3 = RAY_AABB_2_io_pop & RAY_AABB_2_io_valid_out ? RAY_AABB_2_io_hitT_out : 32'h0; // @[Top_AO.scala 393:53 Top_AO.scala 395:54 Top_AO.scala 399:54]
  assign Arbitration_2_2_io_valid_2_3 = RAY_AABB_2_io_pop & RAY_AABB_2_io_valid_out; // @[Top_AO.scala 393:27]
  assign Arbitration_3_clock = clock;
  assign Arbitration_3_reset = reset;
  assign Arbitration_3_io_node_id_3_0 = Triangle_io_pop_3 & Triangle_io_RAY_AABB_1_out_IST3 ? $signed(_T_150) : $signed(32'sh0
    ); // @[Top_AO.scala 571:62 Top_AO.scala 572:43 Top_AO.scala 577:43]
  assign Arbitration_3_io_ray_id_3_0 = Triangle_io_pop_3 & Triangle_io_RAY_AABB_1_out_IST3 ? Triangle_io_ray_id_ist3 : 32'h0
    ; // @[Top_AO.scala 571:62 Top_AO.scala 573:46 Top_AO.scala 578:46]
  assign Arbitration_3_io_hit_3_0 = Triangle_io_pop_3 & Triangle_io_RAY_AABB_1_out_IST3 ? Triangle_io_hiT_out_3 : 32'h0; // @[Top_AO.scala 571:62 Top_AO.scala 574:50 Top_AO.scala 579:50]
  assign Arbitration_3_io_valid_3_0 = Triangle_io_pop_3 & Triangle_io_RAY_AABB_1_out_IST3; // @[Top_AO.scala 571:28]
  assign Arbitration_3_io_node_id_3_1 = Triangle_io_pop_2 & Triangle_io_RAY_AABB_1_out_IST2 ? $signed(_T_142) : $signed(32'sh0
    ); // @[Top_AO.scala 547:61 Top_AO.scala 548:43 Top_AO.scala 553:43]
  assign Arbitration_3_io_ray_id_3_1 = Triangle_io_pop_2 & Triangle_io_RAY_AABB_1_out_IST2 ? Triangle_io_ray_id_ist2 : 32'h0
    ; // @[Top_AO.scala 547:61 Top_AO.scala 549:46 Top_AO.scala 554:46]
  assign Arbitration_3_io_hit_3_1 = Triangle_io_pop_2 & Triangle_io_RAY_AABB_1_out_IST2 ? Triangle_io_hiT_out_2 : 32'h0; // @[Top_AO.scala 547:61 Top_AO.scala 550:50 Top_AO.scala 555:50]
  assign Arbitration_3_io_valid_3_1 = Triangle_io_pop_2 & Triangle_io_RAY_AABB_1_out_IST2; // @[Top_AO.scala 547:27]
  assign Arbitration_3_io_node_id_3_2 = Triangle_io_pop_1 & Triangle_io_RAY_AABB_1_out_IST1 ? $signed(_T_134) : $signed(32'sh0
    ); // @[Top_AO.scala 522:59 Top_AO.scala 523:43 Top_AO.scala 528:43]
  assign Arbitration_3_io_ray_id_3_2 = Triangle_io_pop_1 & Triangle_io_RAY_AABB_1_out_IST1 ? Triangle_io_ray_id_ist1 : 32'h0
    ; // @[Top_AO.scala 522:59 Top_AO.scala 524:46 Top_AO.scala 529:46]
  assign Arbitration_3_io_hit_3_2 = Triangle_io_pop_1 & Triangle_io_RAY_AABB_1_out_IST1 ? Triangle_io_hiT_out_1 : 32'h0; // @[Top_AO.scala 522:59 Top_AO.scala 525:50 Top_AO.scala 530:50]
  assign Arbitration_3_io_valid_3_2 = Triangle_io_pop_1 & Triangle_io_RAY_AABB_1_out_IST1; // @[Top_AO.scala 522:25]
  assign Arbitration_3_io_node_id_3_3 = ~_T_102 & Stack_manage_io_pop_valid ? $signed(_T_115) : $signed(32'sh0); // @[Top_AO.scala 462:87 Top_AO.scala 463:44 Top_AO.scala 472:44]
  assign Arbitration_3_io_ray_id_3_3 = ~_T_102 & Stack_manage_io_pop_valid ? Stack_manage_io_ray_id_out : 32'h0; // @[Top_AO.scala 462:87 Top_AO.scala 464:47 Top_AO.scala 473:47]
  assign Arbitration_3_io_hit_3_3 = ~_T_102 & Stack_manage_io_pop_valid ? Stack_manage_io_hitT_out : 32'h0; // @[Top_AO.scala 462:87 Top_AO.scala 465:52 Top_AO.scala 474:52]
  assign Arbitration_3_io_valid_3_3 = ~_T_102 & Stack_manage_io_pop_valid; // @[Top_AO.scala 462:59]
  assign Arbitration_3_io_node_id_3_4 = RAY_AABB_io_leaf & RAY_AABB_io_valid_out ? $signed(_T_94) : $signed(32'sh0); // @[Top_AO.scala 432:50 Top_AO.scala 433:45 Top_AO.scala 438:45]
  assign Arbitration_3_io_ray_id_3_4 = RAY_AABB_io_leaf & RAY_AABB_io_valid_out ? RAY_AABB_io_rayid_out : 32'h0; // @[Top_AO.scala 432:50 Top_AO.scala 434:48 Top_AO.scala 439:48]
  assign Arbitration_3_io_hit_3_4 = RAY_AABB_io_leaf & RAY_AABB_io_valid_out ? RAY_AABB_io_hitT_out : 32'h0; // @[Top_AO.scala 432:50 Top_AO.scala 435:52 Top_AO.scala 440:52]
  assign Arbitration_3_io_valid_3_4 = RAY_AABB_io_leaf & RAY_AABB_io_valid_out; // @[Top_AO.scala 432:26]
  assign Arbitration_3_2_clock = clock;
  assign Arbitration_3_2_reset = reset;
  assign Arbitration_3_2_io_node_id_3_0 = Triangle_io_pop_3 & Triangle_io_RAY_AABB_2_out_IST3 ? $signed(_T_150) :
    $signed(32'sh0); // @[Top_AO.scala 582:61 Top_AO.scala 583:45 Top_AO.scala 588:45]
  assign Arbitration_3_2_io_ray_id_3_0 = Triangle_io_pop_3 & Triangle_io_RAY_AABB_2_out_IST3 ? Triangle_io_ray_id_ist3
     : 32'h0; // @[Top_AO.scala 582:61 Top_AO.scala 584:48 Top_AO.scala 589:48]
  assign Arbitration_3_2_io_hit_3_0 = Triangle_io_pop_3 & Triangle_io_RAY_AABB_2_out_IST3 ? Triangle_io_hiT_out_3 : 32'h0
    ; // @[Top_AO.scala 582:61 Top_AO.scala 585:52 Top_AO.scala 590:52]
  assign Arbitration_3_2_io_valid_3_0 = Triangle_io_pop_3 & Triangle_io_RAY_AABB_2_out_IST3; // @[Top_AO.scala 582:27]
  assign Arbitration_3_2_io_node_id_3_1 = Triangle_io_pop_2 & Triangle_io_RAY_AABB_2_out_IST2 ? $signed(_T_142) :
    $signed(32'sh0); // @[Top_AO.scala 558:61 Top_AO.scala 559:45 Top_AO.scala 564:45]
  assign Arbitration_3_2_io_ray_id_3_1 = Triangle_io_pop_2 & Triangle_io_RAY_AABB_2_out_IST2 ? Triangle_io_ray_id_ist2
     : 32'h0; // @[Top_AO.scala 558:61 Top_AO.scala 560:48 Top_AO.scala 565:48]
  assign Arbitration_3_2_io_hit_3_1 = Triangle_io_pop_2 & Triangle_io_RAY_AABB_2_out_IST2 ? Triangle_io_hiT_out_2 : 32'h0
    ; // @[Top_AO.scala 558:61 Top_AO.scala 561:52 Top_AO.scala 566:52]
  assign Arbitration_3_2_io_valid_3_1 = Triangle_io_pop_2 & Triangle_io_RAY_AABB_2_out_IST2; // @[Top_AO.scala 558:27]
  assign Arbitration_3_2_io_node_id_3_2 = Triangle_io_pop_1 & Triangle_io_RAY_AABB_2_out_IST1 ? $signed(_T_134) :
    $signed(32'sh0); // @[Top_AO.scala 534:61 Top_AO.scala 535:45 Top_AO.scala 540:45]
  assign Arbitration_3_2_io_ray_id_3_2 = Triangle_io_pop_1 & Triangle_io_RAY_AABB_2_out_IST1 ? Triangle_io_ray_id_ist1
     : 32'h0; // @[Top_AO.scala 534:61 Top_AO.scala 536:48 Top_AO.scala 541:48]
  assign Arbitration_3_2_io_hit_3_2 = Triangle_io_pop_1 & Triangle_io_RAY_AABB_2_out_IST1 ? Triangle_io_hiT_out_1 : 32'h0
    ; // @[Top_AO.scala 534:61 Top_AO.scala 537:52 Top_AO.scala 542:52]
  assign Arbitration_3_2_io_valid_3_2 = Triangle_io_pop_1 & Triangle_io_RAY_AABB_2_out_IST1; // @[Top_AO.scala 534:27]
  assign Arbitration_3_2_io_node_id_3_3 = ~_T_117 & Stack_manage_2_io_pop_valid ? $signed(_T_130) : $signed(32'sh0); // @[Top_AO.scala 482:91 Top_AO.scala 483:46 Top_AO.scala 492:46]
  assign Arbitration_3_2_io_ray_id_3_3 = ~_T_117 & Stack_manage_2_io_pop_valid ? Stack_manage_2_io_ray_id_out : 32'h0; // @[Top_AO.scala 482:91 Top_AO.scala 484:49 Top_AO.scala 493:49]
  assign Arbitration_3_2_io_hit_3_3 = ~_T_117 & Stack_manage_2_io_pop_valid ? Stack_manage_2_io_hitT_out : 32'h0; // @[Top_AO.scala 482:91 Top_AO.scala 485:54 Top_AO.scala 494:54]
  assign Arbitration_3_2_io_valid_3_3 = ~_T_117 & Stack_manage_2_io_pop_valid; // @[Top_AO.scala 482:61]
  assign Arbitration_3_2_io_node_id_3_4 = RAY_AABB_2_io_leaf & RAY_AABB_2_io_valid_out ? $signed(_T_100) : $signed(32'sh0
    ); // @[Top_AO.scala 443:54 Top_AO.scala 444:47 Top_AO.scala 449:47]
  assign Arbitration_3_2_io_ray_id_3_4 = RAY_AABB_2_io_leaf & RAY_AABB_2_io_valid_out ? RAY_AABB_2_io_rayid_out : 32'h0; // @[Top_AO.scala 443:54 Top_AO.scala 445:50 Top_AO.scala 450:50]
  assign Arbitration_3_2_io_hit_3_4 = RAY_AABB_2_io_leaf & RAY_AABB_2_io_valid_out ? RAY_AABB_2_io_hitT_out : 32'h0; // @[Top_AO.scala 443:54 Top_AO.scala 446:54 Top_AO.scala 451:54]
  assign Arbitration_3_2_io_valid_3_4 = RAY_AABB_2_io_leaf & RAY_AABB_2_io_valid_out; // @[Top_AO.scala 443:28]
  assign Arbitration_4_clock = clock;
  assign Arbitration_4_reset = reset;
  assign Arbitration_4_io_node_id_4_0 = Arbitration_3_io_valid_out ? $signed(Arbitration_3_io_node_id_out) : $signed(32'sh0
    ); // @[Top_AO.scala 498:37 Top_AO.scala 499:43 Top_AO.scala 504:43]
  assign Arbitration_4_io_ray_id_4_0 = Arbitration_3_io_valid_out ? Arbitration_3_io_ray_id_out : 32'h0; // @[Top_AO.scala 498:37 Top_AO.scala 500:46 Top_AO.scala 505:46]
  assign Arbitration_4_io_hit_4_0 = Arbitration_3_io_valid_out ? Arbitration_3_io_hit_out : 32'h0; // @[Top_AO.scala 498:37 Top_AO.scala 501:50 Top_AO.scala 506:50]
  assign Arbitration_4_io_valid_4_0 = Arbitration_3_io_valid_out; // @[Top_AO.scala 498:37 Top_AO.scala 502:47 Top_AO.scala 507:48]
  assign Arbitration_4_io_node_id_4_1 = Arbitration_3_2_io_valid_out ? $signed(Arbitration_3_2_io_node_id_out) :
    $signed(32'sh0); // @[Top_AO.scala 510:39 Top_AO.scala 511:43 Top_AO.scala 516:43]
  assign Arbitration_4_io_ray_id_4_1 = Arbitration_3_2_io_valid_out ? Arbitration_3_2_io_ray_id_out : 32'h0; // @[Top_AO.scala 510:39 Top_AO.scala 512:46 Top_AO.scala 517:46]
  assign Arbitration_4_io_hit_4_1 = Arbitration_3_2_io_valid_out ? Arbitration_3_2_io_hit_out : 32'h0; // @[Top_AO.scala 510:39 Top_AO.scala 513:50 Top_AO.scala 518:50]
  assign Arbitration_4_io_valid_4_1 = Arbitration_3_2_io_valid_out; // @[Top_AO.scala 510:39 Top_AO.scala 514:47 Top_AO.scala 519:47]
  assign Stack_manage_clock = clock;
  assign Stack_manage_reset = reset;
  assign Stack_manage_io_push = RAY_AABB_io_push & RAY_AABB_io_valid_out; // @[Top_AO.scala 407:26]
  assign Stack_manage_io_push_en = RAY_AABB_io_push & RAY_AABB_io_valid_out; // @[Top_AO.scala 407:26]
  assign Stack_manage_io_pop = Arbitration_2_io_valid_out; // @[Top_AO.scala 761:46]
  assign Stack_manage_io_pop_en = Arbitration_2_io_valid_out; // @[Top_AO.scala 762:42]
  assign Stack_manage_io_ray_id_push = RAY_AABB_io_push & RAY_AABB_io_valid_out ? RAY_AABB_io_rayid_out : 32'h0; // @[Top_AO.scala 407:50 Top_AO.scala 411:52 Top_AO.scala 416:53]
  assign Stack_manage_io_ray_id_pop = Arbitration_2_io_ray_id_out; // @[Top_AO.scala 763:38]
  assign Stack_manage_io_node_id_push_in = RAY_AABB_io_push & RAY_AABB_io_valid_out ? $signed(RAY_AABB_io_nodeIdx_0) :
    $signed(32'sh0); // @[Top_AO.scala 407:50 Top_AO.scala 410:45 Top_AO.scala 415:47]
  assign Stack_manage_io_hitT_in = Arbitration_2_io_hit_out; // @[Top_AO.scala 764:44]
  assign Stack_manage_io_clear = Triangle_io_hitIndex_en & Triangle_io_RAY_AABB_1_out_IST3; // @[Top_AO.scala 89:54]
  assign Stack_manage_2_clock = clock;
  assign Stack_manage_2_reset = reset;
  assign Stack_manage_2_io_push = RAY_AABB_2_io_push & RAY_AABB_2_io_valid_out; // @[Top_AO.scala 419:28]
  assign Stack_manage_2_io_push_en = RAY_AABB_2_io_push & RAY_AABB_2_io_valid_out; // @[Top_AO.scala 419:28]
  assign Stack_manage_2_io_pop = Arbitration_2_2_io_valid_out; // @[Top_AO.scala 766:48]
  assign Stack_manage_2_io_pop_en = Arbitration_2_2_io_valid_out; // @[Top_AO.scala 767:44]
  assign Stack_manage_2_io_ray_id_push = RAY_AABB_2_io_push & RAY_AABB_2_io_valid_out ? RAY_AABB_2_io_rayid_out : 32'h0; // @[Top_AO.scala 419:54 Top_AO.scala 423:54 Top_AO.scala 428:55]
  assign Stack_manage_2_io_ray_id_pop = Arbitration_2_2_io_ray_id_out; // @[Top_AO.scala 768:40]
  assign Stack_manage_2_io_node_id_push_in = RAY_AABB_2_io_push & RAY_AABB_2_io_valid_out ? $signed(
    RAY_AABB_2_io_nodeIdx_0) : $signed(32'sh0); // @[Top_AO.scala 419:54 Top_AO.scala 422:47 Top_AO.scala 427:49]
  assign Stack_manage_2_io_hitT_in = Arbitration_2_2_io_hit_out; // @[Top_AO.scala 769:46]
  assign Stack_manage_2_io_clear = Triangle_io_hitIndex_en & Triangle_io_RAY_AABB_2_out_IST3; // @[Top_AO.scala 90:56]
  assign Triangle_clock = clock;
  assign Triangle_reset = reset;
  assign Triangle_io_To_IST0_enable = leaf_memory_valid; // @[Top_AO.scala 704:34 Top_AO.scala 705:42 Top_AO.scala 732:42]
  assign Triangle_io_nodeid_leaf = leaf_memory_valid ? $signed(leaf_node_id_temp) : $signed(32'sh0); // @[Top_AO.scala 704:34 Top_AO.scala 706:47 Top_AO.scala 733:47]
  assign Triangle_io_rayid_leaf = leaf_memory_valid ? ray_leaf_temp : 32'h0; // @[Top_AO.scala 704:34 Top_AO.scala 707:50 Top_AO.scala 734:50]
  assign Triangle_io_hiT_in = leaf_memory_valid ? hitT_temp : 32'h0; // @[Top_AO.scala 704:34 Top_AO.scala 708:54 Top_AO.scala 735:54]
  assign Triangle_io_v00_in_x = leaf_memory_valid ? TRI_RAM_x_io_v00_out : 32'h0; // @[Top_AO.scala 704:34 Top_AO.scala 709:52 Top_AO.scala 736:52]
  assign Triangle_io_v00_in_y = leaf_memory_valid ? TRI_RAM_y_io_v00_out : 32'h0; // @[Top_AO.scala 704:34 Top_AO.scala 711:52 Top_AO.scala 738:52]
  assign Triangle_io_v00_in_z = leaf_memory_valid ? TRI_RAM_z_io_v00_out : 32'h0; // @[Top_AO.scala 704:34 Top_AO.scala 712:52 Top_AO.scala 739:52]
  assign Triangle_io_v00_in_w = leaf_memory_valid ? TRI_RAM_w_io_v00_out : 32'h0; // @[Top_AO.scala 704:34 Top_AO.scala 713:51 Top_AO.scala 740:51]
  assign Triangle_io_v11_in_x = leaf_memory_valid ? TRI_RAM_x_io_v11_out : 32'h0; // @[Top_AO.scala 704:34 Top_AO.scala 714:52 Top_AO.scala 741:52]
  assign Triangle_io_v11_in_y = leaf_memory_valid ? TRI_RAM_y_io_v11_out : 32'h0; // @[Top_AO.scala 704:34 Top_AO.scala 715:52 Top_AO.scala 742:52]
  assign Triangle_io_v11_in_z = leaf_memory_valid ? TRI_RAM_z_io_v11_out : 32'h0; // @[Top_AO.scala 704:34 Top_AO.scala 716:52 Top_AO.scala 743:52]
  assign Triangle_io_v11_in_w = leaf_memory_valid ? TRI_RAM_w_io_v11_out : 32'h0; // @[Top_AO.scala 704:34 Top_AO.scala 717:51 Top_AO.scala 744:51]
  assign Triangle_io_v22_in_x = leaf_memory_valid ? TRI_RAM_x_io_v22_out : 32'h0; // @[Top_AO.scala 704:34 Top_AO.scala 718:52 Top_AO.scala 745:52]
  assign Triangle_io_v22_in_y = leaf_memory_valid ? TRI_RAM_y_io_v22_out : 32'h0; // @[Top_AO.scala 704:34 Top_AO.scala 719:52 Top_AO.scala 746:52]
  assign Triangle_io_v22_in_z = leaf_memory_valid ? TRI_RAM_z_io_v22_out : 32'h0; // @[Top_AO.scala 704:34 Top_AO.scala 720:52 Top_AO.scala 747:52]
  assign Triangle_io_v22_in_w = leaf_memory_valid ? TRI_RAM_w_io_v22_out : 32'h0; // @[Top_AO.scala 704:34 Top_AO.scala 721:51 Top_AO.scala 748:51]
  assign Triangle_io_ray_o_in_x = leaf_memory_valid ? Ray_origx_io_Ray_out : 32'h0; // @[Top_AO.scala 704:34 Top_AO.scala 722:50 Top_AO.scala 749:50]
  assign Triangle_io_ray_o_in_y = leaf_memory_valid ? Ray_origy_io_Ray_out : 32'h0; // @[Top_AO.scala 704:34 Top_AO.scala 723:50 Top_AO.scala 750:50]
  assign Triangle_io_ray_o_in_z = leaf_memory_valid ? Ray_origz_io_Ray_out : 32'h0; // @[Top_AO.scala 704:34 Top_AO.scala 724:50 Top_AO.scala 751:50]
  assign Triangle_io_ray_d_in_x = leaf_memory_valid ? Ray_dirx_io_Ray_out : 32'h0; // @[Top_AO.scala 704:34 Top_AO.scala 725:50 Top_AO.scala 752:50]
  assign Triangle_io_ray_d_in_y = leaf_memory_valid ? Ray_diry_io_Ray_out : 32'h0; // @[Top_AO.scala 704:34 Top_AO.scala 726:50 Top_AO.scala 753:50]
  assign Triangle_io_ray_d_in_z = leaf_memory_valid ? Ray_dirz_io_Ray_out : 32'h0; // @[Top_AO.scala 704:34 Top_AO.scala 727:50 Top_AO.scala 754:50]
  assign Triangle_io_break_in = leaf_memory_valid & TRI_RAM_x_io_valid == 32'h80000000; // @[Top_AO.scala 704:34 Top_AO.scala 710:51 Top_AO.scala 737:51]
  assign Triangle_io_RAY_AABB_1 = leaf_memory_valid & ray_aabb; // @[Top_AO.scala 704:34 Top_AO.scala 728:45 Top_AO.scala 755:45]
  assign Triangle_io_RAY_AABB_2 = leaf_memory_valid & ray_aabb_2; // @[Top_AO.scala 704:34 Top_AO.scala 729:45 Top_AO.scala 756:45]
  always @(posedge clock) begin
    if (reset) begin // @[Top_AO.scala 80:42]
      clock_counter <= 64'h0; // @[Top_AO.scala 80:42]
    end else begin
      clock_counter <= _T_1; // @[Top_AO.scala 81:36]
    end
    if (reset) begin // @[Top_AO.scala 135:54]
      memory_valid <= 1'h0; // @[Top_AO.scala 135:54]
    end else begin
      memory_valid <= _GEN_31;
    end
    if (reset) begin // @[Top_AO.scala 136:61]
      hit_temp <= 32'h0; // @[Top_AO.scala 136:61]
    end else if (Arbitration_1_io_valid_out & Arbitration_1_io_hit_out != 32'h0) begin // @[Top_AO.scala 140:70]
      hit_temp <= Arbitration_1_io_hit_out; // @[Top_AO.scala 148:51]
    end else begin
      hit_temp <= 32'h0;
    end
    if (reset) begin // @[Top_AO.scala 137:57]
      ray_id_temp <= 32'h0; // @[Top_AO.scala 137:57]
    end else if (Arbitration_1_io_valid_out & Arbitration_1_io_hit_out != 32'h0) begin // @[Top_AO.scala 140:70]
      ray_id_temp <= Arbitration_1_io_ray_id_out; // @[Top_AO.scala 163:59]
    end else if (Arbitration_1_io_valid_out & Arbitration_1_io_hit_out == 32'h0) begin // @[Top_AO.scala 165:76]
      ray_id_temp <= Arbitration_1_io_ray_id_out; // @[Top_AO.scala 189:59]
    end
    if (reset) begin // @[Top_AO.scala 138:57]
      hit_from_arb <= 1'h0; // @[Top_AO.scala 138:57]
    end else begin
      hit_from_arb <= _T_14;
    end
    if (reset) begin // @[Top_AO.scala 139:64]
      TRV_1 <= 64'h0; // @[Top_AO.scala 139:64]
    end else if (memory_valid) begin // @[Top_AO.scala 196:29]
      TRV_1 <= _T_48; // @[Top_AO.scala 228:70]
    end
    if (reset) begin // @[Top_AO.scala 270:56]
      memory_valid_2 <= 1'h0; // @[Top_AO.scala 270:56]
    end else begin
      memory_valid_2 <= _GEN_98;
    end
    if (reset) begin // @[Top_AO.scala 271:63]
      hit_temp_2 <= 32'h0; // @[Top_AO.scala 271:63]
    end else if (Arbitration_1_2_io_valid_out & Arbitration_1_2_io_hit_out != 32'h0) begin // @[Top_AO.scala 275:74]
      hit_temp_2 <= Arbitration_1_2_io_hit_out; // @[Top_AO.scala 285:65]
    end else begin
      hit_temp_2 <= 32'h0;
    end
    if (reset) begin // @[Top_AO.scala 272:59]
      ray_id_temp_2 <= 32'h0; // @[Top_AO.scala 272:59]
    end else if (Arbitration_1_2_io_valid_out & Arbitration_1_2_io_hit_out != 32'h0) begin // @[Top_AO.scala 275:74]
      ray_id_temp_2 <= Arbitration_1_2_io_ray_id_out; // @[Top_AO.scala 300:61]
    end else if (Arbitration_1_2_io_valid_out & Arbitration_1_2_io_hit_out == 32'h0) begin // @[Top_AO.scala 302:80]
      ray_id_temp_2 <= Arbitration_1_2_io_ray_id_out; // @[Top_AO.scala 328:61]
    end
    if (reset) begin // @[Top_AO.scala 273:59]
      hit_from_arb_2 <= 1'h0; // @[Top_AO.scala 273:59]
    end else begin
      hit_from_arb_2 <= _T_51;
    end
    if (reset) begin // @[Top_AO.scala 274:70]
      TRV_2 <= 64'h0; // @[Top_AO.scala 274:70]
    end else if (memory_valid_2) begin // @[Top_AO.scala 335:31]
      TRV_2 <= _T_85; // @[Top_AO.scala 364:76]
    end
    if (reset) begin // @[Top_AO.scala 672:58]
      leaf_memory_valid <= 1'h0; // @[Top_AO.scala 672:58]
    end else begin
      leaf_memory_valid <= _GEN_239;
    end
    if (reset) begin // @[Top_AO.scala 673:68]
      hitT_temp <= 32'h0; // @[Top_AO.scala 673:68]
    end else if (Arbitration_4_io_valid_out) begin // @[Top_AO.scala 679:37]
      hitT_temp <= Arbitration_4_io_hit_out; // @[Top_AO.scala 691:55]
    end else begin
      hitT_temp <= 32'h0; // @[Top_AO.scala 698:61]
    end
    if (reset) begin // @[Top_AO.scala 674:64]
      ray_leaf_temp <= 32'h0; // @[Top_AO.scala 674:64]
    end else if (Arbitration_4_io_valid_out) begin // @[Top_AO.scala 679:37]
      ray_leaf_temp <= Arbitration_4_io_ray_id_out; // @[Top_AO.scala 692:55]
    end else begin
      ray_leaf_temp <= 32'h0; // @[Top_AO.scala 699:57]
    end
    if (reset) begin // @[Top_AO.scala 675:57]
      leaf_node_id_temp <= 32'sh0; // @[Top_AO.scala 675:57]
    end else if (Arbitration_4_io_valid_out) begin // @[Top_AO.scala 679:37]
      leaf_node_id_temp <= Arbitration_4_io_node_id_out; // @[Top_AO.scala 693:55]
    end else begin
      leaf_node_id_temp <= 32'sh0; // @[Top_AO.scala 700:50]
    end
    if (reset) begin // @[Top_AO.scala 676:69]
      ray_aabb <= 1'h0; // @[Top_AO.scala 676:69]
    end else begin
      ray_aabb <= _GEN_245;
    end
    if (reset) begin // @[Top_AO.scala 677:71]
      ray_aabb_2 <= 1'h0; // @[Top_AO.scala 677:71]
    end else begin
      ray_aabb_2 <= _GEN_246;
    end
    if (reset) begin // @[Top_AO.scala 678:75]
      IST_1 <= 64'h0; // @[Top_AO.scala 678:75]
    end else if (leaf_memory_valid) begin // @[Top_AO.scala 704:34]
      IST_1 <= _T_165; // @[Top_AO.scala 730:67]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  clock_counter = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  memory_valid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  hit_temp = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  ray_id_temp = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  hit_from_arb = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  TRV_1 = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  memory_valid_2 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  hit_temp_2 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  ray_id_temp_2 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  hit_from_arb_2 = _RAND_9[0:0];
  _RAND_10 = {2{`RANDOM}};
  TRV_2 = _RAND_10[63:0];
  _RAND_11 = {1{`RANDOM}};
  leaf_memory_valid = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  hitT_temp = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  ray_leaf_temp = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  leaf_node_id_temp = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  ray_aabb = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  ray_aabb_2 = _RAND_16[0:0];
  _RAND_17 = {2{`RANDOM}};
  IST_1 = _RAND_17[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
