module ray_dispatch(
  input         clock,
  input         reset,
  input         io_dispatch,
  input         io_dispatch_2,
  output [31:0] io_rayid_id,
  output [31:0] io_rayid_id_2,
  output        io_ray_out,
  output        io_ray_out_2,
  output        io_ray_finish
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] count; // @[ray_dispatch.scala 21:37]
  reg [31:0] ray_id; // @[ray_dispatch.scala 22:37]
  reg [31:0] ray_id_2; // @[ray_dispatch.scala 23:33]
  reg  ray_out; // @[ray_dispatch.scala 25:35]
  reg  ray_out_2; // @[ray_dispatch.scala 26:32]
  reg [31:0] base; // @[ray_dispatch.scala 28:38]
  wire [31:0] _T_2 = count - 32'h2; // @[ray_dispatch.scala 33:39]
  wire [31:0] _T_5 = base + 32'h1; // @[ray_dispatch.scala 39:38]
  wire [31:0] _T_7 = base + 32'h2; // @[ray_dispatch.scala 40:35]
  wire  _GEN_5 = count >= 32'h1 | ray_out; // @[ray_dispatch.scala 38:27 ray_dispatch.scala 44:29 ray_dispatch.scala 25:35]
  wire  _GEN_6 = count >= 32'h1 | ray_out_2; // @[ray_dispatch.scala 38:27 ray_dispatch.scala 45:26 ray_dispatch.scala 26:32]
  wire  _GEN_11 = count == 32'h46 | _GEN_5; // @[ray_dispatch.scala 30:23 ray_dispatch.scala 35:29]
  wire  _GEN_12 = count == 32'h46 | _GEN_6; // @[ray_dispatch.scala 30:23 ray_dispatch.scala 36:26]
  wire [20:0] _T_17 = 21'h1e8480 - 21'h1; // @[ray_dispatch.scala 49:80]
  wire [31:0] _GEN_47 = {{11'd0}, _T_17}; // @[ray_dispatch.scala 49:67]
  wire  _T_18 = ray_id < _GEN_47; // @[ray_dispatch.scala 49:67]
  wire  _T_41 = io_dispatch & io_dispatch_2 & _T_18; // @[ray_dispatch.scala 65:63]
  wire [31:0] _GEN_19 = io_dispatch & io_dispatch_2 & _T_18 ? _T_5 : ray_id; // @[ray_dispatch.scala 65:91 ray_dispatch.scala 66:30]
  wire [31:0] _GEN_20 = io_dispatch & io_dispatch_2 & _T_18 ? _T_7 : ray_id_2; // @[ray_dispatch.scala 65:91 ray_dispatch.scala 67:27]
  wire [31:0] _GEN_21 = io_dispatch & io_dispatch_2 & _T_18 ? _T_7 : base; // @[ray_dispatch.scala 65:91 ray_dispatch.scala 68:31]
  wire  _GEN_29 = ~io_dispatch & io_dispatch_2 & _T_18 ? 1'h0 : _T_41; // @[ray_dispatch.scala 57:91 ray_dispatch.scala 62:28]
  wire  _GEN_30 = ~io_dispatch & io_dispatch_2 & _T_18 | _T_41; // @[ray_dispatch.scala 57:91 ray_dispatch.scala 63:26]
  wire  _GEN_36 = io_dispatch & ~io_dispatch_2 & ray_id < _GEN_47 | _GEN_29; // @[ray_dispatch.scala 49:85 ray_dispatch.scala 54:28]
  assign io_rayid_id = ray_id; // @[ray_dispatch.scala 104:25]
  assign io_rayid_id_2 = ray_id_2; // @[ray_dispatch.scala 105:22]
  assign io_ray_out = ray_out; // @[ray_dispatch.scala 107:25]
  assign io_ray_out_2 = ray_out_2; // @[ray_dispatch.scala 108:22]
  assign io_ray_finish = ray_id == 32'h1e8480; // @[ray_dispatch.scala 98:17]
  always @(posedge clock) begin
    if (reset) begin // @[ray_dispatch.scala 21:37]
      count <= 32'h46; // @[ray_dispatch.scala 21:37]
    end else if (count == 32'h46) begin // @[ray_dispatch.scala 30:23]
      count <= _T_2; // @[ray_dispatch.scala 33:30]
    end else if (count >= 32'h1) begin // @[ray_dispatch.scala 38:27]
      count <= _T_2; // @[ray_dispatch.scala 42:30]
    end
    if (reset) begin // @[ray_dispatch.scala 22:37]
      ray_id <= 32'h0; // @[ray_dispatch.scala 22:37]
    end else if (count == 32'h0) begin // @[ray_dispatch.scala 48:23]
      if (io_dispatch & ~io_dispatch_2 & ray_id < _GEN_47) begin // @[ray_dispatch.scala 49:85]
        ray_id <= _T_5; // @[ray_dispatch.scala 50:30]
      end else if (!(~io_dispatch & io_dispatch_2 & _T_18)) begin // @[ray_dispatch.scala 57:91]
        ray_id <= _GEN_19;
      end
    end else if (count == 32'h46) begin // @[ray_dispatch.scala 30:23]
      ray_id <= 32'h0; // @[ray_dispatch.scala 31:30]
    end else if (count >= 32'h1) begin // @[ray_dispatch.scala 38:27]
      ray_id <= _T_5; // @[ray_dispatch.scala 39:30]
    end
    if (reset) begin // @[ray_dispatch.scala 23:33]
      ray_id_2 <= 32'h0; // @[ray_dispatch.scala 23:33]
    end else if (count == 32'h0) begin // @[ray_dispatch.scala 48:23]
      if (!(io_dispatch & ~io_dispatch_2 & ray_id < _GEN_47)) begin // @[ray_dispatch.scala 49:85]
        if (~io_dispatch & io_dispatch_2 & _T_18) begin // @[ray_dispatch.scala 57:91]
          ray_id_2 <= _T_5; // @[ray_dispatch.scala 59:27]
        end else begin
          ray_id_2 <= _GEN_20;
        end
      end
    end else if (count == 32'h46) begin // @[ray_dispatch.scala 30:23]
      ray_id_2 <= 32'h1; // @[ray_dispatch.scala 32:27]
    end else if (count >= 32'h1) begin // @[ray_dispatch.scala 38:27]
      ray_id_2 <= _T_7; // @[ray_dispatch.scala 40:27]
    end
    if (reset) begin // @[ray_dispatch.scala 25:35]
      ray_out <= 1'h0; // @[ray_dispatch.scala 25:35]
    end else if (count == 32'h0) begin // @[ray_dispatch.scala 48:23]
      ray_out <= _GEN_36;
    end else begin
      ray_out <= _GEN_11;
    end
    if (reset) begin // @[ray_dispatch.scala 26:32]
      ray_out_2 <= 1'h0; // @[ray_dispatch.scala 26:32]
    end else if (count == 32'h0) begin // @[ray_dispatch.scala 48:23]
      if (io_dispatch & ~io_dispatch_2 & ray_id < _GEN_47) begin // @[ray_dispatch.scala 49:85]
        ray_out_2 <= 1'h0; // @[ray_dispatch.scala 55:25]
      end else begin
        ray_out_2 <= _GEN_30;
      end
    end else begin
      ray_out_2 <= _GEN_12;
    end
    if (reset) begin // @[ray_dispatch.scala 28:38]
      base <= 32'h0; // @[ray_dispatch.scala 28:38]
    end else if (count == 32'h0) begin // @[ray_dispatch.scala 48:23]
      if (io_dispatch & ~io_dispatch_2 & ray_id < _GEN_47) begin // @[ray_dispatch.scala 49:85]
        base <= _T_5; // @[ray_dispatch.scala 52:31]
      end else if (~io_dispatch & io_dispatch_2 & _T_18) begin // @[ray_dispatch.scala 57:91]
        base <= _T_5; // @[ray_dispatch.scala 60:31]
      end else begin
        base <= _GEN_21;
      end
    end else if (count == 32'h46) begin // @[ray_dispatch.scala 30:23]
      base <= 32'h1; // @[ray_dispatch.scala 37:33]
    end else if (count >= 32'h1) begin // @[ray_dispatch.scala 38:27]
      base <= _T_7; // @[ray_dispatch.scala 41:31]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  ray_id = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  ray_id_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  ray_out = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  ray_out_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  base = _RAND_5[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ray_memory(
  input         clock,
  input  [31:0] io_Ray_id,
  input  [31:0] io_Ray_id_2,
  output [31:0] io_Ray_out,
  output [31:0] io_Ray_out_2
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] mem [0:2073599]; // @[ray_memory.scala 16:26]
  wire [31:0] mem_MPORT_data; // @[ray_memory.scala 16:26]
  wire [20:0] mem_MPORT_addr; // @[ray_memory.scala 16:26]
  wire [31:0] mem_MPORT_1_data; // @[ray_memory.scala 16:26]
  wire [20:0] mem_MPORT_1_addr; // @[ray_memory.scala 16:26]
  wire [31:0] mem_MPORT_2_data; // @[ray_memory.scala 16:26]
  wire [20:0] mem_MPORT_2_addr; // @[ray_memory.scala 16:26]
  wire  mem_MPORT_2_mask; // @[ray_memory.scala 16:26]
  wire  mem_MPORT_2_en; // @[ray_memory.scala 16:26]
  reg [20:0] mem_MPORT_addr_pipe_0;
  reg [20:0] mem_MPORT_1_addr_pipe_0;
  assign mem_MPORT_addr = mem_MPORT_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_data = mem[mem_MPORT_addr]; // @[ray_memory.scala 16:26]
  `else
  assign mem_MPORT_data = mem_MPORT_addr >= 21'h1fa400 ? _RAND_1[31:0] : mem[mem_MPORT_addr]; // @[ray_memory.scala 16:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_1_addr = mem_MPORT_1_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_1_data = mem[mem_MPORT_1_addr]; // @[ray_memory.scala 16:26]
  `else
  assign mem_MPORT_1_data = mem_MPORT_1_addr >= 21'h1fa400 ? _RAND_2[31:0] : mem[mem_MPORT_1_addr]; // @[ray_memory.scala 16:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_2_data = 32'h0;
  assign mem_MPORT_2_addr = 21'h0;
  assign mem_MPORT_2_mask = 1'h1;
  assign mem_MPORT_2_en = 1'h0;
  assign io_Ray_out = mem_MPORT_data; // @[ray_memory.scala 18:16]
  assign io_Ray_out_2 = mem_MPORT_1_data; // @[ray_memory.scala 19:18]
  always @(posedge clock) begin
    if(mem_MPORT_2_en & mem_MPORT_2_mask) begin
      mem[mem_MPORT_2_addr] <= mem_MPORT_2_data; // @[ray_memory.scala 16:26]
    end
    mem_MPORT_addr_pipe_0 <= io_Ray_id[20:0];
    mem_MPORT_1_addr_pipe_0 <= io_Ray_id_2[20:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {1{`RANDOM}};
  _RAND_2 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2073600; initvar = initvar+1)
    mem[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  mem_MPORT_addr_pipe_0 = _RAND_3[20:0];
  _RAND_4 = {1{`RANDOM}};
  mem_MPORT_1_addr_pipe_0 = _RAND_4[20:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BVH_memory(
  input         clock,
  input  [31:0] io_BVH_id,
  input  [31:0] io_BVH_id_2,
  output [31:0] io_BVH_out,
  output [31:0] io_BVH_out_2
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg /* sparse */ [31:0] mem [0:21005099]; // @[BVH_memory.scala 16:26]
  wire [31:0] mem_MPORT_data; // @[BVH_memory.scala 16:26]
  wire [24:0] mem_MPORT_addr; // @[BVH_memory.scala 16:26]
  wire [31:0] mem_MPORT_1_data; // @[BVH_memory.scala 16:26]
  wire [24:0] mem_MPORT_1_addr; // @[BVH_memory.scala 16:26]
  wire [31:0] mem_MPORT_2_data; // @[BVH_memory.scala 16:26]
  wire [24:0] mem_MPORT_2_addr; // @[BVH_memory.scala 16:26]
  wire  mem_MPORT_2_mask; // @[BVH_memory.scala 16:26]
  wire  mem_MPORT_2_en; // @[BVH_memory.scala 16:26]
  reg [24:0] mem_MPORT_addr_pipe_0;
  reg [24:0] mem_MPORT_1_addr_pipe_0;
  wire [31:0] _T = io_BVH_id; // @[BVH_memory.scala 18:38]
  wire [31:0] _T_2 = io_BVH_id_2; // @[BVH_memory.scala 19:42]
  assign mem_MPORT_addr = mem_MPORT_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_data = mem[mem_MPORT_addr]; // @[BVH_memory.scala 16:26]
  `else
  assign mem_MPORT_data = mem_MPORT_addr >= 25'h140832c ? _RAND_1[31:0] : mem[mem_MPORT_addr]; // @[BVH_memory.scala 16:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_1_addr = mem_MPORT_1_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_1_data = mem[mem_MPORT_1_addr]; // @[BVH_memory.scala 16:26]
  `else
  assign mem_MPORT_1_data = mem_MPORT_1_addr >= 25'h140832c ? _RAND_2[31:0] : mem[mem_MPORT_1_addr]; // @[BVH_memory.scala 16:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_2_data = 32'h0;
  assign mem_MPORT_2_addr = 25'h0;
  assign mem_MPORT_2_mask = 1'h1;
  assign mem_MPORT_2_en = 1'h0;
  assign io_BVH_out = mem_MPORT_data; // @[BVH_memory.scala 18:16]
  assign io_BVH_out_2 = mem_MPORT_1_data; // @[BVH_memory.scala 19:18]
  always @(posedge clock) begin
    if(mem_MPORT_2_en & mem_MPORT_2_mask) begin
      mem[mem_MPORT_2_addr] <= mem_MPORT_2_data; // @[BVH_memory.scala 16:26]
    end
    mem_MPORT_addr_pipe_0 <= _T[24:0];
    mem_MPORT_1_addr_pipe_0 <= _T_2[24:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {1{`RANDOM}};
  _RAND_2 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 21005100; initvar = initvar+1)
    mem[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  mem_MPORT_addr_pipe_0 = _RAND_3[24:0];
  _RAND_4 = {1{`RANDOM}};
  mem_MPORT_1_addr_pipe_0 = _RAND_4[24:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BVH_memory_0(
  input         clock,
  input  [31:0] io_BVH_id,
  input  [31:0] io_BVH_id_2,
  output [31:0] io_BVH_out,
  output [31:0] io_BVH_out_2
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg /* sparse */ [31:0] mem [0:21005099]; // @[BVH_memory_0.scala 16:26]
  wire [31:0] mem_MPORT_data; // @[BVH_memory_0.scala 16:26]
  wire [24:0] mem_MPORT_addr; // @[BVH_memory_0.scala 16:26]
  wire [31:0] mem_MPORT_1_data; // @[BVH_memory_0.scala 16:26]
  wire [24:0] mem_MPORT_1_addr; // @[BVH_memory_0.scala 16:26]
  wire [31:0] mem_MPORT_2_data; // @[BVH_memory_0.scala 16:26]
  wire [24:0] mem_MPORT_2_addr; // @[BVH_memory_0.scala 16:26]
  wire  mem_MPORT_2_mask; // @[BVH_memory_0.scala 16:26]
  wire  mem_MPORT_2_en; // @[BVH_memory_0.scala 16:26]
  reg [24:0] mem_MPORT_addr_pipe_0;
  reg [24:0] mem_MPORT_1_addr_pipe_0;
  wire [31:0] _T = io_BVH_id; // @[BVH_memory_0.scala 18:38]
  wire [31:0] _T_2 = io_BVH_id_2; // @[BVH_memory_0.scala 19:42]
  assign mem_MPORT_addr = mem_MPORT_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_data = mem[mem_MPORT_addr]; // @[BVH_memory_0.scala 16:26]
  `else
  assign mem_MPORT_data = mem_MPORT_addr >= 25'h140832c ? _RAND_1[31:0] : mem[mem_MPORT_addr]; // @[BVH_memory_0.scala 16:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_1_addr = mem_MPORT_1_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_1_data = mem[mem_MPORT_1_addr]; // @[BVH_memory_0.scala 16:26]
  `else
  assign mem_MPORT_1_data = mem_MPORT_1_addr >= 25'h140832c ? _RAND_2[31:0] : mem[mem_MPORT_1_addr]; // @[BVH_memory_0.scala 16:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_2_data = 32'sh0;
  assign mem_MPORT_2_addr = 25'h0;
  assign mem_MPORT_2_mask = 1'h1;
  assign mem_MPORT_2_en = 1'h0;
  assign io_BVH_out = mem_MPORT_data; // @[BVH_memory_0.scala 18:16]
  assign io_BVH_out_2 = mem_MPORT_1_data; // @[BVH_memory_0.scala 19:18]
  always @(posedge clock) begin
    if(mem_MPORT_2_en & mem_MPORT_2_mask) begin
      mem[mem_MPORT_2_addr] <= mem_MPORT_2_data; // @[BVH_memory_0.scala 16:26]
    end
    mem_MPORT_addr_pipe_0 <= _T[24:0];
    mem_MPORT_1_addr_pipe_0 <= _T_2[24:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {1{`RANDOM}};
  _RAND_2 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 21005100; initvar = initvar+1)
    mem[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  mem_MPORT_addr_pipe_0 = _RAND_3[24:0];
  _RAND_4 = {1{`RANDOM}};
  mem_MPORT_1_addr_pipe_0 = _RAND_4[24:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Triangle_memory_valid(
  input         clock,
  input  [31:0] io_Triangle_id,
  output [31:0] io_v00_out,
  output [31:0] io_v11_out,
  output [31:0] io_v22_out,
  output [31:0] io_valid
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg /* sparse */ [31:0] mem [0:21005099]; // @[Triangle_memory_valid.scala 18:26]
  wire [31:0] mem_MPORT_data; // @[Triangle_memory_valid.scala 18:26]
  wire [24:0] mem_MPORT_addr; // @[Triangle_memory_valid.scala 18:26]
  wire [31:0] mem_MPORT_1_data; // @[Triangle_memory_valid.scala 18:26]
  wire [24:0] mem_MPORT_1_addr; // @[Triangle_memory_valid.scala 18:26]
  wire [31:0] mem_MPORT_2_data; // @[Triangle_memory_valid.scala 18:26]
  wire [24:0] mem_MPORT_2_addr; // @[Triangle_memory_valid.scala 18:26]
  wire [31:0] mem_MPORT_3_data; // @[Triangle_memory_valid.scala 18:26]
  wire [24:0] mem_MPORT_3_addr; // @[Triangle_memory_valid.scala 18:26]
  wire [31:0] mem_MPORT_4_data; // @[Triangle_memory_valid.scala 18:26]
  wire [24:0] mem_MPORT_4_addr; // @[Triangle_memory_valid.scala 18:26]
  wire  mem_MPORT_4_mask; // @[Triangle_memory_valid.scala 18:26]
  wire  mem_MPORT_4_en; // @[Triangle_memory_valid.scala 18:26]
  reg [24:0] mem_MPORT_addr_pipe_0;
  reg [24:0] mem_MPORT_1_addr_pipe_0;
  reg [24:0] mem_MPORT_2_addr_pipe_0;
  reg [24:0] mem_MPORT_3_addr_pipe_0;
  wire [31:0] _T = io_Triangle_id; // @[Triangle_memory_valid.scala 20:43]
  wire [31:0] _T_4 = io_Triangle_id + 32'h1; // @[Triangle_memory_valid.scala 21:49]
  wire [31:0] _T_8 = io_Triangle_id + 32'h2; // @[Triangle_memory_valid.scala 22:49]
  wire [31:0] _T_12 = io_Triangle_id + 32'h3; // @[Triangle_memory_valid.scala 23:47]
  assign mem_MPORT_addr = mem_MPORT_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_data = mem[mem_MPORT_addr]; // @[Triangle_memory_valid.scala 18:26]
  `else
  assign mem_MPORT_data = mem_MPORT_addr >= 25'h140832c ? _RAND_1[31:0] : mem[mem_MPORT_addr]; // @[Triangle_memory_valid.scala 18:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_1_addr = mem_MPORT_1_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_1_data = mem[mem_MPORT_1_addr]; // @[Triangle_memory_valid.scala 18:26]
  `else
  assign mem_MPORT_1_data = mem_MPORT_1_addr >= 25'h140832c ? _RAND_2[31:0] : mem[mem_MPORT_1_addr]; // @[Triangle_memory_valid.scala 18:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_2_addr = mem_MPORT_2_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_2_data = mem[mem_MPORT_2_addr]; // @[Triangle_memory_valid.scala 18:26]
  `else
  assign mem_MPORT_2_data = mem_MPORT_2_addr >= 25'h140832c ? _RAND_3[31:0] : mem[mem_MPORT_2_addr]; // @[Triangle_memory_valid.scala 18:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_3_addr = mem_MPORT_3_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_3_data = mem[mem_MPORT_3_addr]; // @[Triangle_memory_valid.scala 18:26]
  `else
  assign mem_MPORT_3_data = mem_MPORT_3_addr >= 25'h140832c ? _RAND_4[31:0] : mem[mem_MPORT_3_addr]; // @[Triangle_memory_valid.scala 18:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_4_data = 32'h0;
  assign mem_MPORT_4_addr = 25'h0;
  assign mem_MPORT_4_mask = 1'h1;
  assign mem_MPORT_4_en = 1'h0;
  assign io_v00_out = mem_MPORT_data; // @[Triangle_memory_valid.scala 20:16]
  assign io_v11_out = mem_MPORT_1_data; // @[Triangle_memory_valid.scala 21:16]
  assign io_v22_out = mem_MPORT_2_data; // @[Triangle_memory_valid.scala 22:16]
  assign io_valid = mem_MPORT_3_data; // @[Triangle_memory_valid.scala 23:14]
  always @(posedge clock) begin
    if(mem_MPORT_4_en & mem_MPORT_4_mask) begin
      mem[mem_MPORT_4_addr] <= mem_MPORT_4_data; // @[Triangle_memory_valid.scala 18:26]
    end
    mem_MPORT_addr_pipe_0 <= _T[24:0];
    mem_MPORT_1_addr_pipe_0 <= _T_4[24:0];
    mem_MPORT_2_addr_pipe_0 <= _T_8[24:0];
    mem_MPORT_3_addr_pipe_0 <= _T_12[24:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {1{`RANDOM}};
  _RAND_2 = {1{`RANDOM}};
  _RAND_3 = {1{`RANDOM}};
  _RAND_4 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 21005100; initvar = initvar+1)
    mem[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  mem_MPORT_addr_pipe_0 = _RAND_5[24:0];
  _RAND_6 = {1{`RANDOM}};
  mem_MPORT_1_addr_pipe_0 = _RAND_6[24:0];
  _RAND_7 = {1{`RANDOM}};
  mem_MPORT_2_addr_pipe_0 = _RAND_7[24:0];
  _RAND_8 = {1{`RANDOM}};
  mem_MPORT_3_addr_pipe_0 = _RAND_8[24:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Triangle_memory(
  input         clock,
  input  [31:0] io_Triangle_id,
  output [31:0] io_v00_out,
  output [31:0] io_v11_out,
  output [31:0] io_v22_out
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg /* sparse */ [31:0] mem [0:21005099]; // @[Triangle_memory.scala 16:26]
  wire [31:0] mem_MPORT_data; // @[Triangle_memory.scala 16:26]
  wire [24:0] mem_MPORT_addr; // @[Triangle_memory.scala 16:26]
  wire [31:0] mem_MPORT_1_data; // @[Triangle_memory.scala 16:26]
  wire [24:0] mem_MPORT_1_addr; // @[Triangle_memory.scala 16:26]
  wire [31:0] mem_MPORT_2_data; // @[Triangle_memory.scala 16:26]
  wire [24:0] mem_MPORT_2_addr; // @[Triangle_memory.scala 16:26]
  wire [31:0] mem_MPORT_3_data; // @[Triangle_memory.scala 16:26]
  wire [24:0] mem_MPORT_3_addr; // @[Triangle_memory.scala 16:26]
  wire  mem_MPORT_3_mask; // @[Triangle_memory.scala 16:26]
  wire  mem_MPORT_3_en; // @[Triangle_memory.scala 16:26]
  reg [24:0] mem_MPORT_addr_pipe_0;
  reg [24:0] mem_MPORT_1_addr_pipe_0;
  reg [24:0] mem_MPORT_2_addr_pipe_0;
  wire [31:0] _T = io_Triangle_id; // @[Triangle_memory.scala 18:43]
  wire [31:0] _T_4 = io_Triangle_id + 32'h1; // @[Triangle_memory.scala 19:49]
  wire [31:0] _T_8 = io_Triangle_id + 32'h2; // @[Triangle_memory.scala 20:49]
  assign mem_MPORT_addr = mem_MPORT_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_data = mem[mem_MPORT_addr]; // @[Triangle_memory.scala 16:26]
  `else
  assign mem_MPORT_data = mem_MPORT_addr >= 25'h140832c ? _RAND_1[31:0] : mem[mem_MPORT_addr]; // @[Triangle_memory.scala 16:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_1_addr = mem_MPORT_1_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_1_data = mem[mem_MPORT_1_addr]; // @[Triangle_memory.scala 16:26]
  `else
  assign mem_MPORT_1_data = mem_MPORT_1_addr >= 25'h140832c ? _RAND_2[31:0] : mem[mem_MPORT_1_addr]; // @[Triangle_memory.scala 16:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_2_addr = mem_MPORT_2_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_2_data = mem[mem_MPORT_2_addr]; // @[Triangle_memory.scala 16:26]
  `else
  assign mem_MPORT_2_data = mem_MPORT_2_addr >= 25'h140832c ? _RAND_3[31:0] : mem[mem_MPORT_2_addr]; // @[Triangle_memory.scala 16:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_3_data = 32'h0;
  assign mem_MPORT_3_addr = 25'h0;
  assign mem_MPORT_3_mask = 1'h1;
  assign mem_MPORT_3_en = 1'h0;
  assign io_v00_out = mem_MPORT_data; // @[Triangle_memory.scala 18:16]
  assign io_v11_out = mem_MPORT_1_data; // @[Triangle_memory.scala 19:16]
  assign io_v22_out = mem_MPORT_2_data; // @[Triangle_memory.scala 20:16]
  always @(posedge clock) begin
    if(mem_MPORT_3_en & mem_MPORT_3_mask) begin
      mem[mem_MPORT_3_addr] <= mem_MPORT_3_data; // @[Triangle_memory.scala 16:26]
    end
    mem_MPORT_addr_pipe_0 <= _T[24:0];
    mem_MPORT_1_addr_pipe_0 <= _T_4[24:0];
    mem_MPORT_2_addr_pipe_0 <= _T_8[24:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {1{`RANDOM}};
  _RAND_2 = {1{`RANDOM}};
  _RAND_3 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 21005100; initvar = initvar+1)
    mem[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  mem_MPORT_addr_pipe_0 = _RAND_4[24:0];
  _RAND_5 = {1{`RANDOM}};
  mem_MPORT_1_addr_pipe_0 = _RAND_5[24:0];
  _RAND_6 = {1{`RANDOM}};
  mem_MPORT_2_addr_pipe_0 = _RAND_6[24:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MulAddRecFNToRaw_preMul(
  input  [32:0] io_a,
  input  [32:0] io_b,
  input  [32:0] io_c,
  output [23:0] io_mulAddA,
  output [23:0] io_mulAddB,
  output [47:0] io_mulAddC,
  output        io_toPostMul_isSigNaNAny,
  output        io_toPostMul_isNaNAOrB,
  output        io_toPostMul_isInfA,
  output        io_toPostMul_isZeroA,
  output        io_toPostMul_isInfB,
  output        io_toPostMul_isZeroB,
  output        io_toPostMul_signProd,
  output        io_toPostMul_isNaNC,
  output        io_toPostMul_isInfC,
  output        io_toPostMul_isZeroC,
  output [9:0]  io_toPostMul_sExpSum,
  output        io_toPostMul_doSubMags,
  output        io_toPostMul_CIsDominant,
  output [4:0]  io_toPostMul_CDom_CAlignDist,
  output [25:0] io_toPostMul_highAlignedSigC,
  output        io_toPostMul_bit0AlignedSigC
);
  wire  rawA_isZero = io_a[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_4 = io_a[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawA_isNaN = _T_4 & io_a[29]; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawA_sign = io_a[32]; // @[rawFloatFromRecFN.scala 58:25]
  wire [9:0] rawA_sExp = {1'b0,$signed(io_a[31:23])}; // @[rawFloatFromRecFN.scala 59:27]
  wire  hi_lo = ~rawA_isZero; // @[rawFloatFromRecFN.scala 60:39]
  wire [22:0] lo = io_a[22:0]; // @[rawFloatFromRecFN.scala 60:51]
  wire [24:0] rawA_sig = {1'h0,hi_lo,lo}; // @[Cat.scala 30:58]
  wire  rawB_isZero = io_b[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_17 = io_b[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawB_isNaN = _T_17 & io_b[29]; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawB_sign = io_b[32]; // @[rawFloatFromRecFN.scala 58:25]
  wire [9:0] rawB_sExp = {1'b0,$signed(io_b[31:23])}; // @[rawFloatFromRecFN.scala 59:27]
  wire  hi_lo_1 = ~rawB_isZero; // @[rawFloatFromRecFN.scala 60:39]
  wire [22:0] lo_1 = io_b[22:0]; // @[rawFloatFromRecFN.scala 60:51]
  wire [24:0] rawB_sig = {1'h0,hi_lo_1,lo_1}; // @[Cat.scala 30:58]
  wire  rawC_isZero = io_c[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_30 = io_c[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawC_isNaN = _T_30 & io_c[29]; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawC_sign = io_c[32]; // @[rawFloatFromRecFN.scala 58:25]
  wire [9:0] rawC_sExp = {1'b0,$signed(io_c[31:23])}; // @[rawFloatFromRecFN.scala 59:27]
  wire  hi_lo_2 = ~rawC_isZero; // @[rawFloatFromRecFN.scala 60:39]
  wire [22:0] lo_2 = io_c[22:0]; // @[rawFloatFromRecFN.scala 60:51]
  wire [24:0] rawC_sig = {1'h0,hi_lo_2,lo_2}; // @[Cat.scala 30:58]
  wire  signProd = rawA_sign ^ rawB_sign; // @[MulAddRecFN.scala 98:30]
  wire [10:0] _T_41 = $signed(rawA_sExp) + $signed(rawB_sExp); // @[MulAddRecFN.scala 101:19]
  wire [10:0] sExpAlignedProd = $signed(_T_41) - 11'she5; // @[MulAddRecFN.scala 101:32]
  wire  doSubMags = signProd ^ rawC_sign; // @[MulAddRecFN.scala 103:30]
  wire [10:0] _GEN_0 = {{1{rawC_sExp[9]}},rawC_sExp}; // @[MulAddRecFN.scala 107:42]
  wire [10:0] sNatCAlignDist = $signed(sExpAlignedProd) - $signed(_GEN_0); // @[MulAddRecFN.scala 107:42]
  wire [9:0] posNatCAlignDist = sNatCAlignDist[9:0]; // @[MulAddRecFN.scala 108:42]
  wire  isMinCAlign = rawA_isZero | rawB_isZero | $signed(sNatCAlignDist) < 11'sh0; // @[MulAddRecFN.scala 109:50]
  wire  CIsDominant = hi_lo_2 & (isMinCAlign | posNatCAlignDist <= 10'h18); // @[MulAddRecFN.scala 111:23]
  wire [6:0] _T_55 = posNatCAlignDist < 10'h4a ? posNatCAlignDist[6:0] : 7'h4a; // @[MulAddRecFN.scala 115:16]
  wire [6:0] CAlignDist = isMinCAlign ? 7'h0 : _T_55; // @[MulAddRecFN.scala 113:12]
  wire [24:0] _T_56 = ~rawC_sig; // @[MulAddRecFN.scala 121:28]
  wire [24:0] hi_3 = doSubMags ? _T_56 : rawC_sig; // @[MulAddRecFN.scala 121:16]
  wire [52:0] lo_3 = doSubMags ? 53'h1fffffffffffff : 53'h0; // @[Bitwise.scala 72:12]
  wire [77:0] _T_59 = {hi_3,lo_3}; // @[MulAddRecFN.scala 123:11]
  wire [77:0] mainAlignedSigC = $signed(_T_59) >>> CAlignDist; // @[MulAddRecFN.scala 123:17]
  wire [26:0] _T_60 = {rawC_sig, 2'h0}; // @[MulAddRecFN.scala 125:30]
  wire  _T_62 = |_T_60[3:0]; // @[primitives.scala 121:54]
  wire  _T_64 = |_T_60[7:4]; // @[primitives.scala 121:54]
  wire  _T_66 = |_T_60[11:8]; // @[primitives.scala 121:54]
  wire  _T_68 = |_T_60[15:12]; // @[primitives.scala 121:54]
  wire  _T_70 = |_T_60[19:16]; // @[primitives.scala 121:54]
  wire  _T_72 = |_T_60[23:20]; // @[primitives.scala 121:54]
  wire  _T_74 = |_T_60[26:24]; // @[primitives.scala 124:57]
  wire [6:0] _T_75 = {_T_74,_T_72,_T_70,_T_68,_T_66,_T_64,_T_62}; // @[primitives.scala 125:20]
  wire [32:0] _T_77 = 33'sh100000000 >>> CAlignDist[6:2]; // @[primitives.scala 77:58]
  wire  hi_5 = _T_77[14]; // @[Bitwise.scala 109:18]
  wire  lo_5 = _T_77[15]; // @[Bitwise.scala 109:44]
  wire  hi_7 = _T_77[16]; // @[Bitwise.scala 109:18]
  wire  lo_6 = _T_77[17]; // @[Bitwise.scala 109:44]
  wire  hi_9 = _T_77[18]; // @[Bitwise.scala 109:18]
  wire  lo_8 = _T_77[19]; // @[Bitwise.scala 109:44]
  wire [5:0] _T_83 = {hi_5,lo_5,hi_7,lo_6,hi_9,lo_8}; // @[Cat.scala 30:58]
  wire [6:0] _GEN_1 = {{1'd0}, _T_83}; // @[MulAddRecFN.scala 125:68]
  wire [6:0] _T_84 = _T_75 & _GEN_1; // @[MulAddRecFN.scala 125:68]
  wire  reduced4CExtra = |_T_84; // @[MulAddRecFN.scala 133:11]
  wire  _T_89 = &mainAlignedSigC[2:0] & ~reduced4CExtra; // @[MulAddRecFN.scala 137:44]
  wire  _T_92 = |mainAlignedSigC[2:0] | reduced4CExtra; // @[MulAddRecFN.scala 138:44]
  wire  lo_10 = doSubMags ? _T_89 : _T_92; // @[MulAddRecFN.scala 136:16]
  wire [74:0] hi_10 = mainAlignedSigC[77:3]; // @[Cat.scala 30:58]
  wire [75:0] alignedSigC = {hi_10,lo_10}; // @[Cat.scala 30:58]
  wire  _T_96 = rawA_isNaN & ~rawA_sig[22]; // @[common.scala 81:46]
  wire  _T_99 = rawB_isNaN & ~rawB_sig[22]; // @[common.scala 81:46]
  wire  _T_103 = rawC_isNaN & ~rawC_sig[22]; // @[common.scala 81:46]
  wire [10:0] _T_108 = $signed(sExpAlignedProd) - 11'sh18; // @[MulAddRecFN.scala 161:53]
  wire [10:0] _T_109 = CIsDominant ? $signed({{1{rawC_sExp[9]}},rawC_sExp}) : $signed(_T_108); // @[MulAddRecFN.scala 161:12]
  assign io_mulAddA = rawA_sig[23:0]; // @[MulAddRecFN.scala 144:16]
  assign io_mulAddB = rawB_sig[23:0]; // @[MulAddRecFN.scala 145:16]
  assign io_mulAddC = alignedSigC[48:1]; // @[MulAddRecFN.scala 146:30]
  assign io_toPostMul_isSigNaNAny = _T_96 | _T_99 | _T_103; // @[MulAddRecFN.scala 149:58]
  assign io_toPostMul_isNaNAOrB = rawA_isNaN | rawB_isNaN; // @[MulAddRecFN.scala 151:42]
  assign io_toPostMul_isInfA = _T_4 & ~io_a[29]; // @[rawFloatFromRecFN.scala 56:33]
  assign io_toPostMul_isZeroA = io_a[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign io_toPostMul_isInfB = _T_17 & ~io_b[29]; // @[rawFloatFromRecFN.scala 56:33]
  assign io_toPostMul_isZeroB = io_b[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign io_toPostMul_signProd = rawA_sign ^ rawB_sign; // @[MulAddRecFN.scala 98:30]
  assign io_toPostMul_isNaNC = _T_30 & io_c[29]; // @[rawFloatFromRecFN.scala 55:33]
  assign io_toPostMul_isInfC = _T_30 & ~io_c[29]; // @[rawFloatFromRecFN.scala 56:33]
  assign io_toPostMul_isZeroC = io_c[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign io_toPostMul_sExpSum = _T_109[9:0]; // @[MulAddRecFN.scala 160:28]
  assign io_toPostMul_doSubMags = signProd ^ rawC_sign; // @[MulAddRecFN.scala 103:30]
  assign io_toPostMul_CIsDominant = hi_lo_2 & (isMinCAlign | posNatCAlignDist <= 10'h18); // @[MulAddRecFN.scala 111:23]
  assign io_toPostMul_CDom_CAlignDist = CAlignDist[4:0]; // @[MulAddRecFN.scala 164:47]
  assign io_toPostMul_highAlignedSigC = alignedSigC[74:49]; // @[MulAddRecFN.scala 166:20]
  assign io_toPostMul_bit0AlignedSigC = alignedSigC[0]; // @[MulAddRecFN.scala 167:48]
endmodule
module MulAddRecFNToRaw_postMul(
  input         io_fromPreMul_isSigNaNAny,
  input         io_fromPreMul_isNaNAOrB,
  input         io_fromPreMul_isInfA,
  input         io_fromPreMul_isZeroA,
  input         io_fromPreMul_isInfB,
  input         io_fromPreMul_isZeroB,
  input         io_fromPreMul_signProd,
  input         io_fromPreMul_isNaNC,
  input         io_fromPreMul_isInfC,
  input         io_fromPreMul_isZeroC,
  input  [9:0]  io_fromPreMul_sExpSum,
  input         io_fromPreMul_doSubMags,
  input         io_fromPreMul_CIsDominant,
  input  [4:0]  io_fromPreMul_CDom_CAlignDist,
  input  [25:0] io_fromPreMul_highAlignedSigC,
  input         io_fromPreMul_bit0AlignedSigC,
  input  [48:0] io_mulAddResult,
  output        io_invalidExc,
  output        io_rawOut_isNaN,
  output        io_rawOut_isInf,
  output        io_rawOut_isZero,
  output        io_rawOut_sign,
  output [9:0]  io_rawOut_sExp,
  output [26:0] io_rawOut_sig
);
  wire  CDom_sign = io_fromPreMul_signProd ^ io_fromPreMul_doSubMags; // @[MulAddRecFN.scala 192:42]
  wire [25:0] _T_2 = io_fromPreMul_highAlignedSigC + 26'h1; // @[MulAddRecFN.scala 195:47]
  wire [25:0] hi_hi = io_mulAddResult[48] ? _T_2 : io_fromPreMul_highAlignedSigC; // @[MulAddRecFN.scala 194:16]
  wire [47:0] hi_lo = io_mulAddResult[47:0]; // @[MulAddRecFN.scala 198:28]
  wire [74:0] sigSum = {hi_hi,hi_lo,io_fromPreMul_bit0AlignedSigC}; // @[Cat.scala 30:58]
  wire [1:0] _T_3 = {1'b0,$signed(io_fromPreMul_doSubMags)}; // @[MulAddRecFN.scala 205:69]
  wire [9:0] _GEN_0 = {{8{_T_3[1]}},_T_3}; // @[MulAddRecFN.scala 205:43]
  wire [9:0] CDom_sExp = $signed(io_fromPreMul_sExpSum) - $signed(_GEN_0); // @[MulAddRecFN.scala 205:43]
  wire [49:0] _T_7 = ~sigSum[74:25]; // @[MulAddRecFN.scala 208:13]
  wire [1:0] hi_lo_1 = io_fromPreMul_highAlignedSigC[25:24]; // @[MulAddRecFN.scala 211:46]
  wire [46:0] lo = sigSum[72:26]; // @[MulAddRecFN.scala 212:23]
  wire [49:0] _T_8 = {1'h0,hi_lo_1,lo}; // @[Cat.scala 30:58]
  wire [49:0] CDom_absSigSum = io_fromPreMul_doSubMags ? _T_7 : _T_8; // @[MulAddRecFN.scala 207:12]
  wire [23:0] _T_10 = ~sigSum[24:1]; // @[MulAddRecFN.scala 217:14]
  wire  _T_11 = |_T_10; // @[MulAddRecFN.scala 217:36]
  wire  _T_13 = |sigSum[25:1]; // @[MulAddRecFN.scala 218:37]
  wire  CDom_absSigSumExtra = io_fromPreMul_doSubMags ? _T_11 : _T_13; // @[MulAddRecFN.scala 216:12]
  wire [80:0] _GEN_1 = {{31'd0}, CDom_absSigSum}; // @[MulAddRecFN.scala 221:24]
  wire [80:0] _T_14 = _GEN_1 << io_fromPreMul_CDom_CAlignDist; // @[MulAddRecFN.scala 221:24]
  wire [28:0] CDom_mainSig = _T_14[49:21]; // @[MulAddRecFN.scala 221:56]
  wire [26:0] _T_16 = {CDom_absSigSum[23:0], 3'h0}; // @[MulAddRecFN.scala 224:53]
  wire  _T_18 = |_T_16[3:0]; // @[primitives.scala 121:54]
  wire  _T_20 = |_T_16[7:4]; // @[primitives.scala 121:54]
  wire  _T_22 = |_T_16[11:8]; // @[primitives.scala 121:54]
  wire  _T_24 = |_T_16[15:12]; // @[primitives.scala 121:54]
  wire  _T_26 = |_T_16[19:16]; // @[primitives.scala 121:54]
  wire  _T_28 = |_T_16[23:20]; // @[primitives.scala 121:54]
  wire  _T_30 = |_T_16[26:24]; // @[primitives.scala 124:57]
  wire [6:0] _T_31 = {_T_30,_T_28,_T_26,_T_24,_T_22,_T_20,_T_18}; // @[primitives.scala 125:20]
  wire [2:0] _T_33 = ~io_fromPreMul_CDom_CAlignDist[4:2]; // @[primitives.scala 51:21]
  wire [8:0] _T_34 = 9'sh100 >>> _T_33; // @[primitives.scala 77:58]
  wire  hi_3 = _T_34[1]; // @[Bitwise.scala 109:18]
  wire  lo_2 = _T_34[2]; // @[Bitwise.scala 109:44]
  wire  hi_5 = _T_34[3]; // @[Bitwise.scala 109:18]
  wire  lo_3 = _T_34[4]; // @[Bitwise.scala 109:44]
  wire  hi_7 = _T_34[5]; // @[Bitwise.scala 109:18]
  wire  lo_5 = _T_34[6]; // @[Bitwise.scala 109:44]
  wire [5:0] _T_40 = {hi_3,lo_2,hi_5,lo_3,hi_7,lo_5}; // @[Cat.scala 30:58]
  wire [6:0] _GEN_2 = {{1'd0}, _T_40}; // @[MulAddRecFN.scala 224:72]
  wire [6:0] _T_41 = _T_31 & _GEN_2; // @[MulAddRecFN.scala 224:72]
  wire  CDom_reduced4SigExtra = |_T_41; // @[MulAddRecFN.scala 225:73]
  wire [25:0] hi_8 = CDom_mainSig[28:3]; // @[MulAddRecFN.scala 227:25]
  wire  lo_7 = |CDom_mainSig[2:0] | CDom_reduced4SigExtra | CDom_absSigSumExtra; // @[MulAddRecFN.scala 228:61]
  wire [26:0] CDom_sig = {hi_8,lo_7}; // @[Cat.scala 30:58]
  wire  notCDom_signSigSum = sigSum[51]; // @[MulAddRecFN.scala 234:36]
  wire [50:0] _T_46 = ~sigSum[50:0]; // @[MulAddRecFN.scala 237:13]
  wire [50:0] _GEN_3 = {{50'd0}, io_fromPreMul_doSubMags}; // @[MulAddRecFN.scala 238:41]
  wire [50:0] _T_49 = sigSum[50:0] + _GEN_3; // @[MulAddRecFN.scala 238:41]
  wire [50:0] notCDom_absSigSum = notCDom_signSigSum ? _T_46 : _T_49; // @[MulAddRecFN.scala 236:12]
  wire  _T_51 = |notCDom_absSigSum[1:0]; // @[primitives.scala 104:54]
  wire  _T_53 = |notCDom_absSigSum[3:2]; // @[primitives.scala 104:54]
  wire  _T_55 = |notCDom_absSigSum[5:4]; // @[primitives.scala 104:54]
  wire  _T_57 = |notCDom_absSigSum[7:6]; // @[primitives.scala 104:54]
  wire  _T_59 = |notCDom_absSigSum[9:8]; // @[primitives.scala 104:54]
  wire  _T_61 = |notCDom_absSigSum[11:10]; // @[primitives.scala 104:54]
  wire  _T_63 = |notCDom_absSigSum[13:12]; // @[primitives.scala 104:54]
  wire  _T_65 = |notCDom_absSigSum[15:14]; // @[primitives.scala 104:54]
  wire  _T_67 = |notCDom_absSigSum[17:16]; // @[primitives.scala 104:54]
  wire  _T_69 = |notCDom_absSigSum[19:18]; // @[primitives.scala 104:54]
  wire  _T_71 = |notCDom_absSigSum[21:20]; // @[primitives.scala 104:54]
  wire  _T_73 = |notCDom_absSigSum[23:22]; // @[primitives.scala 104:54]
  wire  _T_75 = |notCDom_absSigSum[25:24]; // @[primitives.scala 104:54]
  wire  _T_77 = |notCDom_absSigSum[27:26]; // @[primitives.scala 104:54]
  wire  _T_79 = |notCDom_absSigSum[29:28]; // @[primitives.scala 104:54]
  wire  _T_81 = |notCDom_absSigSum[31:30]; // @[primitives.scala 104:54]
  wire  _T_83 = |notCDom_absSigSum[33:32]; // @[primitives.scala 104:54]
  wire  _T_85 = |notCDom_absSigSum[35:34]; // @[primitives.scala 104:54]
  wire  _T_87 = |notCDom_absSigSum[37:36]; // @[primitives.scala 104:54]
  wire  _T_89 = |notCDom_absSigSum[39:38]; // @[primitives.scala 104:54]
  wire  _T_91 = |notCDom_absSigSum[41:40]; // @[primitives.scala 104:54]
  wire  _T_93 = |notCDom_absSigSum[43:42]; // @[primitives.scala 104:54]
  wire  _T_95 = |notCDom_absSigSum[45:44]; // @[primitives.scala 104:54]
  wire  _T_97 = |notCDom_absSigSum[47:46]; // @[primitives.scala 104:54]
  wire  _T_99 = |notCDom_absSigSum[49:48]; // @[primitives.scala 104:54]
  wire  _T_101 = |notCDom_absSigSum[50]; // @[primitives.scala 107:57]
  wire [5:0] lo_lo = {_T_61,_T_59,_T_57,_T_55,_T_53,_T_51}; // @[primitives.scala 108:20]
  wire [12:0] lo_8 = {_T_75,_T_73,_T_71,_T_69,_T_67,_T_65,_T_63,lo_lo}; // @[primitives.scala 108:20]
  wire [5:0] hi_lo_3 = {_T_87,_T_85,_T_83,_T_81,_T_79,_T_77}; // @[primitives.scala 108:20]
  wire [25:0] notCDom_reduced2AbsSigSum = {_T_101,_T_99,_T_97,_T_95,_T_93,_T_91,_T_89,hi_lo_3,lo_8}; // @[primitives.scala 108:20]
  wire [4:0] _T_128 = notCDom_reduced2AbsSigSum[1] ? 5'h18 : 5'h19; // @[Mux.scala 47:69]
  wire [4:0] _T_129 = notCDom_reduced2AbsSigSum[2] ? 5'h17 : _T_128; // @[Mux.scala 47:69]
  wire [4:0] _T_130 = notCDom_reduced2AbsSigSum[3] ? 5'h16 : _T_129; // @[Mux.scala 47:69]
  wire [4:0] _T_131 = notCDom_reduced2AbsSigSum[4] ? 5'h15 : _T_130; // @[Mux.scala 47:69]
  wire [4:0] _T_132 = notCDom_reduced2AbsSigSum[5] ? 5'h14 : _T_131; // @[Mux.scala 47:69]
  wire [4:0] _T_133 = notCDom_reduced2AbsSigSum[6] ? 5'h13 : _T_132; // @[Mux.scala 47:69]
  wire [4:0] _T_134 = notCDom_reduced2AbsSigSum[7] ? 5'h12 : _T_133; // @[Mux.scala 47:69]
  wire [4:0] _T_135 = notCDom_reduced2AbsSigSum[8] ? 5'h11 : _T_134; // @[Mux.scala 47:69]
  wire [4:0] _T_136 = notCDom_reduced2AbsSigSum[9] ? 5'h10 : _T_135; // @[Mux.scala 47:69]
  wire [4:0] _T_137 = notCDom_reduced2AbsSigSum[10] ? 5'hf : _T_136; // @[Mux.scala 47:69]
  wire [4:0] _T_138 = notCDom_reduced2AbsSigSum[11] ? 5'he : _T_137; // @[Mux.scala 47:69]
  wire [4:0] _T_139 = notCDom_reduced2AbsSigSum[12] ? 5'hd : _T_138; // @[Mux.scala 47:69]
  wire [4:0] _T_140 = notCDom_reduced2AbsSigSum[13] ? 5'hc : _T_139; // @[Mux.scala 47:69]
  wire [4:0] _T_141 = notCDom_reduced2AbsSigSum[14] ? 5'hb : _T_140; // @[Mux.scala 47:69]
  wire [4:0] _T_142 = notCDom_reduced2AbsSigSum[15] ? 5'ha : _T_141; // @[Mux.scala 47:69]
  wire [4:0] _T_143 = notCDom_reduced2AbsSigSum[16] ? 5'h9 : _T_142; // @[Mux.scala 47:69]
  wire [4:0] _T_144 = notCDom_reduced2AbsSigSum[17] ? 5'h8 : _T_143; // @[Mux.scala 47:69]
  wire [4:0] _T_145 = notCDom_reduced2AbsSigSum[18] ? 5'h7 : _T_144; // @[Mux.scala 47:69]
  wire [4:0] _T_146 = notCDom_reduced2AbsSigSum[19] ? 5'h6 : _T_145; // @[Mux.scala 47:69]
  wire [4:0] _T_147 = notCDom_reduced2AbsSigSum[20] ? 5'h5 : _T_146; // @[Mux.scala 47:69]
  wire [4:0] _T_148 = notCDom_reduced2AbsSigSum[21] ? 5'h4 : _T_147; // @[Mux.scala 47:69]
  wire [4:0] _T_149 = notCDom_reduced2AbsSigSum[22] ? 5'h3 : _T_148; // @[Mux.scala 47:69]
  wire [4:0] _T_150 = notCDom_reduced2AbsSigSum[23] ? 5'h2 : _T_149; // @[Mux.scala 47:69]
  wire [4:0] _T_151 = notCDom_reduced2AbsSigSum[24] ? 5'h1 : _T_150; // @[Mux.scala 47:69]
  wire [4:0] notCDom_normDistReduced2 = notCDom_reduced2AbsSigSum[25] ? 5'h0 : _T_151; // @[Mux.scala 47:69]
  wire [5:0] notCDom_nearNormDist = {notCDom_normDistReduced2, 1'h0}; // @[MulAddRecFN.scala 242:56]
  wire [6:0] _T_152 = {1'b0,$signed(notCDom_nearNormDist)}; // @[MulAddRecFN.scala 243:69]
  wire [9:0] _GEN_4 = {{3{_T_152[6]}},_T_152}; // @[MulAddRecFN.scala 243:46]
  wire [9:0] notCDom_sExp = $signed(io_fromPreMul_sExpSum) - $signed(_GEN_4); // @[MulAddRecFN.scala 243:46]
  wire [113:0] _GEN_5 = {{63'd0}, notCDom_absSigSum}; // @[MulAddRecFN.scala 245:27]
  wire [113:0] _T_155 = _GEN_5 << notCDom_nearNormDist; // @[MulAddRecFN.scala 245:27]
  wire [28:0] notCDom_mainSig = _T_155[51:23]; // @[MulAddRecFN.scala 245:50]
  wire  _T_159 = |notCDom_reduced2AbsSigSum[1:0]; // @[primitives.scala 104:54]
  wire  _T_161 = |notCDom_reduced2AbsSigSum[3:2]; // @[primitives.scala 104:54]
  wire  _T_163 = |notCDom_reduced2AbsSigSum[5:4]; // @[primitives.scala 104:54]
  wire  _T_165 = |notCDom_reduced2AbsSigSum[7:6]; // @[primitives.scala 104:54]
  wire  _T_167 = |notCDom_reduced2AbsSigSum[9:8]; // @[primitives.scala 104:54]
  wire  _T_169 = |notCDom_reduced2AbsSigSum[11:10]; // @[primitives.scala 104:54]
  wire  _T_171 = |notCDom_reduced2AbsSigSum[12]; // @[primitives.scala 107:57]
  wire [6:0] _T_172 = {_T_171,_T_169,_T_167,_T_165,_T_163,_T_161,_T_159}; // @[primitives.scala 108:20]
  wire [3:0] _T_174 = ~notCDom_normDistReduced2[4:1]; // @[primitives.scala 51:21]
  wire [16:0] _T_175 = 17'sh10000 >>> _T_174; // @[primitives.scala 77:58]
  wire  hi_11 = _T_175[1]; // @[Bitwise.scala 109:18]
  wire  lo_10 = _T_175[2]; // @[Bitwise.scala 109:44]
  wire  hi_13 = _T_175[3]; // @[Bitwise.scala 109:18]
  wire  lo_11 = _T_175[4]; // @[Bitwise.scala 109:44]
  wire  hi_15 = _T_175[5]; // @[Bitwise.scala 109:18]
  wire  lo_13 = _T_175[6]; // @[Bitwise.scala 109:44]
  wire [5:0] _T_181 = {hi_11,lo_10,hi_13,lo_11,hi_15,lo_13}; // @[Cat.scala 30:58]
  wire [6:0] _GEN_6 = {{1'd0}, _T_181}; // @[MulAddRecFN.scala 249:78]
  wire [6:0] _T_182 = _T_172 & _GEN_6; // @[MulAddRecFN.scala 249:78]
  wire  notCDom_reduced4SigExtra = |_T_182; // @[MulAddRecFN.scala 251:11]
  wire [25:0] hi_16 = notCDom_mainSig[28:3]; // @[MulAddRecFN.scala 253:28]
  wire  lo_15 = |notCDom_mainSig[2:0] | notCDom_reduced4SigExtra; // @[MulAddRecFN.scala 254:39]
  wire [26:0] notCDom_sig = {hi_16,lo_15}; // @[Cat.scala 30:58]
  wire  notCDom_completeCancellation = notCDom_sig[26:25] == 2'h0; // @[MulAddRecFN.scala 257:50]
  wire  _T_186 = io_fromPreMul_signProd ^ notCDom_signSigSum; // @[MulAddRecFN.scala 261:36]
  wire  notCDom_sign = notCDom_completeCancellation ? 1'h0 : _T_186; // @[MulAddRecFN.scala 259:12]
  wire  notNaN_isInfProd = io_fromPreMul_isInfA | io_fromPreMul_isInfB; // @[MulAddRecFN.scala 266:49]
  wire  notNaN_isInfOut = notNaN_isInfProd | io_fromPreMul_isInfC; // @[MulAddRecFN.scala 267:44]
  wire  notNaN_addZeros = (io_fromPreMul_isZeroA | io_fromPreMul_isZeroB) & io_fromPreMul_isZeroC; // @[MulAddRecFN.scala 269:58]
  wire  _T_188 = io_fromPreMul_isInfA & io_fromPreMul_isZeroB; // @[MulAddRecFN.scala 274:31]
  wire  _T_189 = io_fromPreMul_isSigNaNAny | _T_188; // @[MulAddRecFN.scala 273:35]
  wire  _T_190 = io_fromPreMul_isZeroA & io_fromPreMul_isInfB; // @[MulAddRecFN.scala 275:32]
  wire  _T_191 = _T_189 | _T_190; // @[MulAddRecFN.scala 274:57]
  wire  _T_194 = ~io_fromPreMul_isNaNAOrB & notNaN_isInfProd; // @[MulAddRecFN.scala 276:36]
  wire  _T_195 = _T_194 & io_fromPreMul_isInfC; // @[MulAddRecFN.scala 277:61]
  wire  _T_196 = _T_195 & io_fromPreMul_doSubMags; // @[MulAddRecFN.scala 278:35]
  wire  _T_200 = ~io_fromPreMul_CIsDominant & notCDom_completeCancellation; // @[MulAddRecFN.scala 285:42]
  wire  _T_203 = io_fromPreMul_isInfC & CDom_sign; // @[MulAddRecFN.scala 288:31]
  wire  _T_204 = notNaN_isInfProd & io_fromPreMul_signProd | _T_203; // @[MulAddRecFN.scala 287:54]
  wire  _T_207 = notNaN_addZeros & io_fromPreMul_signProd; // @[MulAddRecFN.scala 289:48]
  wire  _T_208 = _T_207 & CDom_sign; // @[MulAddRecFN.scala 290:36]
  wire  _T_209 = _T_204 | _T_208; // @[MulAddRecFN.scala 288:43]
  wire  _T_217 = io_fromPreMul_CIsDominant ? CDom_sign : notCDom_sign; // @[MulAddRecFN.scala 294:17]
  wire  _T_218 = ~notNaN_isInfOut & ~notNaN_addZeros & _T_217; // @[MulAddRecFN.scala 293:49]
  assign io_invalidExc = _T_191 | _T_196; // @[MulAddRecFN.scala 275:57]
  assign io_rawOut_isNaN = io_fromPreMul_isNaNAOrB | io_fromPreMul_isNaNC; // @[MulAddRecFN.scala 280:48]
  assign io_rawOut_isInf = notNaN_isInfProd | io_fromPreMul_isInfC; // @[MulAddRecFN.scala 267:44]
  assign io_rawOut_isZero = notNaN_addZeros | _T_200; // @[MulAddRecFN.scala 284:25]
  assign io_rawOut_sign = _T_209 | _T_218; // @[MulAddRecFN.scala 292:50]
  assign io_rawOut_sExp = io_fromPreMul_CIsDominant ? $signed(CDom_sExp) : $signed(notCDom_sExp); // @[MulAddRecFN.scala 295:26]
  assign io_rawOut_sig = io_fromPreMul_CIsDominant ? CDom_sig : notCDom_sig; // @[MulAddRecFN.scala 296:25]
endmodule
module RoundAnyRawFNToRecFN(
  input         io_invalidExc,
  input         io_in_isNaN,
  input         io_in_isInf,
  input         io_in_isZero,
  input         io_in_sign,
  input  [9:0]  io_in_sExp,
  input  [26:0] io_in_sig,
  output [32:0] io_out
);
  wire  doShiftSigDown1 = io_in_sig[26]; // @[RoundAnyRawFNToRecFN.scala 118:61]
  wire [8:0] _T_4 = ~io_in_sExp[8:0]; // @[primitives.scala 51:21]
  wire [64:0] _T_11 = 65'sh10000000000000000 >>> _T_4[5:0]; // @[primitives.scala 77:58]
  wire [15:0] _T_17 = {{8'd0}, _T_11[57:50]}; // @[Bitwise.scala 103:31]
  wire [15:0] _T_19 = {_T_11[49:42], 8'h0}; // @[Bitwise.scala 103:65]
  wire [15:0] _T_21 = _T_19 & 16'hff00; // @[Bitwise.scala 103:75]
  wire [15:0] _T_22 = _T_17 | _T_21; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_0 = {{4'd0}, _T_22[15:4]}; // @[Bitwise.scala 103:31]
  wire [15:0] _T_27 = _GEN_0 & 16'hf0f; // @[Bitwise.scala 103:31]
  wire [15:0] _T_29 = {_T_22[11:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [15:0] _T_31 = _T_29 & 16'hf0f0; // @[Bitwise.scala 103:75]
  wire [15:0] _T_32 = _T_27 | _T_31; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_1 = {{2'd0}, _T_32[15:2]}; // @[Bitwise.scala 103:31]
  wire [15:0] _T_37 = _GEN_1 & 16'h3333; // @[Bitwise.scala 103:31]
  wire [15:0] _T_39 = {_T_32[13:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [15:0] _T_41 = _T_39 & 16'hcccc; // @[Bitwise.scala 103:75]
  wire [15:0] _T_42 = _T_37 | _T_41; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_2 = {{1'd0}, _T_42[15:1]}; // @[Bitwise.scala 103:31]
  wire [15:0] _T_47 = _GEN_2 & 16'h5555; // @[Bitwise.scala 103:31]
  wire [15:0] _T_49 = {_T_42[14:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [15:0] _T_51 = _T_49 & 16'haaaa; // @[Bitwise.scala 103:75]
  wire [15:0] hi = _T_47 | _T_51; // @[Bitwise.scala 103:39]
  wire  hi_1 = _T_11[58]; // @[Bitwise.scala 109:18]
  wire  lo = _T_11[59]; // @[Bitwise.scala 109:44]
  wire  hi_3 = _T_11[60]; // @[Bitwise.scala 109:18]
  wire  lo_1 = _T_11[61]; // @[Bitwise.scala 109:44]
  wire  hi_5 = _T_11[62]; // @[Bitwise.scala 109:18]
  wire  lo_3 = _T_11[63]; // @[Bitwise.scala 109:44]
  wire [21:0] _T_57 = {hi,hi_1,lo,hi_3,lo_1,hi_5,lo_3}; // @[Cat.scala 30:58]
  wire [21:0] _T_58 = ~_T_57; // @[primitives.scala 74:36]
  wire [21:0] _T_59 = _T_4[6] ? 22'h0 : _T_58; // @[primitives.scala 74:21]
  wire [21:0] hi_6 = ~_T_59; // @[primitives.scala 74:17]
  wire [24:0] _T_60 = {hi_6,3'h7}; // @[Cat.scala 30:58]
  wire  hi_7 = _T_11[0]; // @[Bitwise.scala 109:18]
  wire  lo_6 = _T_11[1]; // @[Bitwise.scala 109:44]
  wire  lo_7 = _T_11[2]; // @[Bitwise.scala 109:44]
  wire [2:0] _T_66 = {hi_7,lo_6,lo_7}; // @[Cat.scala 30:58]
  wire [2:0] _T_67 = _T_4[6] ? _T_66 : 3'h0; // @[primitives.scala 61:24]
  wire [24:0] _T_68 = _T_4[7] ? _T_60 : {{22'd0}, _T_67}; // @[primitives.scala 66:24]
  wire [24:0] _T_69 = _T_4[8] ? _T_68 : 25'h0; // @[primitives.scala 61:24]
  wire [24:0] _GEN_3 = {{24'd0}, doShiftSigDown1}; // @[RoundAnyRawFNToRecFN.scala 157:23]
  wire [24:0] hi_9 = _T_69 | _GEN_3; // @[RoundAnyRawFNToRecFN.scala 157:23]
  wire [26:0] _T_70 = {hi_9,2'h3}; // @[Cat.scala 30:58]
  wire [25:0] lo_8 = _T_70[26:1]; // @[RoundAnyRawFNToRecFN.scala 160:57]
  wire [26:0] _T_71 = {1'h0,lo_8}; // @[Cat.scala 30:58]
  wire [26:0] _T_72 = ~_T_71; // @[RoundAnyRawFNToRecFN.scala 161:28]
  wire [26:0] _T_73 = _T_72 & _T_70; // @[RoundAnyRawFNToRecFN.scala 161:46]
  wire [26:0] _T_74 = io_in_sig & _T_73; // @[RoundAnyRawFNToRecFN.scala 162:40]
  wire  _T_75 = |_T_74; // @[RoundAnyRawFNToRecFN.scala 162:56]
  wire [26:0] _T_76 = io_in_sig & _T_71; // @[RoundAnyRawFNToRecFN.scala 163:42]
  wire  _T_77 = |_T_76; // @[RoundAnyRawFNToRecFN.scala 163:62]
  wire [26:0] _T_83 = io_in_sig | _T_70; // @[RoundAnyRawFNToRecFN.scala 172:32]
  wire [25:0] _T_85 = _T_83[26:2] + 25'h1; // @[RoundAnyRawFNToRecFN.scala 172:49]
  wire  _T_87 = ~_T_77; // @[RoundAnyRawFNToRecFN.scala 174:30]
  wire [25:0] _T_90 = _T_75 & _T_87 ? lo_8 : 26'h0; // @[RoundAnyRawFNToRecFN.scala 173:25]
  wire [25:0] _T_91 = ~_T_90; // @[RoundAnyRawFNToRecFN.scala 173:21]
  wire [25:0] _T_92 = _T_85 & _T_91; // @[RoundAnyRawFNToRecFN.scala 172:61]
  wire [26:0] _T_93 = ~_T_70; // @[RoundAnyRawFNToRecFN.scala 178:32]
  wire [26:0] _T_94 = io_in_sig & _T_93; // @[RoundAnyRawFNToRecFN.scala 178:30]
  wire [25:0] _T_99 = {{1'd0}, _T_94[26:2]}; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [25:0] _T_100 = _T_75 ? _T_92 : _T_99; // @[RoundAnyRawFNToRecFN.scala 171:16]
  wire [2:0] _T_102 = {1'b0,$signed(_T_100[25:24])}; // @[RoundAnyRawFNToRecFN.scala 183:69]
  wire [9:0] _GEN_4 = {{7{_T_102[2]}},_T_102}; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [10:0] _T_103 = $signed(io_in_sExp) + $signed(_GEN_4); // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [8:0] common_expOut = _T_103[8:0]; // @[RoundAnyRawFNToRecFN.scala 185:37]
  wire [22:0] common_fractOut = doShiftSigDown1 ? _T_100[23:1] : _T_100[22:0]; // @[RoundAnyRawFNToRecFN.scala 187:16]
  wire [3:0] _T_108 = _T_103[10:7]; // @[RoundAnyRawFNToRecFN.scala 194:30]
  wire  common_overflow = $signed(_T_108) >= 4'sh3; // @[RoundAnyRawFNToRecFN.scala 194:50]
  wire  common_totalUnderflow = $signed(_T_103) < 11'sh6b; // @[RoundAnyRawFNToRecFN.scala 198:31]
  wire  isNaNOut = io_invalidExc | io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 233:34]
  wire  commonCase = ~isNaNOut & ~io_in_isInf & ~io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 235:61]
  wire  overflow = commonCase & common_overflow; // @[RoundAnyRawFNToRecFN.scala 236:32]
  wire  notNaN_isInfOut = io_in_isInf | overflow; // @[RoundAnyRawFNToRecFN.scala 246:32]
  wire  signOut = isNaNOut ? 1'h0 : io_in_sign; // @[RoundAnyRawFNToRecFN.scala 248:22]
  wire [8:0] _T_157 = io_in_isZero | common_totalUnderflow ? 9'h1c0 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 251:18]
  wire [8:0] _T_158 = ~_T_157; // @[RoundAnyRawFNToRecFN.scala 251:14]
  wire [8:0] _T_159 = common_expOut & _T_158; // @[RoundAnyRawFNToRecFN.scala 250:24]
  wire [8:0] _T_167 = notNaN_isInfOut ? 9'h40 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 263:18]
  wire [8:0] _T_168 = ~_T_167; // @[RoundAnyRawFNToRecFN.scala 263:14]
  wire [8:0] _T_169 = _T_159 & _T_168; // @[RoundAnyRawFNToRecFN.scala 262:17]
  wire [8:0] _T_174 = notNaN_isInfOut ? 9'h180 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 275:16]
  wire [8:0] _T_175 = _T_169 | _T_174; // @[RoundAnyRawFNToRecFN.scala 274:15]
  wire [8:0] _T_176 = isNaNOut ? 9'h1c0 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 276:16]
  wire [8:0] expOut = _T_175 | _T_176; // @[RoundAnyRawFNToRecFN.scala 275:77]
  wire [22:0] _T_179 = isNaNOut ? 23'h400000 : 23'h0; // @[RoundAnyRawFNToRecFN.scala 279:16]
  wire [22:0] fractOut = isNaNOut | io_in_isZero | common_totalUnderflow ? _T_179 : common_fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12]
  wire [9:0] hi_10 = {signOut,expOut}; // @[Cat.scala 30:58]
  assign io_out = {hi_10,fractOut}; // @[Cat.scala 30:58]
endmodule
module RoundRawFNToRecFN(
  input         io_invalidExc,
  input         io_in_isNaN,
  input         io_in_isInf,
  input         io_in_isZero,
  input         io_in_sign,
  input  [9:0]  io_in_sExp,
  input  [26:0] io_in_sig,
  output [32:0] io_out
);
  wire  roundAnyRawFNToRecFN_io_invalidExc; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_sign; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [9:0] roundAnyRawFNToRecFN_io_in_sExp; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [26:0] roundAnyRawFNToRecFN_io_in_sig; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [32:0] roundAnyRawFNToRecFN_io_out; // @[RoundAnyRawFNToRecFN.scala 307:15]
  RoundAnyRawFNToRecFN roundAnyRawFNToRecFN ( // @[RoundAnyRawFNToRecFN.scala 307:15]
    .io_invalidExc(roundAnyRawFNToRecFN_io_invalidExc),
    .io_in_isNaN(roundAnyRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundAnyRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundAnyRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundAnyRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundAnyRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundAnyRawFNToRecFN_io_in_sig),
    .io_out(roundAnyRawFNToRecFN_io_out)
  );
  assign io_out = roundAnyRawFNToRecFN_io_out; // @[RoundAnyRawFNToRecFN.scala 315:23]
  assign roundAnyRawFNToRecFN_io_invalidExc = io_invalidExc; // @[RoundAnyRawFNToRecFN.scala 310:44]
  assign roundAnyRawFNToRecFN_io_in_isNaN = io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_isInf = io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_isZero = io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_sign = io_in_sign; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_sExp = io_in_sExp; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_sig = io_in_sig; // @[RoundAnyRawFNToRecFN.scala 312:44]
endmodule
module MY_MULADD(
  input         clock,
  input         reset,
  input  [31:0] io_a,
  input  [31:0] io_b,
  input  [31:0] io_c,
  output [31:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_REG_INIT
  wire [32:0] mulAddRecFNToRaw_preMul_io_a; // @[FMULADD_1G_2.scala 36:15]
  wire [32:0] mulAddRecFNToRaw_preMul_io_b; // @[FMULADD_1G_2.scala 36:15]
  wire [32:0] mulAddRecFNToRaw_preMul_io_c; // @[FMULADD_1G_2.scala 36:15]
  wire [23:0] mulAddRecFNToRaw_preMul_io_mulAddA; // @[FMULADD_1G_2.scala 36:15]
  wire [23:0] mulAddRecFNToRaw_preMul_io_mulAddB; // @[FMULADD_1G_2.scala 36:15]
  wire [47:0] mulAddRecFNToRaw_preMul_io_mulAddC; // @[FMULADD_1G_2.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny; // @[FMULADD_1G_2.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB; // @[FMULADD_1G_2.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfA; // @[FMULADD_1G_2.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA; // @[FMULADD_1G_2.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfB; // @[FMULADD_1G_2.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB; // @[FMULADD_1G_2.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_signProd; // @[FMULADD_1G_2.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC; // @[FMULADD_1G_2.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfC; // @[FMULADD_1G_2.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC; // @[FMULADD_1G_2.scala 36:15]
  wire [9:0] mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum; // @[FMULADD_1G_2.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags; // @[FMULADD_1G_2.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant; // @[FMULADD_1G_2.scala 36:15]
  wire [4:0] mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist; // @[FMULADD_1G_2.scala 36:15]
  wire [25:0] mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC; // @[FMULADD_1G_2.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC; // @[FMULADD_1G_2.scala 36:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny; // @[FMULADD_1G_2.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB; // @[FMULADD_1G_2.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA; // @[FMULADD_1G_2.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA; // @[FMULADD_1G_2.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB; // @[FMULADD_1G_2.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB; // @[FMULADD_1G_2.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_signProd; // @[FMULADD_1G_2.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC; // @[FMULADD_1G_2.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC; // @[FMULADD_1G_2.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC; // @[FMULADD_1G_2.scala 116:15]
  wire [9:0] mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum; // @[FMULADD_1G_2.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags; // @[FMULADD_1G_2.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant; // @[FMULADD_1G_2.scala 116:15]
  wire [4:0] mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist; // @[FMULADD_1G_2.scala 116:15]
  wire [25:0] mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC; // @[FMULADD_1G_2.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC; // @[FMULADD_1G_2.scala 116:15]
  wire [48:0] mulAddRecFNToRaw_postMul_io_mulAddResult; // @[FMULADD_1G_2.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_invalidExc; // @[FMULADD_1G_2.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isNaN; // @[FMULADD_1G_2.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isInf; // @[FMULADD_1G_2.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isZero; // @[FMULADD_1G_2.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_sign; // @[FMULADD_1G_2.scala 116:15]
  wire [9:0] mulAddRecFNToRaw_postMul_io_rawOut_sExp; // @[FMULADD_1G_2.scala 116:15]
  wire [26:0] mulAddRecFNToRaw_postMul_io_rawOut_sig; // @[FMULADD_1G_2.scala 116:15]
  wire  roundRawFNToRecFN_io_invalidExc; // @[FMULADD_1G_2.scala 137:15]
  wire  roundRawFNToRecFN_io_in_isNaN; // @[FMULADD_1G_2.scala 137:15]
  wire  roundRawFNToRecFN_io_in_isInf; // @[FMULADD_1G_2.scala 137:15]
  wire  roundRawFNToRecFN_io_in_isZero; // @[FMULADD_1G_2.scala 137:15]
  wire  roundRawFNToRecFN_io_in_sign; // @[FMULADD_1G_2.scala 137:15]
  wire [9:0] roundRawFNToRecFN_io_in_sExp; // @[FMULADD_1G_2.scala 137:15]
  wire [26:0] roundRawFNToRecFN_io_in_sig; // @[FMULADD_1G_2.scala 137:15]
  wire [32:0] roundRawFNToRecFN_io_out; // @[FMULADD_1G_2.scala 137:15]
  reg [23:0] premul_a; // @[FMULADD_1G_2.scala 15:37]
  reg [23:0] premul_b; // @[FMULADD_1G_2.scala 16:37]
  reg [47:0] premul_c; // @[FMULADD_1G_2.scala 17:37]
  reg  isSigNaNAny; // @[FMULADD_1G_2.scala 18:33]
  reg  isNaNAOrB; // @[FMULADD_1G_2.scala 19:34]
  reg  isInfA; // @[FMULADD_1G_2.scala 20:43]
  reg  isZeroA; // @[FMULADD_1G_2.scala 21:40]
  reg  isInfB; // @[FMULADD_1G_2.scala 22:43]
  reg  isZeroB; // @[FMULADD_1G_2.scala 23:40]
  reg  signProd; // @[FMULADD_1G_2.scala 24:38]
  reg  isNaNC; // @[FMULADD_1G_2.scala 25:39]
  reg  isInfC; // @[FMULADD_1G_2.scala 26:42]
  reg  isZeroC; // @[FMULADD_1G_2.scala 27:39]
  reg [9:0] sExpSum; // @[FMULADD_1G_2.scala 28:36]
  reg  doSubMags; // @[FMULADD_1G_2.scala 29:33]
  reg  CIsDominant; // @[FMULADD_1G_2.scala 30:33]
  reg [4:0] CDom_CAlignDist; // @[FMULADD_1G_2.scala 31:34]
  reg [25:0] highAlignedSigC; // @[FMULADD_1G_2.scala 32:37]
  reg  bit0AlignedSigC; // @[FMULADD_1G_2.scala 33:38]
  wire  _T_3 = io_a[30:23] == 8'h0; // @[rawFloatFromFN.scala 50:34]
  wire  _T_4 = io_a[22:0] == 23'h0; // @[rawFloatFromFN.scala 51:38]
  wire [4:0] _T_28 = io_a[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:69]
  wire [4:0] _T_29 = io_a[2] ? 5'h14 : _T_28; // @[Mux.scala 47:69]
  wire [4:0] _T_30 = io_a[3] ? 5'h13 : _T_29; // @[Mux.scala 47:69]
  wire [4:0] _T_31 = io_a[4] ? 5'h12 : _T_30; // @[Mux.scala 47:69]
  wire [4:0] _T_32 = io_a[5] ? 5'h11 : _T_31; // @[Mux.scala 47:69]
  wire [4:0] _T_33 = io_a[6] ? 5'h10 : _T_32; // @[Mux.scala 47:69]
  wire [4:0] _T_34 = io_a[7] ? 5'hf : _T_33; // @[Mux.scala 47:69]
  wire [4:0] _T_35 = io_a[8] ? 5'he : _T_34; // @[Mux.scala 47:69]
  wire [4:0] _T_36 = io_a[9] ? 5'hd : _T_35; // @[Mux.scala 47:69]
  wire [4:0] _T_37 = io_a[10] ? 5'hc : _T_36; // @[Mux.scala 47:69]
  wire [4:0] _T_38 = io_a[11] ? 5'hb : _T_37; // @[Mux.scala 47:69]
  wire [4:0] _T_39 = io_a[12] ? 5'ha : _T_38; // @[Mux.scala 47:69]
  wire [4:0] _T_40 = io_a[13] ? 5'h9 : _T_39; // @[Mux.scala 47:69]
  wire [4:0] _T_41 = io_a[14] ? 5'h8 : _T_40; // @[Mux.scala 47:69]
  wire [4:0] _T_42 = io_a[15] ? 5'h7 : _T_41; // @[Mux.scala 47:69]
  wire [4:0] _T_43 = io_a[16] ? 5'h6 : _T_42; // @[Mux.scala 47:69]
  wire [4:0] _T_44 = io_a[17] ? 5'h5 : _T_43; // @[Mux.scala 47:69]
  wire [4:0] _T_45 = io_a[18] ? 5'h4 : _T_44; // @[Mux.scala 47:69]
  wire [4:0] _T_46 = io_a[19] ? 5'h3 : _T_45; // @[Mux.scala 47:69]
  wire [4:0] _T_47 = io_a[20] ? 5'h2 : _T_46; // @[Mux.scala 47:69]
  wire [4:0] _T_48 = io_a[21] ? 5'h1 : _T_47; // @[Mux.scala 47:69]
  wire [4:0] _T_49 = io_a[22] ? 5'h0 : _T_48; // @[Mux.scala 47:69]
  wire [53:0] _GEN_0 = {{31'd0}, io_a[22:0]}; // @[rawFloatFromFN.scala 54:36]
  wire [53:0] _T_50 = _GEN_0 << _T_49; // @[rawFloatFromFN.scala 54:36]
  wire [22:0] _T_52 = {_T_50[21:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  wire [8:0] _GEN_1 = {{4'd0}, _T_49}; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_53 = _GEN_1 ^ 9'h1ff; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_54 = _T_3 ? _T_53 : {{1'd0}, io_a[30:23]}; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_55 = _T_3 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  wire [7:0] _GEN_2 = {{6'd0}, _T_55}; // @[rawFloatFromFN.scala 60:22]
  wire [7:0] _T_56 = 8'h80 | _GEN_2; // @[rawFloatFromFN.scala 60:22]
  wire [8:0] _GEN_3 = {{1'd0}, _T_56}; // @[rawFloatFromFN.scala 59:15]
  wire [8:0] _T_58 = _T_54 + _GEN_3; // @[rawFloatFromFN.scala 59:15]
  wire  _T_59 = _T_3 & _T_4; // @[rawFloatFromFN.scala 62:34]
  wire  _T_61 = _T_58[8:7] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  wire  _T_63 = _T_61 & ~_T_4; // @[rawFloatFromFN.scala 66:33]
  wire [9:0] _T_66 = {1'b0,$signed(_T_58)}; // @[rawFloatFromFN.scala 70:48]
  wire  hi_lo = ~_T_59; // @[rawFloatFromFN.scala 72:29]
  wire [22:0] lo = _T_3 ? _T_52 : io_a[22:0]; // @[rawFloatFromFN.scala 72:42]
  wire [24:0] _T_67 = {1'h0,hi_lo,lo}; // @[Cat.scala 30:58]
  wire [2:0] _T_69 = _T_59 ? 3'h0 : _T_66[8:6]; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_4 = {{2'd0}, _T_63}; // @[recFNFromFN.scala 48:79]
  wire [2:0] hi_lo_1 = _T_69 | _GEN_4; // @[recFNFromFN.scala 48:79]
  wire [5:0] lo_hi = _T_66[5:0]; // @[recFNFromFN.scala 50:23]
  wire [22:0] lo_lo = _T_67[22:0]; // @[recFNFromFN.scala 51:22]
  wire [28:0] lo_1 = {lo_hi,lo_lo}; // @[Cat.scala 30:58]
  wire [3:0] hi_1 = {io_a[31],hi_lo_1}; // @[Cat.scala 30:58]
  wire  _T_75 = io_b[30:23] == 8'h0; // @[rawFloatFromFN.scala 50:34]
  wire  _T_76 = io_b[22:0] == 23'h0; // @[rawFloatFromFN.scala 51:38]
  wire [4:0] _T_100 = io_b[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:69]
  wire [4:0] _T_101 = io_b[2] ? 5'h14 : _T_100; // @[Mux.scala 47:69]
  wire [4:0] _T_102 = io_b[3] ? 5'h13 : _T_101; // @[Mux.scala 47:69]
  wire [4:0] _T_103 = io_b[4] ? 5'h12 : _T_102; // @[Mux.scala 47:69]
  wire [4:0] _T_104 = io_b[5] ? 5'h11 : _T_103; // @[Mux.scala 47:69]
  wire [4:0] _T_105 = io_b[6] ? 5'h10 : _T_104; // @[Mux.scala 47:69]
  wire [4:0] _T_106 = io_b[7] ? 5'hf : _T_105; // @[Mux.scala 47:69]
  wire [4:0] _T_107 = io_b[8] ? 5'he : _T_106; // @[Mux.scala 47:69]
  wire [4:0] _T_108 = io_b[9] ? 5'hd : _T_107; // @[Mux.scala 47:69]
  wire [4:0] _T_109 = io_b[10] ? 5'hc : _T_108; // @[Mux.scala 47:69]
  wire [4:0] _T_110 = io_b[11] ? 5'hb : _T_109; // @[Mux.scala 47:69]
  wire [4:0] _T_111 = io_b[12] ? 5'ha : _T_110; // @[Mux.scala 47:69]
  wire [4:0] _T_112 = io_b[13] ? 5'h9 : _T_111; // @[Mux.scala 47:69]
  wire [4:0] _T_113 = io_b[14] ? 5'h8 : _T_112; // @[Mux.scala 47:69]
  wire [4:0] _T_114 = io_b[15] ? 5'h7 : _T_113; // @[Mux.scala 47:69]
  wire [4:0] _T_115 = io_b[16] ? 5'h6 : _T_114; // @[Mux.scala 47:69]
  wire [4:0] _T_116 = io_b[17] ? 5'h5 : _T_115; // @[Mux.scala 47:69]
  wire [4:0] _T_117 = io_b[18] ? 5'h4 : _T_116; // @[Mux.scala 47:69]
  wire [4:0] _T_118 = io_b[19] ? 5'h3 : _T_117; // @[Mux.scala 47:69]
  wire [4:0] _T_119 = io_b[20] ? 5'h2 : _T_118; // @[Mux.scala 47:69]
  wire [4:0] _T_120 = io_b[21] ? 5'h1 : _T_119; // @[Mux.scala 47:69]
  wire [4:0] _T_121 = io_b[22] ? 5'h0 : _T_120; // @[Mux.scala 47:69]
  wire [53:0] _GEN_5 = {{31'd0}, io_b[22:0]}; // @[rawFloatFromFN.scala 54:36]
  wire [53:0] _T_122 = _GEN_5 << _T_121; // @[rawFloatFromFN.scala 54:36]
  wire [22:0] _T_124 = {_T_122[21:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  wire [8:0] _GEN_6 = {{4'd0}, _T_121}; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_125 = _GEN_6 ^ 9'h1ff; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_126 = _T_75 ? _T_125 : {{1'd0}, io_b[30:23]}; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_127 = _T_75 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  wire [7:0] _GEN_7 = {{6'd0}, _T_127}; // @[rawFloatFromFN.scala 60:22]
  wire [7:0] _T_128 = 8'h80 | _GEN_7; // @[rawFloatFromFN.scala 60:22]
  wire [8:0] _GEN_8 = {{1'd0}, _T_128}; // @[rawFloatFromFN.scala 59:15]
  wire [8:0] _T_130 = _T_126 + _GEN_8; // @[rawFloatFromFN.scala 59:15]
  wire  _T_131 = _T_75 & _T_76; // @[rawFloatFromFN.scala 62:34]
  wire  _T_133 = _T_130[8:7] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  wire  _T_135 = _T_133 & ~_T_76; // @[rawFloatFromFN.scala 66:33]
  wire [9:0] _T_138 = {1'b0,$signed(_T_130)}; // @[rawFloatFromFN.scala 70:48]
  wire  hi_lo_2 = ~_T_131; // @[rawFloatFromFN.scala 72:29]
  wire [22:0] lo_2 = _T_75 ? _T_124 : io_b[22:0]; // @[rawFloatFromFN.scala 72:42]
  wire [24:0] _T_139 = {1'h0,hi_lo_2,lo_2}; // @[Cat.scala 30:58]
  wire [2:0] _T_141 = _T_131 ? 3'h0 : _T_138[8:6]; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_9 = {{2'd0}, _T_135}; // @[recFNFromFN.scala 48:79]
  wire [2:0] hi_lo_3 = _T_141 | _GEN_9; // @[recFNFromFN.scala 48:79]
  wire [5:0] lo_hi_1 = _T_138[5:0]; // @[recFNFromFN.scala 50:23]
  wire [22:0] lo_lo_1 = _T_139[22:0]; // @[recFNFromFN.scala 51:22]
  wire [28:0] lo_3 = {lo_hi_1,lo_lo_1}; // @[Cat.scala 30:58]
  wire [3:0] hi_3 = {io_b[31],hi_lo_3}; // @[Cat.scala 30:58]
  wire  _T_147 = io_c[30:23] == 8'h0; // @[rawFloatFromFN.scala 50:34]
  wire  _T_148 = io_c[22:0] == 23'h0; // @[rawFloatFromFN.scala 51:38]
  wire [4:0] _T_172 = io_c[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:69]
  wire [4:0] _T_173 = io_c[2] ? 5'h14 : _T_172; // @[Mux.scala 47:69]
  wire [4:0] _T_174 = io_c[3] ? 5'h13 : _T_173; // @[Mux.scala 47:69]
  wire [4:0] _T_175 = io_c[4] ? 5'h12 : _T_174; // @[Mux.scala 47:69]
  wire [4:0] _T_176 = io_c[5] ? 5'h11 : _T_175; // @[Mux.scala 47:69]
  wire [4:0] _T_177 = io_c[6] ? 5'h10 : _T_176; // @[Mux.scala 47:69]
  wire [4:0] _T_178 = io_c[7] ? 5'hf : _T_177; // @[Mux.scala 47:69]
  wire [4:0] _T_179 = io_c[8] ? 5'he : _T_178; // @[Mux.scala 47:69]
  wire [4:0] _T_180 = io_c[9] ? 5'hd : _T_179; // @[Mux.scala 47:69]
  wire [4:0] _T_181 = io_c[10] ? 5'hc : _T_180; // @[Mux.scala 47:69]
  wire [4:0] _T_182 = io_c[11] ? 5'hb : _T_181; // @[Mux.scala 47:69]
  wire [4:0] _T_183 = io_c[12] ? 5'ha : _T_182; // @[Mux.scala 47:69]
  wire [4:0] _T_184 = io_c[13] ? 5'h9 : _T_183; // @[Mux.scala 47:69]
  wire [4:0] _T_185 = io_c[14] ? 5'h8 : _T_184; // @[Mux.scala 47:69]
  wire [4:0] _T_186 = io_c[15] ? 5'h7 : _T_185; // @[Mux.scala 47:69]
  wire [4:0] _T_187 = io_c[16] ? 5'h6 : _T_186; // @[Mux.scala 47:69]
  wire [4:0] _T_188 = io_c[17] ? 5'h5 : _T_187; // @[Mux.scala 47:69]
  wire [4:0] _T_189 = io_c[18] ? 5'h4 : _T_188; // @[Mux.scala 47:69]
  wire [4:0] _T_190 = io_c[19] ? 5'h3 : _T_189; // @[Mux.scala 47:69]
  wire [4:0] _T_191 = io_c[20] ? 5'h2 : _T_190; // @[Mux.scala 47:69]
  wire [4:0] _T_192 = io_c[21] ? 5'h1 : _T_191; // @[Mux.scala 47:69]
  wire [4:0] _T_193 = io_c[22] ? 5'h0 : _T_192; // @[Mux.scala 47:69]
  wire [53:0] _GEN_10 = {{31'd0}, io_c[22:0]}; // @[rawFloatFromFN.scala 54:36]
  wire [53:0] _T_194 = _GEN_10 << _T_193; // @[rawFloatFromFN.scala 54:36]
  wire [22:0] _T_196 = {_T_194[21:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  wire [8:0] _GEN_11 = {{4'd0}, _T_193}; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_197 = _GEN_11 ^ 9'h1ff; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_198 = _T_147 ? _T_197 : {{1'd0}, io_c[30:23]}; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_199 = _T_147 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  wire [7:0] _GEN_12 = {{6'd0}, _T_199}; // @[rawFloatFromFN.scala 60:22]
  wire [7:0] _T_200 = 8'h80 | _GEN_12; // @[rawFloatFromFN.scala 60:22]
  wire [8:0] _GEN_13 = {{1'd0}, _T_200}; // @[rawFloatFromFN.scala 59:15]
  wire [8:0] _T_202 = _T_198 + _GEN_13; // @[rawFloatFromFN.scala 59:15]
  wire  _T_203 = _T_147 & _T_148; // @[rawFloatFromFN.scala 62:34]
  wire  _T_205 = _T_202[8:7] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  wire  _T_207 = _T_205 & ~_T_148; // @[rawFloatFromFN.scala 66:33]
  wire [9:0] _T_210 = {1'b0,$signed(_T_202)}; // @[rawFloatFromFN.scala 70:48]
  wire  hi_lo_4 = ~_T_203; // @[rawFloatFromFN.scala 72:29]
  wire [22:0] lo_4 = _T_147 ? _T_196 : io_c[22:0]; // @[rawFloatFromFN.scala 72:42]
  wire [24:0] _T_211 = {1'h0,hi_lo_4,lo_4}; // @[Cat.scala 30:58]
  wire [2:0] _T_213 = _T_203 ? 3'h0 : _T_210[8:6]; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_14 = {{2'd0}, _T_207}; // @[recFNFromFN.scala 48:79]
  wire [2:0] hi_lo_5 = _T_213 | _GEN_14; // @[recFNFromFN.scala 48:79]
  wire [5:0] lo_hi_2 = _T_210[5:0]; // @[recFNFromFN.scala 50:23]
  wire [22:0] lo_lo_2 = _T_211[22:0]; // @[recFNFromFN.scala 51:22]
  wire [28:0] lo_5 = {lo_hi_2,lo_lo_2}; // @[Cat.scala 30:58]
  wire [3:0] hi_5 = {io_c[31],hi_lo_5}; // @[Cat.scala 30:58]
  wire [47:0] _T_216 = premul_a * premul_b; // @[FMULADD_1G_2.scala 113:19]
  wire  _T_219 = roundRawFNToRecFN_io_out[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_221 = roundRawFNToRecFN_io_out[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  wire  _T_223 = _T_221 & roundRawFNToRecFN_io_out[29]; // @[rawFloatFromRecFN.scala 55:33]
  wire  _T_226 = _T_221 & ~roundRawFNToRecFN_io_out[29]; // @[rawFloatFromRecFN.scala 56:33]
  wire [9:0] _T_228 = {1'b0,$signed(roundRawFNToRecFN_io_out[31:23])}; // @[rawFloatFromRecFN.scala 59:27]
  wire  hi_lo_6 = ~_T_219; // @[rawFloatFromRecFN.scala 60:39]
  wire [22:0] lo_6 = roundRawFNToRecFN_io_out[22:0]; // @[rawFloatFromRecFN.scala 60:51]
  wire [24:0] _T_229 = {1'h0,hi_lo_6,lo_6}; // @[Cat.scala 30:58]
  wire  _T_230 = $signed(_T_228) < 10'sh82; // @[fNFromRecFN.scala 50:39]
  wire [4:0] _T_233 = 5'h1 - _T_228[4:0]; // @[fNFromRecFN.scala 51:39]
  wire [23:0] _T_235 = _T_229[24:1] >> _T_233; // @[fNFromRecFN.scala 52:42]
  wire [7:0] _T_239 = _T_228[7:0] - 8'h81; // @[fNFromRecFN.scala 57:45]
  wire [7:0] _T_240 = _T_230 ? 8'h0 : _T_239; // @[fNFromRecFN.scala 55:16]
  wire  _T_241 = _T_223 | _T_226; // @[fNFromRecFN.scala 59:44]
  wire [7:0] _T_243 = _T_241 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] hi_lo_7 = _T_240 | _T_243; // @[fNFromRecFN.scala 59:15]
  wire [22:0] _T_245 = _T_226 ? 23'h0 : _T_229[22:0]; // @[fNFromRecFN.scala 63:20]
  wire [22:0] lo_7 = _T_230 ? _T_235[22:0] : _T_245; // @[fNFromRecFN.scala 61:16]
  wire [8:0] hi_7 = {roundRawFNToRecFN_io_out[32],hi_lo_7}; // @[Cat.scala 30:58]
  MulAddRecFNToRaw_preMul mulAddRecFNToRaw_preMul ( // @[FMULADD_1G_2.scala 36:15]
    .io_a(mulAddRecFNToRaw_preMul_io_a),
    .io_b(mulAddRecFNToRaw_preMul_io_b),
    .io_c(mulAddRecFNToRaw_preMul_io_c),
    .io_mulAddA(mulAddRecFNToRaw_preMul_io_mulAddA),
    .io_mulAddB(mulAddRecFNToRaw_preMul_io_mulAddB),
    .io_mulAddC(mulAddRecFNToRaw_preMul_io_mulAddC),
    .io_toPostMul_isSigNaNAny(mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny),
    .io_toPostMul_isNaNAOrB(mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB),
    .io_toPostMul_isInfA(mulAddRecFNToRaw_preMul_io_toPostMul_isInfA),
    .io_toPostMul_isZeroA(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA),
    .io_toPostMul_isInfB(mulAddRecFNToRaw_preMul_io_toPostMul_isInfB),
    .io_toPostMul_isZeroB(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB),
    .io_toPostMul_signProd(mulAddRecFNToRaw_preMul_io_toPostMul_signProd),
    .io_toPostMul_isNaNC(mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC),
    .io_toPostMul_isInfC(mulAddRecFNToRaw_preMul_io_toPostMul_isInfC),
    .io_toPostMul_isZeroC(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC),
    .io_toPostMul_sExpSum(mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum),
    .io_toPostMul_doSubMags(mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags),
    .io_toPostMul_CIsDominant(mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant),
    .io_toPostMul_CDom_CAlignDist(mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist),
    .io_toPostMul_highAlignedSigC(mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC),
    .io_toPostMul_bit0AlignedSigC(mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC)
  );
  MulAddRecFNToRaw_postMul mulAddRecFNToRaw_postMul ( // @[FMULADD_1G_2.scala 116:15]
    .io_fromPreMul_isSigNaNAny(mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny),
    .io_fromPreMul_isNaNAOrB(mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB),
    .io_fromPreMul_isInfA(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA),
    .io_fromPreMul_isZeroA(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA),
    .io_fromPreMul_isInfB(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB),
    .io_fromPreMul_isZeroB(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB),
    .io_fromPreMul_signProd(mulAddRecFNToRaw_postMul_io_fromPreMul_signProd),
    .io_fromPreMul_isNaNC(mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC),
    .io_fromPreMul_isInfC(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC),
    .io_fromPreMul_isZeroC(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC),
    .io_fromPreMul_sExpSum(mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum),
    .io_fromPreMul_doSubMags(mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags),
    .io_fromPreMul_CIsDominant(mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant),
    .io_fromPreMul_CDom_CAlignDist(mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist),
    .io_fromPreMul_highAlignedSigC(mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC),
    .io_fromPreMul_bit0AlignedSigC(mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC),
    .io_mulAddResult(mulAddRecFNToRaw_postMul_io_mulAddResult),
    .io_invalidExc(mulAddRecFNToRaw_postMul_io_invalidExc),
    .io_rawOut_isNaN(mulAddRecFNToRaw_postMul_io_rawOut_isNaN),
    .io_rawOut_isInf(mulAddRecFNToRaw_postMul_io_rawOut_isInf),
    .io_rawOut_isZero(mulAddRecFNToRaw_postMul_io_rawOut_isZero),
    .io_rawOut_sign(mulAddRecFNToRaw_postMul_io_rawOut_sign),
    .io_rawOut_sExp(mulAddRecFNToRaw_postMul_io_rawOut_sExp),
    .io_rawOut_sig(mulAddRecFNToRaw_postMul_io_rawOut_sig)
  );
  RoundRawFNToRecFN roundRawFNToRecFN ( // @[FMULADD_1G_2.scala 137:15]
    .io_invalidExc(roundRawFNToRecFN_io_invalidExc),
    .io_in_isNaN(roundRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundRawFNToRecFN_io_in_sig),
    .io_out(roundRawFNToRecFN_io_out)
  );
  assign io_out = {hi_7,lo_7}; // @[Cat.scala 30:58]
  assign mulAddRecFNToRaw_preMul_io_a = {hi_1,lo_1}; // @[Cat.scala 30:58]
  assign mulAddRecFNToRaw_preMul_io_b = {hi_3,lo_3}; // @[Cat.scala 30:58]
  assign mulAddRecFNToRaw_preMul_io_c = {hi_5,lo_5}; // @[Cat.scala 30:58]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny = isSigNaNAny; // @[FMULADD_1G_2.scala 119:84]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB = isNaNAOrB; // @[FMULADD_1G_2.scala 120:86]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA = isInfA; // @[FMULADD_1G_2.scala 121:94]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA = isZeroA; // @[FMULADD_1G_2.scala 122:91]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB = isInfB; // @[FMULADD_1G_2.scala 123:94]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB = isZeroB; // @[FMULADD_1G_2.scala 124:91]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_signProd = signProd; // @[FMULADD_1G_2.scala 125:89]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC = isNaNC; // @[FMULADD_1G_2.scala 126:90]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC = isInfC; // @[FMULADD_1G_2.scala 127:94]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC = isZeroC; // @[FMULADD_1G_2.scala 128:91]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum = sExpSum; // @[FMULADD_1G_2.scala 129:88]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags = doSubMags; // @[FMULADD_1G_2.scala 130:85]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant = CIsDominant; // @[FMULADD_1G_2.scala 131:84]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist = CDom_CAlignDist; // @[FMULADD_1G_2.scala 132:78]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC = highAlignedSigC; // @[FMULADD_1G_2.scala 133:80]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC = bit0AlignedSigC; // @[FMULADD_1G_2.scala 134:82]
  assign mulAddRecFNToRaw_postMul_io_mulAddResult = _T_216 + premul_c; // @[FMULADD_1G_2.scala 113:31]
  assign roundRawFNToRecFN_io_invalidExc = mulAddRecFNToRaw_postMul_io_invalidExc; // @[FMULADD_1G_2.scala 138:39]
  assign roundRawFNToRecFN_io_in_isNaN = mulAddRecFNToRaw_postMul_io_rawOut_isNaN; // @[FMULADD_1G_2.scala 140:39]
  assign roundRawFNToRecFN_io_in_isInf = mulAddRecFNToRaw_postMul_io_rawOut_isInf; // @[FMULADD_1G_2.scala 140:39]
  assign roundRawFNToRecFN_io_in_isZero = mulAddRecFNToRaw_postMul_io_rawOut_isZero; // @[FMULADD_1G_2.scala 140:39]
  assign roundRawFNToRecFN_io_in_sign = mulAddRecFNToRaw_postMul_io_rawOut_sign; // @[FMULADD_1G_2.scala 140:39]
  assign roundRawFNToRecFN_io_in_sExp = mulAddRecFNToRaw_postMul_io_rawOut_sExp; // @[FMULADD_1G_2.scala 140:39]
  assign roundRawFNToRecFN_io_in_sig = mulAddRecFNToRaw_postMul_io_rawOut_sig; // @[FMULADD_1G_2.scala 140:39]
  always @(posedge clock) begin
    if (reset) begin // @[FMULADD_1G_2.scala 15:37]
      premul_a <= 24'h0; // @[FMULADD_1G_2.scala 15:37]
    end else begin
      premul_a <= mulAddRecFNToRaw_preMul_io_mulAddA; // @[FMULADD_1G_2.scala 103:63]
    end
    if (reset) begin // @[FMULADD_1G_2.scala 16:37]
      premul_b <= 24'h0; // @[FMULADD_1G_2.scala 16:37]
    end else begin
      premul_b <= mulAddRecFNToRaw_preMul_io_mulAddB; // @[FMULADD_1G_2.scala 104:63]
    end
    if (reset) begin // @[FMULADD_1G_2.scala 17:37]
      premul_c <= 48'h0; // @[FMULADD_1G_2.scala 17:37]
    end else begin
      premul_c <= mulAddRecFNToRaw_preMul_io_mulAddC; // @[FMULADD_1G_2.scala 105:63]
    end
    if (reset) begin // @[FMULADD_1G_2.scala 18:33]
      isSigNaNAny <= 1'h0; // @[FMULADD_1G_2.scala 18:33]
    end else begin
      isSigNaNAny <= mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny; // @[FMULADD_1G_2.scala 43:61]
    end
    if (reset) begin // @[FMULADD_1G_2.scala 19:34]
      isNaNAOrB <= 1'h0; // @[FMULADD_1G_2.scala 19:34]
    end else begin
      isNaNAOrB <= mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB; // @[FMULADD_1G_2.scala 44:62]
    end
    if (reset) begin // @[FMULADD_1G_2.scala 20:43]
      isInfA <= 1'h0; // @[FMULADD_1G_2.scala 20:43]
    end else begin
      isInfA <= mulAddRecFNToRaw_preMul_io_toPostMul_isInfA; // @[FMULADD_1G_2.scala 45:70]
    end
    if (reset) begin // @[FMULADD_1G_2.scala 21:40]
      isZeroA <= 1'h0; // @[FMULADD_1G_2.scala 21:40]
    end else begin
      isZeroA <= mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA; // @[FMULADD_1G_2.scala 46:67]
    end
    if (reset) begin // @[FMULADD_1G_2.scala 22:43]
      isInfB <= 1'h0; // @[FMULADD_1G_2.scala 22:43]
    end else begin
      isInfB <= mulAddRecFNToRaw_preMul_io_toPostMul_isInfB; // @[FMULADD_1G_2.scala 47:70]
    end
    if (reset) begin // @[FMULADD_1G_2.scala 23:40]
      isZeroB <= 1'h0; // @[FMULADD_1G_2.scala 23:40]
    end else begin
      isZeroB <= mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB; // @[FMULADD_1G_2.scala 48:67]
    end
    if (reset) begin // @[FMULADD_1G_2.scala 24:38]
      signProd <= 1'h0; // @[FMULADD_1G_2.scala 24:38]
    end else begin
      signProd <= mulAddRecFNToRaw_preMul_io_toPostMul_signProd; // @[FMULADD_1G_2.scala 49:65]
    end
    if (reset) begin // @[FMULADD_1G_2.scala 25:39]
      isNaNC <= 1'h0; // @[FMULADD_1G_2.scala 25:39]
    end else begin
      isNaNC <= mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC; // @[FMULADD_1G_2.scala 50:66]
    end
    if (reset) begin // @[FMULADD_1G_2.scala 26:42]
      isInfC <= 1'h0; // @[FMULADD_1G_2.scala 26:42]
    end else begin
      isInfC <= mulAddRecFNToRaw_preMul_io_toPostMul_isInfC; // @[FMULADD_1G_2.scala 51:69]
    end
    if (reset) begin // @[FMULADD_1G_2.scala 27:39]
      isZeroC <= 1'h0; // @[FMULADD_1G_2.scala 27:39]
    end else begin
      isZeroC <= mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC; // @[FMULADD_1G_2.scala 52:66]
    end
    if (reset) begin // @[FMULADD_1G_2.scala 28:36]
      sExpSum <= 10'sh0; // @[FMULADD_1G_2.scala 28:36]
    end else begin
      sExpSum <= mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum; // @[FMULADD_1G_2.scala 53:63]
    end
    if (reset) begin // @[FMULADD_1G_2.scala 29:33]
      doSubMags <= 1'h0; // @[FMULADD_1G_2.scala 29:33]
    end else begin
      doSubMags <= mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags; // @[FMULADD_1G_2.scala 54:60]
    end
    if (reset) begin // @[FMULADD_1G_2.scala 30:33]
      CIsDominant <= 1'h0; // @[FMULADD_1G_2.scala 30:33]
    end else begin
      CIsDominant <= mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant; // @[FMULADD_1G_2.scala 55:59]
    end
    if (reset) begin // @[FMULADD_1G_2.scala 31:34]
      CDom_CAlignDist <= 5'h0; // @[FMULADD_1G_2.scala 31:34]
    end else begin
      CDom_CAlignDist <= mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist; // @[FMULADD_1G_2.scala 56:54]
    end
    if (reset) begin // @[FMULADD_1G_2.scala 32:37]
      highAlignedSigC <= 26'h0; // @[FMULADD_1G_2.scala 32:37]
    end else begin
      highAlignedSigC <= mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC; // @[FMULADD_1G_2.scala 57:56]
    end
    if (reset) begin // @[FMULADD_1G_2.scala 33:38]
      bit0AlignedSigC <= 1'h0; // @[FMULADD_1G_2.scala 33:38]
    end else begin
      bit0AlignedSigC <= mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC; // @[FMULADD_1G_2.scala 58:57]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  premul_a = _RAND_0[23:0];
  _RAND_1 = {1{`RANDOM}};
  premul_b = _RAND_1[23:0];
  _RAND_2 = {2{`RANDOM}};
  premul_c = _RAND_2[47:0];
  _RAND_3 = {1{`RANDOM}};
  isSigNaNAny = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  isNaNAOrB = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  isInfA = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  isZeroA = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  isInfB = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  isZeroB = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  signProd = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  isNaNC = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  isInfC = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  isZeroC = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  sExpSum = _RAND_13[9:0];
  _RAND_14 = {1{`RANDOM}};
  doSubMags = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  CIsDominant = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  CDom_CAlignDist = _RAND_16[4:0];
  _RAND_17 = {1{`RANDOM}};
  highAlignedSigC = _RAND_17[25:0];
  _RAND_18 = {1{`RANDOM}};
  bit0AlignedSigC = _RAND_18[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CompareRecFN(
  input  [32:0] io_a,
  input  [32:0] io_b,
  output        io_lt,
  output        io_eq
);
  wire  rawA_isZero = io_a[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_4 = io_a[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawA_isNaN = _T_4 & io_a[29]; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawA_isInf = _T_4 & ~io_a[29]; // @[rawFloatFromRecFN.scala 56:33]
  wire  rawA_sign = io_a[32]; // @[rawFloatFromRecFN.scala 58:25]
  wire [9:0] rawA_sExp = {1'b0,$signed(io_a[31:23])}; // @[rawFloatFromRecFN.scala 59:27]
  wire  hi_lo = ~rawA_isZero; // @[rawFloatFromRecFN.scala 60:39]
  wire [22:0] lo = io_a[22:0]; // @[rawFloatFromRecFN.scala 60:51]
  wire [24:0] rawA_sig = {1'h0,hi_lo,lo}; // @[Cat.scala 30:58]
  wire  rawB_isZero = io_b[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_17 = io_b[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawB_isNaN = _T_17 & io_b[29]; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawB_isInf = _T_17 & ~io_b[29]; // @[rawFloatFromRecFN.scala 56:33]
  wire  rawB_sign = io_b[32]; // @[rawFloatFromRecFN.scala 58:25]
  wire [9:0] rawB_sExp = {1'b0,$signed(io_b[31:23])}; // @[rawFloatFromRecFN.scala 59:27]
  wire  hi_lo_1 = ~rawB_isZero; // @[rawFloatFromRecFN.scala 60:39]
  wire [22:0] lo_1 = io_b[22:0]; // @[rawFloatFromRecFN.scala 60:51]
  wire [24:0] rawB_sig = {1'h0,hi_lo_1,lo_1}; // @[Cat.scala 30:58]
  wire  ordered = ~rawA_isNaN & ~rawB_isNaN; // @[CompareRecFN.scala 57:32]
  wire  bothInfs = rawA_isInf & rawB_isInf; // @[CompareRecFN.scala 58:33]
  wire  bothZeros = rawA_isZero & rawB_isZero; // @[CompareRecFN.scala 59:33]
  wire  eqExps = $signed(rawA_sExp) == $signed(rawB_sExp); // @[CompareRecFN.scala 60:29]
  wire  common_ltMags = $signed(rawA_sExp) < $signed(rawB_sExp) | eqExps & rawA_sig < rawB_sig; // @[CompareRecFN.scala 62:33]
  wire  common_eqMags = eqExps & rawA_sig == rawB_sig; // @[CompareRecFN.scala 63:32]
  wire  _T_33 = ~rawB_sign; // @[CompareRecFN.scala 67:28]
  wire  _T_41 = _T_33 & common_ltMags; // @[CompareRecFN.scala 70:41]
  wire  _T_42 = rawA_sign & ~common_ltMags & ~common_eqMags | _T_41; // @[CompareRecFN.scala 69:74]
  wire  _T_43 = ~bothInfs & _T_42; // @[CompareRecFN.scala 68:30]
  wire  _T_44 = rawA_sign & ~rawB_sign | _T_43; // @[CompareRecFN.scala 67:41]
  wire  ordered_lt = ~bothZeros & _T_44; // @[CompareRecFN.scala 66:21]
  wire  ordered_eq = bothZeros | rawA_sign == rawB_sign & (bothInfs | common_eqMags); // @[CompareRecFN.scala 72:19]
  assign io_lt = ordered & ordered_lt; // @[CompareRecFN.scala 78:22]
  assign io_eq = ordered & ordered_eq; // @[CompareRecFN.scala 79:22]
endmodule
module ValExec_CompareRecF32_le(
  input  [31:0] io_a,
  input  [31:0] io_b,
  output        io_actual_out
);
  wire [32:0] compareRecFN_io_a; // @[ValExec_CompareRecFN.scala 94:30]
  wire [32:0] compareRecFN_io_b; // @[ValExec_CompareRecFN.scala 94:30]
  wire  compareRecFN_io_lt; // @[ValExec_CompareRecFN.scala 94:30]
  wire  compareRecFN_io_eq; // @[ValExec_CompareRecFN.scala 94:30]
  wire  _T_3 = io_a[30:23] == 8'h0; // @[rawFloatFromFN.scala 50:34]
  wire  _T_4 = io_a[22:0] == 23'h0; // @[rawFloatFromFN.scala 51:38]
  wire [4:0] _T_28 = io_a[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:69]
  wire [4:0] _T_29 = io_a[2] ? 5'h14 : _T_28; // @[Mux.scala 47:69]
  wire [4:0] _T_30 = io_a[3] ? 5'h13 : _T_29; // @[Mux.scala 47:69]
  wire [4:0] _T_31 = io_a[4] ? 5'h12 : _T_30; // @[Mux.scala 47:69]
  wire [4:0] _T_32 = io_a[5] ? 5'h11 : _T_31; // @[Mux.scala 47:69]
  wire [4:0] _T_33 = io_a[6] ? 5'h10 : _T_32; // @[Mux.scala 47:69]
  wire [4:0] _T_34 = io_a[7] ? 5'hf : _T_33; // @[Mux.scala 47:69]
  wire [4:0] _T_35 = io_a[8] ? 5'he : _T_34; // @[Mux.scala 47:69]
  wire [4:0] _T_36 = io_a[9] ? 5'hd : _T_35; // @[Mux.scala 47:69]
  wire [4:0] _T_37 = io_a[10] ? 5'hc : _T_36; // @[Mux.scala 47:69]
  wire [4:0] _T_38 = io_a[11] ? 5'hb : _T_37; // @[Mux.scala 47:69]
  wire [4:0] _T_39 = io_a[12] ? 5'ha : _T_38; // @[Mux.scala 47:69]
  wire [4:0] _T_40 = io_a[13] ? 5'h9 : _T_39; // @[Mux.scala 47:69]
  wire [4:0] _T_41 = io_a[14] ? 5'h8 : _T_40; // @[Mux.scala 47:69]
  wire [4:0] _T_42 = io_a[15] ? 5'h7 : _T_41; // @[Mux.scala 47:69]
  wire [4:0] _T_43 = io_a[16] ? 5'h6 : _T_42; // @[Mux.scala 47:69]
  wire [4:0] _T_44 = io_a[17] ? 5'h5 : _T_43; // @[Mux.scala 47:69]
  wire [4:0] _T_45 = io_a[18] ? 5'h4 : _T_44; // @[Mux.scala 47:69]
  wire [4:0] _T_46 = io_a[19] ? 5'h3 : _T_45; // @[Mux.scala 47:69]
  wire [4:0] _T_47 = io_a[20] ? 5'h2 : _T_46; // @[Mux.scala 47:69]
  wire [4:0] _T_48 = io_a[21] ? 5'h1 : _T_47; // @[Mux.scala 47:69]
  wire [4:0] _T_49 = io_a[22] ? 5'h0 : _T_48; // @[Mux.scala 47:69]
  wire [53:0] _GEN_0 = {{31'd0}, io_a[22:0]}; // @[rawFloatFromFN.scala 54:36]
  wire [53:0] _T_50 = _GEN_0 << _T_49; // @[rawFloatFromFN.scala 54:36]
  wire [22:0] _T_52 = {_T_50[21:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  wire [8:0] _GEN_1 = {{4'd0}, _T_49}; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_53 = _GEN_1 ^ 9'h1ff; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_54 = _T_3 ? _T_53 : {{1'd0}, io_a[30:23]}; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_55 = _T_3 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  wire [7:0] _GEN_2 = {{6'd0}, _T_55}; // @[rawFloatFromFN.scala 60:22]
  wire [7:0] _T_56 = 8'h80 | _GEN_2; // @[rawFloatFromFN.scala 60:22]
  wire [8:0] _GEN_3 = {{1'd0}, _T_56}; // @[rawFloatFromFN.scala 59:15]
  wire [8:0] _T_58 = _T_54 + _GEN_3; // @[rawFloatFromFN.scala 59:15]
  wire  _T_59 = _T_3 & _T_4; // @[rawFloatFromFN.scala 62:34]
  wire  _T_61 = _T_58[8:7] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  wire  _T_63 = _T_61 & ~_T_4; // @[rawFloatFromFN.scala 66:33]
  wire [9:0] _T_66 = {1'b0,$signed(_T_58)}; // @[rawFloatFromFN.scala 70:48]
  wire  hi_lo = ~_T_59; // @[rawFloatFromFN.scala 72:29]
  wire [22:0] lo = _T_3 ? _T_52 : io_a[22:0]; // @[rawFloatFromFN.scala 72:42]
  wire [24:0] _T_67 = {1'h0,hi_lo,lo}; // @[Cat.scala 30:58]
  wire [2:0] _T_69 = _T_59 ? 3'h0 : _T_66[8:6]; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_4 = {{2'd0}, _T_63}; // @[recFNFromFN.scala 48:79]
  wire [2:0] hi_lo_1 = _T_69 | _GEN_4; // @[recFNFromFN.scala 48:79]
  wire [5:0] lo_hi = _T_66[5:0]; // @[recFNFromFN.scala 50:23]
  wire [22:0] lo_lo = _T_67[22:0]; // @[recFNFromFN.scala 51:22]
  wire [28:0] lo_1 = {lo_hi,lo_lo}; // @[Cat.scala 30:58]
  wire [3:0] hi_1 = {io_a[31],hi_lo_1}; // @[Cat.scala 30:58]
  wire  _T_75 = io_b[30:23] == 8'h0; // @[rawFloatFromFN.scala 50:34]
  wire  _T_76 = io_b[22:0] == 23'h0; // @[rawFloatFromFN.scala 51:38]
  wire [4:0] _T_100 = io_b[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:69]
  wire [4:0] _T_101 = io_b[2] ? 5'h14 : _T_100; // @[Mux.scala 47:69]
  wire [4:0] _T_102 = io_b[3] ? 5'h13 : _T_101; // @[Mux.scala 47:69]
  wire [4:0] _T_103 = io_b[4] ? 5'h12 : _T_102; // @[Mux.scala 47:69]
  wire [4:0] _T_104 = io_b[5] ? 5'h11 : _T_103; // @[Mux.scala 47:69]
  wire [4:0] _T_105 = io_b[6] ? 5'h10 : _T_104; // @[Mux.scala 47:69]
  wire [4:0] _T_106 = io_b[7] ? 5'hf : _T_105; // @[Mux.scala 47:69]
  wire [4:0] _T_107 = io_b[8] ? 5'he : _T_106; // @[Mux.scala 47:69]
  wire [4:0] _T_108 = io_b[9] ? 5'hd : _T_107; // @[Mux.scala 47:69]
  wire [4:0] _T_109 = io_b[10] ? 5'hc : _T_108; // @[Mux.scala 47:69]
  wire [4:0] _T_110 = io_b[11] ? 5'hb : _T_109; // @[Mux.scala 47:69]
  wire [4:0] _T_111 = io_b[12] ? 5'ha : _T_110; // @[Mux.scala 47:69]
  wire [4:0] _T_112 = io_b[13] ? 5'h9 : _T_111; // @[Mux.scala 47:69]
  wire [4:0] _T_113 = io_b[14] ? 5'h8 : _T_112; // @[Mux.scala 47:69]
  wire [4:0] _T_114 = io_b[15] ? 5'h7 : _T_113; // @[Mux.scala 47:69]
  wire [4:0] _T_115 = io_b[16] ? 5'h6 : _T_114; // @[Mux.scala 47:69]
  wire [4:0] _T_116 = io_b[17] ? 5'h5 : _T_115; // @[Mux.scala 47:69]
  wire [4:0] _T_117 = io_b[18] ? 5'h4 : _T_116; // @[Mux.scala 47:69]
  wire [4:0] _T_118 = io_b[19] ? 5'h3 : _T_117; // @[Mux.scala 47:69]
  wire [4:0] _T_119 = io_b[20] ? 5'h2 : _T_118; // @[Mux.scala 47:69]
  wire [4:0] _T_120 = io_b[21] ? 5'h1 : _T_119; // @[Mux.scala 47:69]
  wire [4:0] _T_121 = io_b[22] ? 5'h0 : _T_120; // @[Mux.scala 47:69]
  wire [53:0] _GEN_5 = {{31'd0}, io_b[22:0]}; // @[rawFloatFromFN.scala 54:36]
  wire [53:0] _T_122 = _GEN_5 << _T_121; // @[rawFloatFromFN.scala 54:36]
  wire [22:0] _T_124 = {_T_122[21:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  wire [8:0] _GEN_6 = {{4'd0}, _T_121}; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_125 = _GEN_6 ^ 9'h1ff; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_126 = _T_75 ? _T_125 : {{1'd0}, io_b[30:23]}; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_127 = _T_75 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  wire [7:0] _GEN_7 = {{6'd0}, _T_127}; // @[rawFloatFromFN.scala 60:22]
  wire [7:0] _T_128 = 8'h80 | _GEN_7; // @[rawFloatFromFN.scala 60:22]
  wire [8:0] _GEN_8 = {{1'd0}, _T_128}; // @[rawFloatFromFN.scala 59:15]
  wire [8:0] _T_130 = _T_126 + _GEN_8; // @[rawFloatFromFN.scala 59:15]
  wire  _T_131 = _T_75 & _T_76; // @[rawFloatFromFN.scala 62:34]
  wire  _T_133 = _T_130[8:7] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  wire  _T_135 = _T_133 & ~_T_76; // @[rawFloatFromFN.scala 66:33]
  wire [9:0] _T_138 = {1'b0,$signed(_T_130)}; // @[rawFloatFromFN.scala 70:48]
  wire  hi_lo_2 = ~_T_131; // @[rawFloatFromFN.scala 72:29]
  wire [22:0] lo_2 = _T_75 ? _T_124 : io_b[22:0]; // @[rawFloatFromFN.scala 72:42]
  wire [24:0] _T_139 = {1'h0,hi_lo_2,lo_2}; // @[Cat.scala 30:58]
  wire [2:0] _T_141 = _T_131 ? 3'h0 : _T_138[8:6]; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_9 = {{2'd0}, _T_135}; // @[recFNFromFN.scala 48:79]
  wire [2:0] hi_lo_3 = _T_141 | _GEN_9; // @[recFNFromFN.scala 48:79]
  wire [5:0] lo_hi_1 = _T_138[5:0]; // @[recFNFromFN.scala 50:23]
  wire [22:0] lo_lo_1 = _T_139[22:0]; // @[recFNFromFN.scala 51:22]
  wire [28:0] lo_3 = {lo_hi_1,lo_lo_1}; // @[Cat.scala 30:58]
  wire [3:0] hi_3 = {io_b[31],hi_lo_3}; // @[Cat.scala 30:58]
  CompareRecFN compareRecFN ( // @[ValExec_CompareRecFN.scala 94:30]
    .io_a(compareRecFN_io_a),
    .io_b(compareRecFN_io_b),
    .io_lt(compareRecFN_io_lt),
    .io_eq(compareRecFN_io_eq)
  );
  assign io_actual_out = compareRecFN_io_lt | compareRecFN_io_eq; // @[ValExec_CompareRecFN.scala 99:41]
  assign compareRecFN_io_a = {hi_1,lo_1}; // @[Cat.scala 30:58]
  assign compareRecFN_io_b = {hi_3,lo_3}; // @[Cat.scala 30:58]
endmodule
module ValExec_CompareRecF32_lt(
  input  [31:0] io_a,
  input  [31:0] io_b,
  output        io_actual_out
);
  wire [32:0] compareRecFN_io_a; // @[ValExec_CompareRecFN.scala 59:30]
  wire [32:0] compareRecFN_io_b; // @[ValExec_CompareRecFN.scala 59:30]
  wire  compareRecFN_io_lt; // @[ValExec_CompareRecFN.scala 59:30]
  wire  compareRecFN_io_eq; // @[ValExec_CompareRecFN.scala 59:30]
  wire  _T_3 = io_a[30:23] == 8'h0; // @[rawFloatFromFN.scala 50:34]
  wire  _T_4 = io_a[22:0] == 23'h0; // @[rawFloatFromFN.scala 51:38]
  wire [4:0] _T_28 = io_a[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:69]
  wire [4:0] _T_29 = io_a[2] ? 5'h14 : _T_28; // @[Mux.scala 47:69]
  wire [4:0] _T_30 = io_a[3] ? 5'h13 : _T_29; // @[Mux.scala 47:69]
  wire [4:0] _T_31 = io_a[4] ? 5'h12 : _T_30; // @[Mux.scala 47:69]
  wire [4:0] _T_32 = io_a[5] ? 5'h11 : _T_31; // @[Mux.scala 47:69]
  wire [4:0] _T_33 = io_a[6] ? 5'h10 : _T_32; // @[Mux.scala 47:69]
  wire [4:0] _T_34 = io_a[7] ? 5'hf : _T_33; // @[Mux.scala 47:69]
  wire [4:0] _T_35 = io_a[8] ? 5'he : _T_34; // @[Mux.scala 47:69]
  wire [4:0] _T_36 = io_a[9] ? 5'hd : _T_35; // @[Mux.scala 47:69]
  wire [4:0] _T_37 = io_a[10] ? 5'hc : _T_36; // @[Mux.scala 47:69]
  wire [4:0] _T_38 = io_a[11] ? 5'hb : _T_37; // @[Mux.scala 47:69]
  wire [4:0] _T_39 = io_a[12] ? 5'ha : _T_38; // @[Mux.scala 47:69]
  wire [4:0] _T_40 = io_a[13] ? 5'h9 : _T_39; // @[Mux.scala 47:69]
  wire [4:0] _T_41 = io_a[14] ? 5'h8 : _T_40; // @[Mux.scala 47:69]
  wire [4:0] _T_42 = io_a[15] ? 5'h7 : _T_41; // @[Mux.scala 47:69]
  wire [4:0] _T_43 = io_a[16] ? 5'h6 : _T_42; // @[Mux.scala 47:69]
  wire [4:0] _T_44 = io_a[17] ? 5'h5 : _T_43; // @[Mux.scala 47:69]
  wire [4:0] _T_45 = io_a[18] ? 5'h4 : _T_44; // @[Mux.scala 47:69]
  wire [4:0] _T_46 = io_a[19] ? 5'h3 : _T_45; // @[Mux.scala 47:69]
  wire [4:0] _T_47 = io_a[20] ? 5'h2 : _T_46; // @[Mux.scala 47:69]
  wire [4:0] _T_48 = io_a[21] ? 5'h1 : _T_47; // @[Mux.scala 47:69]
  wire [4:0] _T_49 = io_a[22] ? 5'h0 : _T_48; // @[Mux.scala 47:69]
  wire [53:0] _GEN_0 = {{31'd0}, io_a[22:0]}; // @[rawFloatFromFN.scala 54:36]
  wire [53:0] _T_50 = _GEN_0 << _T_49; // @[rawFloatFromFN.scala 54:36]
  wire [22:0] _T_52 = {_T_50[21:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  wire [8:0] _GEN_1 = {{4'd0}, _T_49}; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_53 = _GEN_1 ^ 9'h1ff; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_54 = _T_3 ? _T_53 : {{1'd0}, io_a[30:23]}; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_55 = _T_3 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  wire [7:0] _GEN_2 = {{6'd0}, _T_55}; // @[rawFloatFromFN.scala 60:22]
  wire [7:0] _T_56 = 8'h80 | _GEN_2; // @[rawFloatFromFN.scala 60:22]
  wire [8:0] _GEN_3 = {{1'd0}, _T_56}; // @[rawFloatFromFN.scala 59:15]
  wire [8:0] _T_58 = _T_54 + _GEN_3; // @[rawFloatFromFN.scala 59:15]
  wire  _T_59 = _T_3 & _T_4; // @[rawFloatFromFN.scala 62:34]
  wire  _T_61 = _T_58[8:7] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  wire  _T_63 = _T_61 & ~_T_4; // @[rawFloatFromFN.scala 66:33]
  wire [9:0] _T_66 = {1'b0,$signed(_T_58)}; // @[rawFloatFromFN.scala 70:48]
  wire  hi_lo = ~_T_59; // @[rawFloatFromFN.scala 72:29]
  wire [22:0] lo = _T_3 ? _T_52 : io_a[22:0]; // @[rawFloatFromFN.scala 72:42]
  wire [24:0] _T_67 = {1'h0,hi_lo,lo}; // @[Cat.scala 30:58]
  wire [2:0] _T_69 = _T_59 ? 3'h0 : _T_66[8:6]; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_4 = {{2'd0}, _T_63}; // @[recFNFromFN.scala 48:79]
  wire [2:0] hi_lo_1 = _T_69 | _GEN_4; // @[recFNFromFN.scala 48:79]
  wire [5:0] lo_hi = _T_66[5:0]; // @[recFNFromFN.scala 50:23]
  wire [22:0] lo_lo = _T_67[22:0]; // @[recFNFromFN.scala 51:22]
  wire [28:0] lo_1 = {lo_hi,lo_lo}; // @[Cat.scala 30:58]
  wire [3:0] hi_1 = {io_a[31],hi_lo_1}; // @[Cat.scala 30:58]
  wire  _T_75 = io_b[30:23] == 8'h0; // @[rawFloatFromFN.scala 50:34]
  wire  _T_76 = io_b[22:0] == 23'h0; // @[rawFloatFromFN.scala 51:38]
  wire [4:0] _T_100 = io_b[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:69]
  wire [4:0] _T_101 = io_b[2] ? 5'h14 : _T_100; // @[Mux.scala 47:69]
  wire [4:0] _T_102 = io_b[3] ? 5'h13 : _T_101; // @[Mux.scala 47:69]
  wire [4:0] _T_103 = io_b[4] ? 5'h12 : _T_102; // @[Mux.scala 47:69]
  wire [4:0] _T_104 = io_b[5] ? 5'h11 : _T_103; // @[Mux.scala 47:69]
  wire [4:0] _T_105 = io_b[6] ? 5'h10 : _T_104; // @[Mux.scala 47:69]
  wire [4:0] _T_106 = io_b[7] ? 5'hf : _T_105; // @[Mux.scala 47:69]
  wire [4:0] _T_107 = io_b[8] ? 5'he : _T_106; // @[Mux.scala 47:69]
  wire [4:0] _T_108 = io_b[9] ? 5'hd : _T_107; // @[Mux.scala 47:69]
  wire [4:0] _T_109 = io_b[10] ? 5'hc : _T_108; // @[Mux.scala 47:69]
  wire [4:0] _T_110 = io_b[11] ? 5'hb : _T_109; // @[Mux.scala 47:69]
  wire [4:0] _T_111 = io_b[12] ? 5'ha : _T_110; // @[Mux.scala 47:69]
  wire [4:0] _T_112 = io_b[13] ? 5'h9 : _T_111; // @[Mux.scala 47:69]
  wire [4:0] _T_113 = io_b[14] ? 5'h8 : _T_112; // @[Mux.scala 47:69]
  wire [4:0] _T_114 = io_b[15] ? 5'h7 : _T_113; // @[Mux.scala 47:69]
  wire [4:0] _T_115 = io_b[16] ? 5'h6 : _T_114; // @[Mux.scala 47:69]
  wire [4:0] _T_116 = io_b[17] ? 5'h5 : _T_115; // @[Mux.scala 47:69]
  wire [4:0] _T_117 = io_b[18] ? 5'h4 : _T_116; // @[Mux.scala 47:69]
  wire [4:0] _T_118 = io_b[19] ? 5'h3 : _T_117; // @[Mux.scala 47:69]
  wire [4:0] _T_119 = io_b[20] ? 5'h2 : _T_118; // @[Mux.scala 47:69]
  wire [4:0] _T_120 = io_b[21] ? 5'h1 : _T_119; // @[Mux.scala 47:69]
  wire [4:0] _T_121 = io_b[22] ? 5'h0 : _T_120; // @[Mux.scala 47:69]
  wire [53:0] _GEN_5 = {{31'd0}, io_b[22:0]}; // @[rawFloatFromFN.scala 54:36]
  wire [53:0] _T_122 = _GEN_5 << _T_121; // @[rawFloatFromFN.scala 54:36]
  wire [22:0] _T_124 = {_T_122[21:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  wire [8:0] _GEN_6 = {{4'd0}, _T_121}; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_125 = _GEN_6 ^ 9'h1ff; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_126 = _T_75 ? _T_125 : {{1'd0}, io_b[30:23]}; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_127 = _T_75 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  wire [7:0] _GEN_7 = {{6'd0}, _T_127}; // @[rawFloatFromFN.scala 60:22]
  wire [7:0] _T_128 = 8'h80 | _GEN_7; // @[rawFloatFromFN.scala 60:22]
  wire [8:0] _GEN_8 = {{1'd0}, _T_128}; // @[rawFloatFromFN.scala 59:15]
  wire [8:0] _T_130 = _T_126 + _GEN_8; // @[rawFloatFromFN.scala 59:15]
  wire  _T_131 = _T_75 & _T_76; // @[rawFloatFromFN.scala 62:34]
  wire  _T_133 = _T_130[8:7] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  wire  _T_135 = _T_133 & ~_T_76; // @[rawFloatFromFN.scala 66:33]
  wire [9:0] _T_138 = {1'b0,$signed(_T_130)}; // @[rawFloatFromFN.scala 70:48]
  wire  hi_lo_2 = ~_T_131; // @[rawFloatFromFN.scala 72:29]
  wire [22:0] lo_2 = _T_75 ? _T_124 : io_b[22:0]; // @[rawFloatFromFN.scala 72:42]
  wire [24:0] _T_139 = {1'h0,hi_lo_2,lo_2}; // @[Cat.scala 30:58]
  wire [2:0] _T_141 = _T_131 ? 3'h0 : _T_138[8:6]; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_9 = {{2'd0}, _T_135}; // @[recFNFromFN.scala 48:79]
  wire [2:0] hi_lo_3 = _T_141 | _GEN_9; // @[recFNFromFN.scala 48:79]
  wire [5:0] lo_hi_1 = _T_138[5:0]; // @[recFNFromFN.scala 50:23]
  wire [22:0] lo_lo_1 = _T_139[22:0]; // @[recFNFromFN.scala 51:22]
  wire [28:0] lo_3 = {lo_hi_1,lo_lo_1}; // @[Cat.scala 30:58]
  wire [3:0] hi_3 = {io_b[31],hi_lo_3}; // @[Cat.scala 30:58]
  CompareRecFN compareRecFN ( // @[ValExec_CompareRecFN.scala 59:30]
    .io_a(compareRecFN_io_a),
    .io_b(compareRecFN_io_b),
    .io_lt(compareRecFN_io_lt),
    .io_eq(compareRecFN_io_eq)
  );
  assign io_actual_out = compareRecFN_io_lt; // @[ValExec_CompareRecFN.scala 64:19]
  assign compareRecFN_io_a = {hi_1,lo_1}; // @[Cat.scala 30:58]
  assign compareRecFN_io_b = {hi_3,lo_3}; // @[Cat.scala 30:58]
endmodule
module ray_AABB_1(
  input         clock,
  input         reset,
  input  [31:0] io_ray_idir_x,
  input  [31:0] io_ray_idir_y,
  input  [31:0] io_ray_idir_z,
  input  [31:0] io_ray_ood_x,
  input  [31:0] io_ray_ood_y,
  input  [31:0] io_ray_ood_z,
  input  [31:0] io_ray_hitT,
  input  [31:0] io_bvh_n0xy_x,
  input  [31:0] io_bvh_n0xy_y,
  input  [31:0] io_bvh_n0xy_z,
  input  [31:0] io_bvh_n0xy_w,
  input  [31:0] io_bvh_n1xy_x,
  input  [31:0] io_bvh_n1xy_y,
  input  [31:0] io_bvh_n1xy_z,
  input  [31:0] io_bvh_n1xy_w,
  input  [31:0] io_bvh_nz_x,
  input  [31:0] io_bvh_nz_y,
  input  [31:0] io_bvh_nz_z,
  input  [31:0] io_bvh_nz_w,
  input  [31:0] io_bvh_temp_x,
  input  [31:0] io_bvh_temp_y,
  input  [31:0] io_rayid,
  input         io_valid_en,
  output [31:0] io_rayid_out,
  output [31:0] io_nodeIdx_0,
  output [31:0] io_nodeIdx_1,
  output [31:0] io_nodeIdx_2,
  output        io_push,
  output        io_pop,
  output        io_leaf,
  output        io_back,
  output [31:0] io_hitT_out,
  output        io_valid_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
`endif // RANDOMIZE_REG_INIT
  wire  FADD_MUL_1_clock; // @[Ray_AABB_1.scala 80:33]
  wire  FADD_MUL_1_reset; // @[Ray_AABB_1.scala 80:33]
  wire [31:0] FADD_MUL_1_io_a; // @[Ray_AABB_1.scala 80:33]
  wire [31:0] FADD_MUL_1_io_b; // @[Ray_AABB_1.scala 80:33]
  wire [31:0] FADD_MUL_1_io_c; // @[Ray_AABB_1.scala 80:33]
  wire [31:0] FADD_MUL_1_io_out; // @[Ray_AABB_1.scala 80:33]
  wire  FADD_MUL_2_clock; // @[Ray_AABB_1.scala 90:33]
  wire  FADD_MUL_2_reset; // @[Ray_AABB_1.scala 90:33]
  wire [31:0] FADD_MUL_2_io_a; // @[Ray_AABB_1.scala 90:33]
  wire [31:0] FADD_MUL_2_io_b; // @[Ray_AABB_1.scala 90:33]
  wire [31:0] FADD_MUL_2_io_c; // @[Ray_AABB_1.scala 90:33]
  wire [31:0] FADD_MUL_2_io_out; // @[Ray_AABB_1.scala 90:33]
  wire  FADD_MUL_3_clock; // @[Ray_AABB_1.scala 100:33]
  wire  FADD_MUL_3_reset; // @[Ray_AABB_1.scala 100:33]
  wire [31:0] FADD_MUL_3_io_a; // @[Ray_AABB_1.scala 100:33]
  wire [31:0] FADD_MUL_3_io_b; // @[Ray_AABB_1.scala 100:33]
  wire [31:0] FADD_MUL_3_io_c; // @[Ray_AABB_1.scala 100:33]
  wire [31:0] FADD_MUL_3_io_out; // @[Ray_AABB_1.scala 100:33]
  wire  FADD_MUL_4_clock; // @[Ray_AABB_1.scala 110:33]
  wire  FADD_MUL_4_reset; // @[Ray_AABB_1.scala 110:33]
  wire [31:0] FADD_MUL_4_io_a; // @[Ray_AABB_1.scala 110:33]
  wire [31:0] FADD_MUL_4_io_b; // @[Ray_AABB_1.scala 110:33]
  wire [31:0] FADD_MUL_4_io_c; // @[Ray_AABB_1.scala 110:33]
  wire [31:0] FADD_MUL_4_io_out; // @[Ray_AABB_1.scala 110:33]
  wire  FADD_MUL_5_clock; // @[Ray_AABB_1.scala 120:33]
  wire  FADD_MUL_5_reset; // @[Ray_AABB_1.scala 120:33]
  wire [31:0] FADD_MUL_5_io_a; // @[Ray_AABB_1.scala 120:33]
  wire [31:0] FADD_MUL_5_io_b; // @[Ray_AABB_1.scala 120:33]
  wire [31:0] FADD_MUL_5_io_c; // @[Ray_AABB_1.scala 120:33]
  wire [31:0] FADD_MUL_5_io_out; // @[Ray_AABB_1.scala 120:33]
  wire  FADD_MUL_6_clock; // @[Ray_AABB_1.scala 130:33]
  wire  FADD_MUL_6_reset; // @[Ray_AABB_1.scala 130:33]
  wire [31:0] FADD_MUL_6_io_a; // @[Ray_AABB_1.scala 130:33]
  wire [31:0] FADD_MUL_6_io_b; // @[Ray_AABB_1.scala 130:33]
  wire [31:0] FADD_MUL_6_io_c; // @[Ray_AABB_1.scala 130:33]
  wire [31:0] FADD_MUL_6_io_out; // @[Ray_AABB_1.scala 130:33]
  wire  FADD_MUL_7_clock; // @[Ray_AABB_1.scala 140:33]
  wire  FADD_MUL_7_reset; // @[Ray_AABB_1.scala 140:33]
  wire [31:0] FADD_MUL_7_io_a; // @[Ray_AABB_1.scala 140:33]
  wire [31:0] FADD_MUL_7_io_b; // @[Ray_AABB_1.scala 140:33]
  wire [31:0] FADD_MUL_7_io_c; // @[Ray_AABB_1.scala 140:33]
  wire [31:0] FADD_MUL_7_io_out; // @[Ray_AABB_1.scala 140:33]
  wire  FADD_MUL_8_clock; // @[Ray_AABB_1.scala 150:33]
  wire  FADD_MUL_8_reset; // @[Ray_AABB_1.scala 150:33]
  wire [31:0] FADD_MUL_8_io_a; // @[Ray_AABB_1.scala 150:33]
  wire [31:0] FADD_MUL_8_io_b; // @[Ray_AABB_1.scala 150:33]
  wire [31:0] FADD_MUL_8_io_c; // @[Ray_AABB_1.scala 150:33]
  wire [31:0] FADD_MUL_8_io_out; // @[Ray_AABB_1.scala 150:33]
  wire  FADD_MUL_9_clock; // @[Ray_AABB_1.scala 160:33]
  wire  FADD_MUL_9_reset; // @[Ray_AABB_1.scala 160:33]
  wire [31:0] FADD_MUL_9_io_a; // @[Ray_AABB_1.scala 160:33]
  wire [31:0] FADD_MUL_9_io_b; // @[Ray_AABB_1.scala 160:33]
  wire [31:0] FADD_MUL_9_io_c; // @[Ray_AABB_1.scala 160:33]
  wire [31:0] FADD_MUL_9_io_out; // @[Ray_AABB_1.scala 160:33]
  wire  FADD_MUL_10_clock; // @[Ray_AABB_1.scala 170:33]
  wire  FADD_MUL_10_reset; // @[Ray_AABB_1.scala 170:33]
  wire [31:0] FADD_MUL_10_io_a; // @[Ray_AABB_1.scala 170:33]
  wire [31:0] FADD_MUL_10_io_b; // @[Ray_AABB_1.scala 170:33]
  wire [31:0] FADD_MUL_10_io_c; // @[Ray_AABB_1.scala 170:33]
  wire [31:0] FADD_MUL_10_io_out; // @[Ray_AABB_1.scala 170:33]
  wire  FADD_MUL_11_clock; // @[Ray_AABB_1.scala 180:33]
  wire  FADD_MUL_11_reset; // @[Ray_AABB_1.scala 180:33]
  wire [31:0] FADD_MUL_11_io_a; // @[Ray_AABB_1.scala 180:33]
  wire [31:0] FADD_MUL_11_io_b; // @[Ray_AABB_1.scala 180:33]
  wire [31:0] FADD_MUL_11_io_c; // @[Ray_AABB_1.scala 180:33]
  wire [31:0] FADD_MUL_11_io_out; // @[Ray_AABB_1.scala 180:33]
  wire  FADD_MUL_12_clock; // @[Ray_AABB_1.scala 190:33]
  wire  FADD_MUL_12_reset; // @[Ray_AABB_1.scala 190:33]
  wire [31:0] FADD_MUL_12_io_a; // @[Ray_AABB_1.scala 190:33]
  wire [31:0] FADD_MUL_12_io_b; // @[Ray_AABB_1.scala 190:33]
  wire [31:0] FADD_MUL_12_io_c; // @[Ray_AABB_1.scala 190:33]
  wire [31:0] FADD_MUL_12_io_out; // @[Ray_AABB_1.scala 190:33]
  wire [31:0] FCMP_1_io_a; // @[Ray_AABB_1.scala 238:24]
  wire [31:0] FCMP_1_io_b; // @[Ray_AABB_1.scala 238:24]
  wire  FCMP_1_io_actual_out; // @[Ray_AABB_1.scala 238:24]
  wire [31:0] FCMP_2_io_a; // @[Ray_AABB_1.scala 253:24]
  wire [31:0] FCMP_2_io_b; // @[Ray_AABB_1.scala 253:24]
  wire  FCMP_2_io_actual_out; // @[Ray_AABB_1.scala 253:24]
  wire [31:0] FCMP_3_io_a; // @[Ray_AABB_1.scala 266:24]
  wire [31:0] FCMP_3_io_b; // @[Ray_AABB_1.scala 266:24]
  wire  FCMP_3_io_actual_out; // @[Ray_AABB_1.scala 266:24]
  wire [31:0] FCMP_4_io_a; // @[Ray_AABB_1.scala 279:24]
  wire [31:0] FCMP_4_io_b; // @[Ray_AABB_1.scala 279:24]
  wire  FCMP_4_io_actual_out; // @[Ray_AABB_1.scala 279:24]
  wire [31:0] FCMP_5_io_a; // @[Ray_AABB_1.scala 292:25]
  wire [31:0] FCMP_5_io_b; // @[Ray_AABB_1.scala 292:25]
  wire  FCMP_5_io_actual_out; // @[Ray_AABB_1.scala 292:25]
  wire [31:0] FCMP_6_io_a; // @[Ray_AABB_1.scala 305:24]
  wire [31:0] FCMP_6_io_b; // @[Ray_AABB_1.scala 305:24]
  wire  FCMP_6_io_actual_out; // @[Ray_AABB_1.scala 305:24]
  wire [31:0] FCMP_7_io_a; // @[Ray_AABB_1.scala 350:24]
  wire [31:0] FCMP_7_io_b; // @[Ray_AABB_1.scala 350:24]
  wire  FCMP_7_io_actual_out; // @[Ray_AABB_1.scala 350:24]
  wire [31:0] FCMP_8_io_a; // @[Ray_AABB_1.scala 361:24]
  wire [31:0] FCMP_8_io_b; // @[Ray_AABB_1.scala 361:24]
  wire  FCMP_8_io_actual_out; // @[Ray_AABB_1.scala 361:24]
  wire [31:0] FCMP_9_io_a; // @[Ray_AABB_1.scala 372:24]
  wire [31:0] FCMP_9_io_b; // @[Ray_AABB_1.scala 372:24]
  wire  FCMP_9_io_actual_out; // @[Ray_AABB_1.scala 372:24]
  wire [31:0] FCMP_10_io_a; // @[Ray_AABB_1.scala 383:25]
  wire [31:0] FCMP_10_io_b; // @[Ray_AABB_1.scala 383:25]
  wire  FCMP_10_io_actual_out; // @[Ray_AABB_1.scala 383:25]
  wire [31:0] FCMP_11_io_a; // @[Ray_AABB_1.scala 394:25]
  wire [31:0] FCMP_11_io_b; // @[Ray_AABB_1.scala 394:25]
  wire  FCMP_11_io_actual_out; // @[Ray_AABB_1.scala 394:25]
  wire [31:0] FCMP_12_io_a; // @[Ray_AABB_1.scala 405:25]
  wire [31:0] FCMP_12_io_b; // @[Ray_AABB_1.scala 405:25]
  wire  FCMP_12_io_actual_out; // @[Ray_AABB_1.scala 405:25]
  wire [31:0] FCMP_13_io_a; // @[Ray_AABB_1.scala 416:25]
  wire [31:0] FCMP_13_io_b; // @[Ray_AABB_1.scala 416:25]
  wire  FCMP_13_io_actual_out; // @[Ray_AABB_1.scala 416:25]
  wire [31:0] FCMP_14_io_a; // @[Ray_AABB_1.scala 427:25]
  wire [31:0] FCMP_14_io_b; // @[Ray_AABB_1.scala 427:25]
  wire  FCMP_14_io_actual_out; // @[Ray_AABB_1.scala 427:25]
  wire [31:0] FCMP_15_io_a; // @[Ray_AABB_1.scala 465:25]
  wire [31:0] FCMP_15_io_b; // @[Ray_AABB_1.scala 465:25]
  wire  FCMP_15_io_actual_out; // @[Ray_AABB_1.scala 465:25]
  wire [31:0] FCMP_16_io_a; // @[Ray_AABB_1.scala 476:25]
  wire [31:0] FCMP_16_io_b; // @[Ray_AABB_1.scala 476:25]
  wire  FCMP_16_io_actual_out; // @[Ray_AABB_1.scala 476:25]
  wire [31:0] FCMP_17_io_a; // @[Ray_AABB_1.scala 487:25]
  wire [31:0] FCMP_17_io_b; // @[Ray_AABB_1.scala 487:25]
  wire  FCMP_17_io_actual_out; // @[Ray_AABB_1.scala 487:25]
  wire [31:0] FCMP_18_io_a; // @[Ray_AABB_1.scala 498:25]
  wire [31:0] FCMP_18_io_b; // @[Ray_AABB_1.scala 498:25]
  wire  FCMP_18_io_actual_out; // @[Ray_AABB_1.scala 498:25]
  wire [31:0] FCMP_19_io_a; // @[Ray_AABB_1.scala 541:25]
  wire [31:0] FCMP_19_io_b; // @[Ray_AABB_1.scala 541:25]
  wire  FCMP_19_io_actual_out; // @[Ray_AABB_1.scala 541:25]
  wire [31:0] FCMP_20_io_a; // @[Ray_AABB_1.scala 554:25]
  wire [31:0] FCMP_20_io_b; // @[Ray_AABB_1.scala 554:25]
  wire  FCMP_20_io_actual_out; // @[Ray_AABB_1.scala 554:25]
  wire [31:0] FCMP_21_io_a; // @[Ray_AABB_1.scala 567:25]
  wire [31:0] FCMP_21_io_b; // @[Ray_AABB_1.scala 567:25]
  wire  FCMP_21_io_actual_out; // @[Ray_AABB_1.scala 567:25]
  reg  traverseChild0; // @[Ray_AABB_1.scala 32:33]
  reg  traverseChild1; // @[Ray_AABB_1.scala 33:33]
  reg [31:0] c0lox; // @[Ray_AABB_1.scala 35:34]
  reg [31:0] c0hix; // @[Ray_AABB_1.scala 36:34]
  reg [31:0] c0loy; // @[Ray_AABB_1.scala 37:34]
  reg [31:0] c0hiy; // @[Ray_AABB_1.scala 38:33]
  reg [31:0] c0loz; // @[Ray_AABB_1.scala 39:34]
  reg [31:0] c0hiz; // @[Ray_AABB_1.scala 40:34]
  reg [31:0] c1lox; // @[Ray_AABB_1.scala 42:34]
  reg [31:0] c1hix; // @[Ray_AABB_1.scala 43:34]
  reg [31:0] c1loy; // @[Ray_AABB_1.scala 44:34]
  reg [31:0] c1hiy; // @[Ray_AABB_1.scala 45:34]
  reg [31:0] c1loz; // @[Ray_AABB_1.scala 46:34]
  reg [31:0] c1hiz; // @[Ray_AABB_1.scala 47:34]
  reg [31:0] rayid_1; // @[Ray_AABB_1.scala 49:32]
  reg [31:0] hitT_1; // @[Ray_AABB_1.scala 50:33]
  reg [31:0] valid_1; // @[Ray_AABB_1.scala 52:32]
  reg [31:0] cidx_0_1; // @[Ray_AABB_1.scala 53:45]
  reg [31:0] cidx_1_1; // @[Ray_AABB_1.scala 54:45]
  reg [31:0] rayid_temp; // @[Ray_AABB_1.scala 62:35]
  reg [31:0] hitT_temp; // @[Ray_AABB_1.scala 63:36]
  reg [31:0] valid_temp; // @[Ray_AABB_1.scala 65:35]
  reg [31:0] cidx_0_temp; // @[Ray_AABB_1.scala 72:48]
  reg [31:0] cidx_1_temp; // @[Ray_AABB_1.scala 73:48]
  wire  hi = ~io_ray_ood_x[31]; // @[common.scala 90:20]
  wire [30:0] lo = io_ray_ood_x[30:0]; // @[common.scala 90:30]
  wire  hi_2 = ~io_ray_ood_y[31]; // @[common.scala 90:20]
  wire [30:0] lo_2 = io_ray_ood_y[30:0]; // @[common.scala 90:30]
  wire  hi_4 = ~io_ray_ood_z[31]; // @[common.scala 90:20]
  wire [30:0] lo_4 = io_ray_ood_z[30:0]; // @[common.scala 90:30]
  reg [31:0] cidx_0_2; // @[Ray_AABB_1.scala 201:45]
  reg [31:0] cidx_1_2; // @[Ray_AABB_1.scala 202:45]
  reg [31:0] rayid_2; // @[Ray_AABB_1.scala 215:32]
  reg [31:0] hitT_2; // @[Ray_AABB_1.scala 216:33]
  reg [31:0] valid_2; // @[Ray_AABB_1.scala 218:32]
  reg [31:0] cmpMin0_1; // @[Ray_AABB_1.scala 225:28]
  reg [31:0] cmpMin0_2; // @[Ray_AABB_1.scala 226:28]
  reg [31:0] cmpMin0_3; // @[Ray_AABB_1.scala 227:28]
  reg [31:0] cmpMax0_1; // @[Ray_AABB_1.scala 228:28]
  reg [31:0] cmpMax0_2; // @[Ray_AABB_1.scala 229:28]
  reg [31:0] cmpMax0_3; // @[Ray_AABB_1.scala 230:28]
  reg [31:0] cmpMin1_1; // @[Ray_AABB_1.scala 231:28]
  reg [31:0] cmpMin1_2; // @[Ray_AABB_1.scala 232:28]
  reg [31:0] cmpMin1_3; // @[Ray_AABB_1.scala 233:28]
  reg [31:0] cmpMax1_1; // @[Ray_AABB_1.scala 234:28]
  reg [31:0] cmpMax1_2; // @[Ray_AABB_1.scala 235:28]
  reg [31:0] cmpMax1_3; // @[Ray_AABB_1.scala 236:28]
  wire  _T_24 = FCMP_1_io_actual_out; // @[Ray_AABB_1.scala 243:47]
  reg [31:0] c0Min_temp_1; // @[Ray_AABB_1.scala 319:31]
  reg [31:0] c0Min_temp_2; // @[Ray_AABB_1.scala 320:31]
  reg [31:0] c0Max_temp_1; // @[Ray_AABB_1.scala 321:31]
  reg [31:0] c0Max_temp_2; // @[Ray_AABB_1.scala 322:31]
  reg [31:0] c1Min_temp_1; // @[Ray_AABB_1.scala 323:31]
  reg [31:0] c1Min_temp_2; // @[Ray_AABB_1.scala 324:31]
  reg [31:0] c1Max_temp_1; // @[Ray_AABB_1.scala 325:31]
  reg [31:0] c1Max_temp_2; // @[Ray_AABB_1.scala 326:31]
  reg [31:0] cidx_0_3; // @[Ray_AABB_1.scala 328:45]
  reg [31:0] cidx_1_3; // @[Ray_AABB_1.scala 329:45]
  reg [31:0] hitT_3; // @[Ray_AABB_1.scala 343:49]
  reg [31:0] rayid_3; // @[Ray_AABB_1.scala 345:48]
  reg  valid_3; // @[Ray_AABB_1.scala 347:49]
  reg [31:0] c0Min; // @[Ray_AABB_1.scala 438:24]
  reg [31:0] c0Max; // @[Ray_AABB_1.scala 439:24]
  reg [31:0] c1Min; // @[Ray_AABB_1.scala 440:24]
  reg [31:0] c1Max; // @[Ray_AABB_1.scala 441:24]
  reg [31:0] cidx_0_4; // @[Ray_AABB_1.scala 443:45]
  reg [31:0] cidx_1_4; // @[Ray_AABB_1.scala 444:45]
  reg [31:0] hitT_4; // @[Ray_AABB_1.scala 458:49]
  reg [31:0] rayid_4; // @[Ray_AABB_1.scala 460:48]
  reg  valid_4; // @[Ray_AABB_1.scala 462:49]
  reg [31:0] rayid_5; // @[Ray_AABB_1.scala 510:48]
  reg [31:0] hitT_5; // @[Ray_AABB_1.scala 512:49]
  reg  valid_5; // @[Ray_AABB_1.scala 514:49]
  reg [31:0] cidx_0_5; // @[Ray_AABB_1.scala 519:45]
  reg [31:0] cidx_1_5; // @[Ray_AABB_1.scala 520:45]
  reg  swp; // @[Ray_AABB_1.scala 526:49]
  wire  _T_47 = FCMP_21_io_actual_out > 1'h0; // @[Ray_AABB_1.scala 572:36]
  wire  _T_48 = ~traverseChild0; // @[Ray_AABB_1.scala 580:10]
  wire  _T_49 = ~traverseChild1; // @[Ray_AABB_1.scala 580:29]
  wire  _T_60 = ~cidx_1_5[31]; // @[common.scala 100:25]
  wire  _T_62 = ~_T_60; // @[Ray_AABB_1.scala 600:32]
  wire [31:0] _GEN_28 = _T_60 ? $signed(cidx_1_5) : $signed(32'sh0); // @[Ray_AABB_1.scala 609:45 Ray_AABB_1.scala 615:29 Ray_AABB_1.scala 624:29]
  wire  _GEN_31 = ~_T_60 ? 1'h0 : _T_60; // @[Ray_AABB_1.scala 600:39 Ray_AABB_1.scala 604:37]
  wire [31:0] _GEN_33 = ~_T_60 ? $signed(32'sh0) : $signed(_GEN_28); // @[Ray_AABB_1.scala 600:39 Ray_AABB_1.scala 606:30]
  wire [31:0] _GEN_34 = ~_T_60 ? $signed(cidx_1_5) : $signed(32'sh0); // @[Ray_AABB_1.scala 600:39 Ray_AABB_1.scala 607:30]
  wire  _GEN_35 = ~_T_60 | _T_60; // @[Ray_AABB_1.scala 600:39 Ray_AABB_1.scala 608:32]
  wire  _T_73 = ~cidx_0_5[31]; // @[common.scala 100:25]
  wire  _T_75 = ~_T_73; // @[Ray_AABB_1.scala 639:32]
  wire [31:0] _GEN_39 = _T_73 ? $signed(cidx_0_5) : $signed(32'sh0); // @[Ray_AABB_1.scala 648:45 Ray_AABB_1.scala 654:33 Ray_AABB_1.scala 663:33]
  wire  _GEN_42 = ~_T_73 ? 1'h0 : _T_73; // @[Ray_AABB_1.scala 639:39 Ray_AABB_1.scala 643:41]
  wire [31:0] _GEN_44 = ~_T_73 ? $signed(32'sh0) : $signed(_GEN_39); // @[Ray_AABB_1.scala 639:39 Ray_AABB_1.scala 645:34]
  wire [31:0] _GEN_45 = ~_T_73 ? $signed(cidx_0_5) : $signed(32'sh0); // @[Ray_AABB_1.scala 639:39 Ray_AABB_1.scala 646:34]
  wire  _GEN_46 = ~_T_73 | _T_73; // @[Ray_AABB_1.scala 639:39 Ray_AABB_1.scala 647:36]
  wire [31:0] _GEN_49 = _T_60 ? $signed(cidx_0_5) : $signed(32'sh0); // @[Ray_AABB_1.scala 678:49 Ray_AABB_1.scala 683:32 Ray_AABB_1.scala 692:32]
  wire [31:0] _GEN_56 = _T_62 ? $signed(cidx_0_5) : $signed(_GEN_49); // @[Ray_AABB_1.scala 669:43 Ray_AABB_1.scala 674:32]
  wire [31:0] _GEN_61 = _T_73 ? $signed(cidx_1_5) : $signed(32'sh0); // @[Ray_AABB_1.scala 707:49 Ray_AABB_1.scala 712:32 Ray_AABB_1.scala 721:32]
  wire [31:0] _GEN_68 = _T_75 ? $signed(cidx_1_5) : $signed(_GEN_61); // @[Ray_AABB_1.scala 698:43 Ray_AABB_1.scala 703:32]
  wire  _GEN_71 = ~swp & valid_5 & _GEN_46; // @[Ray_AABB_1.scala 697:49 Ray_AABB_1.scala 746:38]
  wire  _GEN_73 = ~swp & valid_5 & _T_75; // @[Ray_AABB_1.scala 697:49 Ray_AABB_1.scala 748:41]
  wire  _GEN_74 = ~swp & valid_5 & _GEN_42; // @[Ray_AABB_1.scala 697:49 Ray_AABB_1.scala 749:39]
  wire [31:0] _GEN_75 = ~swp & valid_5 ? $signed(_GEN_68) : $signed(32'sh0); // @[Ray_AABB_1.scala 697:49 Ray_AABB_1.scala 750:32]
  wire [31:0] _GEN_76 = ~swp & valid_5 ? $signed(_GEN_44) : $signed(32'sh0); // @[Ray_AABB_1.scala 697:49 Ray_AABB_1.scala 751:32]
  wire [31:0] _GEN_77 = ~swp & valid_5 ? $signed(_GEN_45) : $signed(32'sh0); // @[Ray_AABB_1.scala 697:49 Ray_AABB_1.scala 752:32]
  wire  _GEN_78 = swp & valid_5 ? _GEN_35 : _GEN_71; // @[Ray_AABB_1.scala 668:43]
  wire  _GEN_80 = swp & valid_5 ? _T_62 : _GEN_73; // @[Ray_AABB_1.scala 668:43]
  wire  _GEN_81 = swp & valid_5 ? _GEN_31 : _GEN_74; // @[Ray_AABB_1.scala 668:43]
  wire [31:0] _GEN_82 = swp & valid_5 ? $signed(_GEN_56) : $signed(_GEN_75); // @[Ray_AABB_1.scala 668:43]
  wire [31:0] _GEN_83 = swp & valid_5 ? $signed(_GEN_33) : $signed(_GEN_76); // @[Ray_AABB_1.scala 668:43]
  wire [31:0] _GEN_84 = swp & valid_5 ? $signed(_GEN_34) : $signed(_GEN_77); // @[Ray_AABB_1.scala 668:43]
  wire  _GEN_85 = traverseChild0 & traverseChild1 & valid_5 & _GEN_78; // @[Ray_AABB_1.scala 667:84 Ray_AABB_1.scala 756:30]
  wire  _GEN_87 = traverseChild0 & traverseChild1 & valid_5 & _GEN_80; // @[Ray_AABB_1.scala 667:84 Ray_AABB_1.scala 758:33]
  wire  _GEN_88 = traverseChild0 & traverseChild1 & valid_5 & _GEN_81; // @[Ray_AABB_1.scala 667:84 Ray_AABB_1.scala 759:31]
  wire [31:0] _GEN_89 = traverseChild0 & traverseChild1 & valid_5 ? $signed(_GEN_82) : $signed(32'sh0); // @[Ray_AABB_1.scala 667:84 Ray_AABB_1.scala 760:24]
  wire [31:0] _GEN_90 = traverseChild0 & traverseChild1 & valid_5 ? $signed(_GEN_83) : $signed(32'sh0); // @[Ray_AABB_1.scala 667:84 Ray_AABB_1.scala 761:24]
  wire [31:0] _GEN_91 = traverseChild0 & traverseChild1 & valid_5 ? $signed(_GEN_84) : $signed(32'sh0); // @[Ray_AABB_1.scala 667:84 Ray_AABB_1.scala 762:24]
  wire  _GEN_92 = traverseChild0 & _T_49 & valid_5 ? _T_75 : _GEN_87; // @[Ray_AABB_1.scala 628:78]
  wire  _GEN_94 = traverseChild0 & _T_49 & valid_5 ? 1'h0 : _GEN_85; // @[Ray_AABB_1.scala 628:78]
  wire  _GEN_95 = traverseChild0 & _T_49 & valid_5 ? _GEN_42 : _GEN_88; // @[Ray_AABB_1.scala 628:78]
  wire [31:0] _GEN_96 = traverseChild0 & _T_49 & valid_5 ? $signed(32'sh0) : $signed(_GEN_89); // @[Ray_AABB_1.scala 628:78]
  wire [31:0] _GEN_97 = traverseChild0 & _T_49 & valid_5 ? $signed(_GEN_44) : $signed(_GEN_90); // @[Ray_AABB_1.scala 628:78]
  wire [31:0] _GEN_98 = traverseChild0 & _T_49 & valid_5 ? $signed(_GEN_45) : $signed(_GEN_91); // @[Ray_AABB_1.scala 628:78]
  wire  _GEN_99 = traverseChild0 & _T_49 & valid_5 ? _GEN_46 : _GEN_85; // @[Ray_AABB_1.scala 628:78]
  wire  _GEN_100 = _T_48 & traverseChild1 & valid_5 ? _T_62 : _GEN_92; // @[Ray_AABB_1.scala 589:74]
  wire  _GEN_102 = _T_48 & traverseChild1 & valid_5 ? 1'h0 : _GEN_94; // @[Ray_AABB_1.scala 589:74]
  wire  _GEN_103 = _T_48 & traverseChild1 & valid_5 ? _GEN_31 : _GEN_95; // @[Ray_AABB_1.scala 589:74]
  wire [31:0] _GEN_104 = _T_48 & traverseChild1 & valid_5 ? $signed(32'sh0) : $signed(_GEN_96); // @[Ray_AABB_1.scala 589:74]
  wire [31:0] _GEN_105 = _T_48 & traverseChild1 & valid_5 ? $signed(_GEN_33) : $signed(_GEN_97); // @[Ray_AABB_1.scala 589:74]
  wire [31:0] _GEN_106 = _T_48 & traverseChild1 & valid_5 ? $signed(_GEN_34) : $signed(_GEN_98); // @[Ray_AABB_1.scala 589:74]
  wire  _GEN_107 = _T_48 & traverseChild1 & valid_5 ? _GEN_35 : _GEN_99; // @[Ray_AABB_1.scala 589:74]
  MY_MULADD FADD_MUL_1 ( // @[Ray_AABB_1.scala 80:33]
    .clock(FADD_MUL_1_clock),
    .reset(FADD_MUL_1_reset),
    .io_a(FADD_MUL_1_io_a),
    .io_b(FADD_MUL_1_io_b),
    .io_c(FADD_MUL_1_io_c),
    .io_out(FADD_MUL_1_io_out)
  );
  MY_MULADD FADD_MUL_2 ( // @[Ray_AABB_1.scala 90:33]
    .clock(FADD_MUL_2_clock),
    .reset(FADD_MUL_2_reset),
    .io_a(FADD_MUL_2_io_a),
    .io_b(FADD_MUL_2_io_b),
    .io_c(FADD_MUL_2_io_c),
    .io_out(FADD_MUL_2_io_out)
  );
  MY_MULADD FADD_MUL_3 ( // @[Ray_AABB_1.scala 100:33]
    .clock(FADD_MUL_3_clock),
    .reset(FADD_MUL_3_reset),
    .io_a(FADD_MUL_3_io_a),
    .io_b(FADD_MUL_3_io_b),
    .io_c(FADD_MUL_3_io_c),
    .io_out(FADD_MUL_3_io_out)
  );
  MY_MULADD FADD_MUL_4 ( // @[Ray_AABB_1.scala 110:33]
    .clock(FADD_MUL_4_clock),
    .reset(FADD_MUL_4_reset),
    .io_a(FADD_MUL_4_io_a),
    .io_b(FADD_MUL_4_io_b),
    .io_c(FADD_MUL_4_io_c),
    .io_out(FADD_MUL_4_io_out)
  );
  MY_MULADD FADD_MUL_5 ( // @[Ray_AABB_1.scala 120:33]
    .clock(FADD_MUL_5_clock),
    .reset(FADD_MUL_5_reset),
    .io_a(FADD_MUL_5_io_a),
    .io_b(FADD_MUL_5_io_b),
    .io_c(FADD_MUL_5_io_c),
    .io_out(FADD_MUL_5_io_out)
  );
  MY_MULADD FADD_MUL_6 ( // @[Ray_AABB_1.scala 130:33]
    .clock(FADD_MUL_6_clock),
    .reset(FADD_MUL_6_reset),
    .io_a(FADD_MUL_6_io_a),
    .io_b(FADD_MUL_6_io_b),
    .io_c(FADD_MUL_6_io_c),
    .io_out(FADD_MUL_6_io_out)
  );
  MY_MULADD FADD_MUL_7 ( // @[Ray_AABB_1.scala 140:33]
    .clock(FADD_MUL_7_clock),
    .reset(FADD_MUL_7_reset),
    .io_a(FADD_MUL_7_io_a),
    .io_b(FADD_MUL_7_io_b),
    .io_c(FADD_MUL_7_io_c),
    .io_out(FADD_MUL_7_io_out)
  );
  MY_MULADD FADD_MUL_8 ( // @[Ray_AABB_1.scala 150:33]
    .clock(FADD_MUL_8_clock),
    .reset(FADD_MUL_8_reset),
    .io_a(FADD_MUL_8_io_a),
    .io_b(FADD_MUL_8_io_b),
    .io_c(FADD_MUL_8_io_c),
    .io_out(FADD_MUL_8_io_out)
  );
  MY_MULADD FADD_MUL_9 ( // @[Ray_AABB_1.scala 160:33]
    .clock(FADD_MUL_9_clock),
    .reset(FADD_MUL_9_reset),
    .io_a(FADD_MUL_9_io_a),
    .io_b(FADD_MUL_9_io_b),
    .io_c(FADD_MUL_9_io_c),
    .io_out(FADD_MUL_9_io_out)
  );
  MY_MULADD FADD_MUL_10 ( // @[Ray_AABB_1.scala 170:33]
    .clock(FADD_MUL_10_clock),
    .reset(FADD_MUL_10_reset),
    .io_a(FADD_MUL_10_io_a),
    .io_b(FADD_MUL_10_io_b),
    .io_c(FADD_MUL_10_io_c),
    .io_out(FADD_MUL_10_io_out)
  );
  MY_MULADD FADD_MUL_11 ( // @[Ray_AABB_1.scala 180:33]
    .clock(FADD_MUL_11_clock),
    .reset(FADD_MUL_11_reset),
    .io_a(FADD_MUL_11_io_a),
    .io_b(FADD_MUL_11_io_b),
    .io_c(FADD_MUL_11_io_c),
    .io_out(FADD_MUL_11_io_out)
  );
  MY_MULADD FADD_MUL_12 ( // @[Ray_AABB_1.scala 190:33]
    .clock(FADD_MUL_12_clock),
    .reset(FADD_MUL_12_reset),
    .io_a(FADD_MUL_12_io_a),
    .io_b(FADD_MUL_12_io_b),
    .io_c(FADD_MUL_12_io_c),
    .io_out(FADD_MUL_12_io_out)
  );
  ValExec_CompareRecF32_le FCMP_1 ( // @[Ray_AABB_1.scala 238:24]
    .io_a(FCMP_1_io_a),
    .io_b(FCMP_1_io_b),
    .io_actual_out(FCMP_1_io_actual_out)
  );
  ValExec_CompareRecF32_le FCMP_2 ( // @[Ray_AABB_1.scala 253:24]
    .io_a(FCMP_2_io_a),
    .io_b(FCMP_2_io_b),
    .io_actual_out(FCMP_2_io_actual_out)
  );
  ValExec_CompareRecF32_le FCMP_3 ( // @[Ray_AABB_1.scala 266:24]
    .io_a(FCMP_3_io_a),
    .io_b(FCMP_3_io_b),
    .io_actual_out(FCMP_3_io_actual_out)
  );
  ValExec_CompareRecF32_le FCMP_4 ( // @[Ray_AABB_1.scala 279:24]
    .io_a(FCMP_4_io_a),
    .io_b(FCMP_4_io_b),
    .io_actual_out(FCMP_4_io_actual_out)
  );
  ValExec_CompareRecF32_le FCMP_5 ( // @[Ray_AABB_1.scala 292:25]
    .io_a(FCMP_5_io_a),
    .io_b(FCMP_5_io_b),
    .io_actual_out(FCMP_5_io_actual_out)
  );
  ValExec_CompareRecF32_le FCMP_6 ( // @[Ray_AABB_1.scala 305:24]
    .io_a(FCMP_6_io_a),
    .io_b(FCMP_6_io_b),
    .io_actual_out(FCMP_6_io_actual_out)
  );
  ValExec_CompareRecF32_le FCMP_7 ( // @[Ray_AABB_1.scala 350:24]
    .io_a(FCMP_7_io_a),
    .io_b(FCMP_7_io_b),
    .io_actual_out(FCMP_7_io_actual_out)
  );
  ValExec_CompareRecF32_le FCMP_8 ( // @[Ray_AABB_1.scala 361:24]
    .io_a(FCMP_8_io_a),
    .io_b(FCMP_8_io_b),
    .io_actual_out(FCMP_8_io_actual_out)
  );
  ValExec_CompareRecF32_le FCMP_9 ( // @[Ray_AABB_1.scala 372:24]
    .io_a(FCMP_9_io_a),
    .io_b(FCMP_9_io_b),
    .io_actual_out(FCMP_9_io_actual_out)
  );
  ValExec_CompareRecF32_le FCMP_10 ( // @[Ray_AABB_1.scala 383:25]
    .io_a(FCMP_10_io_a),
    .io_b(FCMP_10_io_b),
    .io_actual_out(FCMP_10_io_actual_out)
  );
  ValExec_CompareRecF32_le FCMP_11 ( // @[Ray_AABB_1.scala 394:25]
    .io_a(FCMP_11_io_a),
    .io_b(FCMP_11_io_b),
    .io_actual_out(FCMP_11_io_actual_out)
  );
  ValExec_CompareRecF32_le FCMP_12 ( // @[Ray_AABB_1.scala 405:25]
    .io_a(FCMP_12_io_a),
    .io_b(FCMP_12_io_b),
    .io_actual_out(FCMP_12_io_actual_out)
  );
  ValExec_CompareRecF32_le FCMP_13 ( // @[Ray_AABB_1.scala 416:25]
    .io_a(FCMP_13_io_a),
    .io_b(FCMP_13_io_b),
    .io_actual_out(FCMP_13_io_actual_out)
  );
  ValExec_CompareRecF32_le FCMP_14 ( // @[Ray_AABB_1.scala 427:25]
    .io_a(FCMP_14_io_a),
    .io_b(FCMP_14_io_b),
    .io_actual_out(FCMP_14_io_actual_out)
  );
  ValExec_CompareRecF32_le FCMP_15 ( // @[Ray_AABB_1.scala 465:25]
    .io_a(FCMP_15_io_a),
    .io_b(FCMP_15_io_b),
    .io_actual_out(FCMP_15_io_actual_out)
  );
  ValExec_CompareRecF32_le FCMP_16 ( // @[Ray_AABB_1.scala 476:25]
    .io_a(FCMP_16_io_a),
    .io_b(FCMP_16_io_b),
    .io_actual_out(FCMP_16_io_actual_out)
  );
  ValExec_CompareRecF32_le FCMP_17 ( // @[Ray_AABB_1.scala 487:25]
    .io_a(FCMP_17_io_a),
    .io_b(FCMP_17_io_b),
    .io_actual_out(FCMP_17_io_actual_out)
  );
  ValExec_CompareRecF32_le FCMP_18 ( // @[Ray_AABB_1.scala 498:25]
    .io_a(FCMP_18_io_a),
    .io_b(FCMP_18_io_b),
    .io_actual_out(FCMP_18_io_actual_out)
  );
  ValExec_CompareRecF32_lt FCMP_19 ( // @[Ray_AABB_1.scala 541:25]
    .io_a(FCMP_19_io_a),
    .io_b(FCMP_19_io_b),
    .io_actual_out(FCMP_19_io_actual_out)
  );
  ValExec_CompareRecF32_lt FCMP_20 ( // @[Ray_AABB_1.scala 554:25]
    .io_a(FCMP_20_io_a),
    .io_b(FCMP_20_io_b),
    .io_actual_out(FCMP_20_io_actual_out)
  );
  ValExec_CompareRecF32_lt FCMP_21 ( // @[Ray_AABB_1.scala 567:25]
    .io_a(FCMP_21_io_a),
    .io_b(FCMP_21_io_b),
    .io_actual_out(FCMP_21_io_actual_out)
  );
  assign io_rayid_out = rayid_5; // @[Ray_AABB_1.scala 578:47]
  assign io_nodeIdx_0 = ~traverseChild0 & ~traverseChild1 & valid_5 ? $signed(32'sh0) : $signed(_GEN_104); // @[Ray_AABB_1.scala 580:69 Ray_AABB_1.scala 585:26]
  assign io_nodeIdx_1 = ~traverseChild0 & ~traverseChild1 & valid_5 ? $signed(32'sh0) : $signed(_GEN_105); // @[Ray_AABB_1.scala 580:69 Ray_AABB_1.scala 586:26]
  assign io_nodeIdx_2 = ~traverseChild0 & ~traverseChild1 & valid_5 ? $signed(32'sh0) : $signed(_GEN_106); // @[Ray_AABB_1.scala 580:69 Ray_AABB_1.scala 587:26]
  assign io_push = ~traverseChild0 & ~traverseChild1 & valid_5 ? 1'h0 : _GEN_102; // @[Ray_AABB_1.scala 580:69 Ray_AABB_1.scala 582:32]
  assign io_pop = ~traverseChild0 & ~traverseChild1 & valid_5; // @[Ray_AABB_1.scala 580:51]
  assign io_leaf = ~traverseChild0 & ~traverseChild1 & valid_5 ? 1'h0 : _GEN_100; // @[Ray_AABB_1.scala 580:69 Ray_AABB_1.scala 583:35]
  assign io_back = ~traverseChild0 & ~traverseChild1 & valid_5 ? 1'h0 : _GEN_103; // @[Ray_AABB_1.scala 580:69 Ray_AABB_1.scala 584:33]
  assign io_hitT_out = hitT_5; // @[Ray_AABB_1.scala 579:48]
  assign io_valid_out = ~traverseChild0 & ~traverseChild1 & valid_5 | _GEN_107; // @[Ray_AABB_1.scala 580:69 Ray_AABB_1.scala 588:28]
  assign FADD_MUL_1_clock = clock;
  assign FADD_MUL_1_reset = reset;
  assign FADD_MUL_1_io_a = io_bvh_n0xy_x; // @[Ray_AABB_1.scala 81:21]
  assign FADD_MUL_1_io_b = io_ray_idir_x; // @[Ray_AABB_1.scala 82:21]
  assign FADD_MUL_1_io_c = {hi,lo}; // @[Cat.scala 30:58]
  assign FADD_MUL_2_clock = clock;
  assign FADD_MUL_2_reset = reset;
  assign FADD_MUL_2_io_a = io_bvh_n0xy_y; // @[Ray_AABB_1.scala 91:21]
  assign FADD_MUL_2_io_b = io_ray_idir_x; // @[Ray_AABB_1.scala 92:21]
  assign FADD_MUL_2_io_c = {hi,lo}; // @[Cat.scala 30:58]
  assign FADD_MUL_3_clock = clock;
  assign FADD_MUL_3_reset = reset;
  assign FADD_MUL_3_io_a = io_bvh_n0xy_z; // @[Ray_AABB_1.scala 101:21]
  assign FADD_MUL_3_io_b = io_ray_idir_y; // @[Ray_AABB_1.scala 102:21]
  assign FADD_MUL_3_io_c = {hi_2,lo_2}; // @[Cat.scala 30:58]
  assign FADD_MUL_4_clock = clock;
  assign FADD_MUL_4_reset = reset;
  assign FADD_MUL_4_io_a = io_bvh_n0xy_w; // @[Ray_AABB_1.scala 111:21]
  assign FADD_MUL_4_io_b = io_ray_idir_y; // @[Ray_AABB_1.scala 112:21]
  assign FADD_MUL_4_io_c = {hi_2,lo_2}; // @[Cat.scala 30:58]
  assign FADD_MUL_5_clock = clock;
  assign FADD_MUL_5_reset = reset;
  assign FADD_MUL_5_io_a = io_bvh_nz_x; // @[Ray_AABB_1.scala 121:21]
  assign FADD_MUL_5_io_b = io_ray_idir_z; // @[Ray_AABB_1.scala 122:21]
  assign FADD_MUL_5_io_c = {hi_4,lo_4}; // @[Cat.scala 30:58]
  assign FADD_MUL_6_clock = clock;
  assign FADD_MUL_6_reset = reset;
  assign FADD_MUL_6_io_a = io_bvh_nz_y; // @[Ray_AABB_1.scala 131:21]
  assign FADD_MUL_6_io_b = io_ray_idir_z; // @[Ray_AABB_1.scala 132:21]
  assign FADD_MUL_6_io_c = {hi_4,lo_4}; // @[Cat.scala 30:58]
  assign FADD_MUL_7_clock = clock;
  assign FADD_MUL_7_reset = reset;
  assign FADD_MUL_7_io_a = io_bvh_n1xy_x; // @[Ray_AABB_1.scala 141:21]
  assign FADD_MUL_7_io_b = io_ray_idir_x; // @[Ray_AABB_1.scala 142:21]
  assign FADD_MUL_7_io_c = {hi,lo}; // @[Cat.scala 30:58]
  assign FADD_MUL_8_clock = clock;
  assign FADD_MUL_8_reset = reset;
  assign FADD_MUL_8_io_a = io_bvh_n1xy_y; // @[Ray_AABB_1.scala 151:21]
  assign FADD_MUL_8_io_b = io_ray_idir_x; // @[Ray_AABB_1.scala 152:21]
  assign FADD_MUL_8_io_c = {hi,lo}; // @[Cat.scala 30:58]
  assign FADD_MUL_9_clock = clock;
  assign FADD_MUL_9_reset = reset;
  assign FADD_MUL_9_io_a = io_bvh_n1xy_z; // @[Ray_AABB_1.scala 161:21]
  assign FADD_MUL_9_io_b = io_ray_idir_y; // @[Ray_AABB_1.scala 162:21]
  assign FADD_MUL_9_io_c = {hi_2,lo_2}; // @[Cat.scala 30:58]
  assign FADD_MUL_10_clock = clock;
  assign FADD_MUL_10_reset = reset;
  assign FADD_MUL_10_io_a = io_bvh_n1xy_w; // @[Ray_AABB_1.scala 171:22]
  assign FADD_MUL_10_io_b = io_ray_idir_y; // @[Ray_AABB_1.scala 172:22]
  assign FADD_MUL_10_io_c = {hi_2,lo_2}; // @[Cat.scala 30:58]
  assign FADD_MUL_11_clock = clock;
  assign FADD_MUL_11_reset = reset;
  assign FADD_MUL_11_io_a = io_bvh_nz_z; // @[Ray_AABB_1.scala 181:22]
  assign FADD_MUL_11_io_b = io_ray_idir_z; // @[Ray_AABB_1.scala 182:22]
  assign FADD_MUL_11_io_c = {hi_4,lo_4}; // @[Cat.scala 30:58]
  assign FADD_MUL_12_clock = clock;
  assign FADD_MUL_12_reset = reset;
  assign FADD_MUL_12_io_a = io_bvh_nz_w; // @[Ray_AABB_1.scala 191:22]
  assign FADD_MUL_12_io_b = io_ray_idir_z; // @[Ray_AABB_1.scala 192:22]
  assign FADD_MUL_12_io_c = {hi_4,lo_4}; // @[Cat.scala 30:58]
  assign FCMP_1_io_a = c0lox; // @[Ray_AABB_1.scala 239:21]
  assign FCMP_1_io_b = c0hix; // @[Ray_AABB_1.scala 240:21]
  assign FCMP_2_io_a = c0loy; // @[Ray_AABB_1.scala 254:21]
  assign FCMP_2_io_b = c0hiy; // @[Ray_AABB_1.scala 255:21]
  assign FCMP_3_io_a = c0loz; // @[Ray_AABB_1.scala 267:21]
  assign FCMP_3_io_b = c0hiz; // @[Ray_AABB_1.scala 268:21]
  assign FCMP_4_io_a = c1lox; // @[Ray_AABB_1.scala 280:21]
  assign FCMP_4_io_b = c1hix; // @[Ray_AABB_1.scala 281:21]
  assign FCMP_5_io_a = c1loy; // @[Ray_AABB_1.scala 293:21]
  assign FCMP_5_io_b = c1hiy; // @[Ray_AABB_1.scala 294:21]
  assign FCMP_6_io_a = c1loz; // @[Ray_AABB_1.scala 306:21]
  assign FCMP_6_io_b = c1hiz; // @[Ray_AABB_1.scala 307:21]
  assign FCMP_7_io_a = cmpMin0_1; // @[Ray_AABB_1.scala 351:21]
  assign FCMP_7_io_b = cmpMin0_2; // @[Ray_AABB_1.scala 352:21]
  assign FCMP_8_io_a = cmpMin0_3; // @[Ray_AABB_1.scala 362:21]
  assign FCMP_8_io_b = 32'h0; // @[Ray_AABB_1.scala 363:21]
  assign FCMP_9_io_a = cmpMax0_1; // @[Ray_AABB_1.scala 373:21]
  assign FCMP_9_io_b = cmpMax0_2; // @[Ray_AABB_1.scala 374:21]
  assign FCMP_10_io_a = cmpMax0_3; // @[Ray_AABB_1.scala 384:22]
  assign FCMP_10_io_b = hitT_2; // @[Ray_AABB_1.scala 385:22]
  assign FCMP_11_io_a = cmpMin1_1; // @[Ray_AABB_1.scala 395:22]
  assign FCMP_11_io_b = cmpMin1_2; // @[Ray_AABB_1.scala 396:22]
  assign FCMP_12_io_a = cmpMin1_3; // @[Ray_AABB_1.scala 406:22]
  assign FCMP_12_io_b = 32'h0; // @[Ray_AABB_1.scala 407:22]
  assign FCMP_13_io_a = cmpMax1_1; // @[Ray_AABB_1.scala 417:22]
  assign FCMP_13_io_b = cmpMax1_2; // @[Ray_AABB_1.scala 418:22]
  assign FCMP_14_io_a = cmpMax1_3; // @[Ray_AABB_1.scala 428:22]
  assign FCMP_14_io_b = hitT_2; // @[Ray_AABB_1.scala 429:22]
  assign FCMP_15_io_a = c0Min_temp_1; // @[Ray_AABB_1.scala 466:22]
  assign FCMP_15_io_b = c0Min_temp_2; // @[Ray_AABB_1.scala 467:22]
  assign FCMP_16_io_a = c0Max_temp_1; // @[Ray_AABB_1.scala 477:22]
  assign FCMP_16_io_b = c0Max_temp_2; // @[Ray_AABB_1.scala 478:22]
  assign FCMP_17_io_a = c1Min_temp_1; // @[Ray_AABB_1.scala 488:22]
  assign FCMP_17_io_b = c1Min_temp_2; // @[Ray_AABB_1.scala 489:22]
  assign FCMP_18_io_a = c1Max_temp_1; // @[Ray_AABB_1.scala 499:22]
  assign FCMP_18_io_b = c1Max_temp_2; // @[Ray_AABB_1.scala 500:22]
  assign FCMP_19_io_a = c0Max; // @[Ray_AABB_1.scala 542:22]
  assign FCMP_19_io_b = c0Min; // @[Ray_AABB_1.scala 543:22]
  assign FCMP_20_io_a = c1Max; // @[Ray_AABB_1.scala 555:22]
  assign FCMP_20_io_b = c1Min; // @[Ray_AABB_1.scala 556:22]
  assign FCMP_21_io_a = c1Min; // @[Ray_AABB_1.scala 568:22]
  assign FCMP_21_io_b = c0Min; // @[Ray_AABB_1.scala 569:22]
  always @(posedge clock) begin
    if (reset) begin // @[Ray_AABB_1.scala 32:33]
      traverseChild0 <= 1'h0; // @[Ray_AABB_1.scala 32:33]
    end else if (FCMP_19_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 546:42]
      traverseChild0 <= 1'h0; // @[Ray_AABB_1.scala 547:28]
    end else begin
      traverseChild0 <= 1'h1; // @[Ray_AABB_1.scala 549:28]
    end
    if (reset) begin // @[Ray_AABB_1.scala 33:33]
      traverseChild1 <= 1'h0; // @[Ray_AABB_1.scala 33:33]
    end else if (FCMP_20_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 559:42]
      traverseChild1 <= 1'h0; // @[Ray_AABB_1.scala 560:28]
    end else begin
      traverseChild1 <= 1'h1; // @[Ray_AABB_1.scala 562:28]
    end
    if (reset) begin // @[Ray_AABB_1.scala 35:34]
      c0lox <= 32'h0; // @[Ray_AABB_1.scala 35:34]
    end else begin
      c0lox <= FADD_MUL_1_io_out; // @[Ray_AABB_1.scala 88:37]
    end
    if (reset) begin // @[Ray_AABB_1.scala 36:34]
      c0hix <= 32'h0; // @[Ray_AABB_1.scala 36:34]
    end else begin
      c0hix <= FADD_MUL_2_io_out; // @[Ray_AABB_1.scala 98:37]
    end
    if (reset) begin // @[Ray_AABB_1.scala 37:34]
      c0loy <= 32'h0; // @[Ray_AABB_1.scala 37:34]
    end else begin
      c0loy <= FADD_MUL_3_io_out; // @[Ray_AABB_1.scala 108:37]
    end
    if (reset) begin // @[Ray_AABB_1.scala 38:33]
      c0hiy <= 32'h0; // @[Ray_AABB_1.scala 38:33]
    end else begin
      c0hiy <= FADD_MUL_4_io_out; // @[Ray_AABB_1.scala 118:37]
    end
    if (reset) begin // @[Ray_AABB_1.scala 39:34]
      c0loz <= 32'h0; // @[Ray_AABB_1.scala 39:34]
    end else begin
      c0loz <= FADD_MUL_5_io_out; // @[Ray_AABB_1.scala 128:37]
    end
    if (reset) begin // @[Ray_AABB_1.scala 40:34]
      c0hiz <= 32'h0; // @[Ray_AABB_1.scala 40:34]
    end else begin
      c0hiz <= FADD_MUL_6_io_out; // @[Ray_AABB_1.scala 138:37]
    end
    if (reset) begin // @[Ray_AABB_1.scala 42:34]
      c1lox <= 32'h0; // @[Ray_AABB_1.scala 42:34]
    end else begin
      c1lox <= FADD_MUL_7_io_out; // @[Ray_AABB_1.scala 148:37]
    end
    if (reset) begin // @[Ray_AABB_1.scala 43:34]
      c1hix <= 32'h0; // @[Ray_AABB_1.scala 43:34]
    end else begin
      c1hix <= FADD_MUL_8_io_out; // @[Ray_AABB_1.scala 158:37]
    end
    if (reset) begin // @[Ray_AABB_1.scala 44:34]
      c1loy <= 32'h0; // @[Ray_AABB_1.scala 44:34]
    end else begin
      c1loy <= FADD_MUL_9_io_out; // @[Ray_AABB_1.scala 168:37]
    end
    if (reset) begin // @[Ray_AABB_1.scala 45:34]
      c1hiy <= 32'h0; // @[Ray_AABB_1.scala 45:34]
    end else begin
      c1hiy <= FADD_MUL_10_io_out; // @[Ray_AABB_1.scala 178:37]
    end
    if (reset) begin // @[Ray_AABB_1.scala 46:34]
      c1loz <= 32'h0; // @[Ray_AABB_1.scala 46:34]
    end else begin
      c1loz <= FADD_MUL_11_io_out; // @[Ray_AABB_1.scala 188:37]
    end
    if (reset) begin // @[Ray_AABB_1.scala 47:34]
      c1hiz <= 32'h0; // @[Ray_AABB_1.scala 47:34]
    end else begin
      c1hiz <= FADD_MUL_12_io_out; // @[Ray_AABB_1.scala 198:37]
    end
    if (reset) begin // @[Ray_AABB_1.scala 49:32]
      rayid_1 <= 32'h0; // @[Ray_AABB_1.scala 49:32]
    end else begin
      rayid_1 <= io_rayid; // @[Ray_AABB_1.scala 55:41]
    end
    if (reset) begin // @[Ray_AABB_1.scala 50:33]
      hitT_1 <= 32'h0; // @[Ray_AABB_1.scala 50:33]
    end else begin
      hitT_1 <= io_ray_hitT; // @[Ray_AABB_1.scala 57:43]
    end
    if (reset) begin // @[Ray_AABB_1.scala 52:32]
      valid_1 <= 32'h0; // @[Ray_AABB_1.scala 52:32]
    end else begin
      valid_1 <= {{31'd0}, io_valid_en}; // @[Ray_AABB_1.scala 58:42]
    end
    if (reset) begin // @[Ray_AABB_1.scala 53:45]
      cidx_0_1 <= 32'sh0; // @[Ray_AABB_1.scala 53:45]
    end else begin
      cidx_0_1 <= io_bvh_temp_x; // @[Ray_AABB_1.scala 59:44]
    end
    if (reset) begin // @[Ray_AABB_1.scala 54:45]
      cidx_1_1 <= 32'sh0; // @[Ray_AABB_1.scala 54:45]
    end else begin
      cidx_1_1 <= io_bvh_temp_y; // @[Ray_AABB_1.scala 60:44]
    end
    if (reset) begin // @[Ray_AABB_1.scala 62:35]
      rayid_temp <= 32'h0; // @[Ray_AABB_1.scala 62:35]
    end else begin
      rayid_temp <= rayid_1; // @[Ray_AABB_1.scala 69:31]
    end
    if (reset) begin // @[Ray_AABB_1.scala 63:36]
      hitT_temp <= 32'h0; // @[Ray_AABB_1.scala 63:36]
    end else begin
      hitT_temp <= hitT_1; // @[Ray_AABB_1.scala 67:32]
    end
    if (reset) begin // @[Ray_AABB_1.scala 65:35]
      valid_temp <= 32'h0; // @[Ray_AABB_1.scala 65:35]
    end else begin
      valid_temp <= valid_1; // @[Ray_AABB_1.scala 70:32]
    end
    if (reset) begin // @[Ray_AABB_1.scala 72:48]
      cidx_0_temp <= 32'sh0; // @[Ray_AABB_1.scala 72:48]
    end else begin
      cidx_0_temp <= cidx_0_1; // @[Ray_AABB_1.scala 76:41]
    end
    if (reset) begin // @[Ray_AABB_1.scala 73:48]
      cidx_1_temp <= 32'sh0; // @[Ray_AABB_1.scala 73:48]
    end else begin
      cidx_1_temp <= cidx_1_1; // @[Ray_AABB_1.scala 77:41]
    end
    if (reset) begin // @[Ray_AABB_1.scala 201:45]
      cidx_0_2 <= 32'sh0; // @[Ray_AABB_1.scala 201:45]
    end else begin
      cidx_0_2 <= cidx_0_temp; // @[Ray_AABB_1.scala 208:38]
    end
    if (reset) begin // @[Ray_AABB_1.scala 202:45]
      cidx_1_2 <= 32'sh0; // @[Ray_AABB_1.scala 202:45]
    end else begin
      cidx_1_2 <= cidx_1_temp; // @[Ray_AABB_1.scala 209:38]
    end
    if (reset) begin // @[Ray_AABB_1.scala 215:32]
      rayid_2 <= 32'h0; // @[Ray_AABB_1.scala 215:32]
    end else begin
      rayid_2 <= rayid_temp; // @[Ray_AABB_1.scala 222:28]
    end
    if (reset) begin // @[Ray_AABB_1.scala 216:33]
      hitT_2 <= 32'h0; // @[Ray_AABB_1.scala 216:33]
    end else begin
      hitT_2 <= hitT_temp; // @[Ray_AABB_1.scala 220:29]
    end
    if (reset) begin // @[Ray_AABB_1.scala 218:32]
      valid_2 <= 32'h0; // @[Ray_AABB_1.scala 218:32]
    end else begin
      valid_2 <= valid_temp; // @[Ray_AABB_1.scala 223:29]
    end
    if (reset) begin // @[Ray_AABB_1.scala 225:28]
      cmpMin0_1 <= 32'h0; // @[Ray_AABB_1.scala 225:28]
    end else if (FCMP_1_io_actual_out) begin // @[Ray_AABB_1.scala 243:25]
      cmpMin0_1 <= c0lox;
    end else begin
      cmpMin0_1 <= c0hix;
    end
    if (reset) begin // @[Ray_AABB_1.scala 226:28]
      cmpMin0_2 <= 32'h0; // @[Ray_AABB_1.scala 226:28]
    end else if (FCMP_2_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 258:41]
      cmpMin0_2 <= c0loy; // @[Ray_AABB_1.scala 259:23]
    end else begin
      cmpMin0_2 <= c0hiy; // @[Ray_AABB_1.scala 262:23]
    end
    if (reset) begin // @[Ray_AABB_1.scala 227:28]
      cmpMin0_3 <= 32'h0; // @[Ray_AABB_1.scala 227:28]
    end else if (FCMP_3_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 271:41]
      cmpMin0_3 <= c0loz; // @[Ray_AABB_1.scala 272:23]
    end else begin
      cmpMin0_3 <= c0hiz; // @[Ray_AABB_1.scala 275:23]
    end
    if (reset) begin // @[Ray_AABB_1.scala 228:28]
      cmpMax0_1 <= 32'h0; // @[Ray_AABB_1.scala 228:28]
    end else if (_T_24) begin // @[Ray_AABB_1.scala 244:25]
      cmpMax0_1 <= c0hix;
    end else begin
      cmpMax0_1 <= c0lox;
    end
    if (reset) begin // @[Ray_AABB_1.scala 229:28]
      cmpMax0_2 <= 32'h0; // @[Ray_AABB_1.scala 229:28]
    end else if (FCMP_2_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 258:41]
      cmpMax0_2 <= c0hiy; // @[Ray_AABB_1.scala 260:23]
    end else begin
      cmpMax0_2 <= c0loy; // @[Ray_AABB_1.scala 263:23]
    end
    if (reset) begin // @[Ray_AABB_1.scala 230:28]
      cmpMax0_3 <= 32'h0; // @[Ray_AABB_1.scala 230:28]
    end else if (FCMP_3_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 271:41]
      cmpMax0_3 <= c0hiz; // @[Ray_AABB_1.scala 273:23]
    end else begin
      cmpMax0_3 <= c0loz; // @[Ray_AABB_1.scala 276:23]
    end
    if (reset) begin // @[Ray_AABB_1.scala 231:28]
      cmpMin1_1 <= 32'h0; // @[Ray_AABB_1.scala 231:28]
    end else if (FCMP_4_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 284:41]
      cmpMin1_1 <= c1lox; // @[Ray_AABB_1.scala 285:23]
    end else begin
      cmpMin1_1 <= c1hix; // @[Ray_AABB_1.scala 288:23]
    end
    if (reset) begin // @[Ray_AABB_1.scala 232:28]
      cmpMin1_2 <= 32'h0; // @[Ray_AABB_1.scala 232:28]
    end else if (FCMP_5_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 297:41]
      cmpMin1_2 <= c1loy; // @[Ray_AABB_1.scala 298:23]
    end else begin
      cmpMin1_2 <= c1hiy; // @[Ray_AABB_1.scala 301:23]
    end
    if (reset) begin // @[Ray_AABB_1.scala 233:28]
      cmpMin1_3 <= 32'h0; // @[Ray_AABB_1.scala 233:28]
    end else if (FCMP_6_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 310:41]
      cmpMin1_3 <= c1loz; // @[Ray_AABB_1.scala 311:23]
    end else begin
      cmpMin1_3 <= c1hiz; // @[Ray_AABB_1.scala 314:23]
    end
    if (reset) begin // @[Ray_AABB_1.scala 234:28]
      cmpMax1_1 <= 32'h0; // @[Ray_AABB_1.scala 234:28]
    end else if (FCMP_4_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 284:41]
      cmpMax1_1 <= c1hix; // @[Ray_AABB_1.scala 286:23]
    end else begin
      cmpMax1_1 <= c1lox; // @[Ray_AABB_1.scala 289:23]
    end
    if (reset) begin // @[Ray_AABB_1.scala 235:28]
      cmpMax1_2 <= 32'h0; // @[Ray_AABB_1.scala 235:28]
    end else if (FCMP_5_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 297:41]
      cmpMax1_2 <= c1hiy; // @[Ray_AABB_1.scala 299:23]
    end else begin
      cmpMax1_2 <= c1loy; // @[Ray_AABB_1.scala 302:23]
    end
    if (reset) begin // @[Ray_AABB_1.scala 236:28]
      cmpMax1_3 <= 32'h0; // @[Ray_AABB_1.scala 236:28]
    end else if (FCMP_6_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 310:41]
      cmpMax1_3 <= c1hiz; // @[Ray_AABB_1.scala 312:23]
    end else begin
      cmpMax1_3 <= c1loz; // @[Ray_AABB_1.scala 315:23]
    end
    if (reset) begin // @[Ray_AABB_1.scala 319:31]
      c0Min_temp_1 <= 32'h0; // @[Ray_AABB_1.scala 319:31]
    end else if (FCMP_7_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 355:41]
      c0Min_temp_1 <= cmpMin0_2; // @[Ray_AABB_1.scala 356:26]
    end else begin
      c0Min_temp_1 <= cmpMin0_1; // @[Ray_AABB_1.scala 358:26]
    end
    if (reset) begin // @[Ray_AABB_1.scala 320:31]
      c0Min_temp_2 <= 32'h0; // @[Ray_AABB_1.scala 320:31]
    end else if (FCMP_8_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 366:41]
      c0Min_temp_2 <= 32'h0; // @[Ray_AABB_1.scala 367:26]
    end else begin
      c0Min_temp_2 <= cmpMin0_3; // @[Ray_AABB_1.scala 369:26]
    end
    if (reset) begin // @[Ray_AABB_1.scala 321:31]
      c0Max_temp_1 <= 32'h0; // @[Ray_AABB_1.scala 321:31]
    end else if (FCMP_9_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 377:41]
      c0Max_temp_1 <= cmpMax0_1; // @[Ray_AABB_1.scala 378:26]
    end else begin
      c0Max_temp_1 <= cmpMax0_2; // @[Ray_AABB_1.scala 380:26]
    end
    if (reset) begin // @[Ray_AABB_1.scala 322:31]
      c0Max_temp_2 <= 32'h0; // @[Ray_AABB_1.scala 322:31]
    end else if (FCMP_10_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 388:42]
      c0Max_temp_2 <= cmpMax0_3; // @[Ray_AABB_1.scala 389:26]
    end else begin
      c0Max_temp_2 <= hitT_2; // @[Ray_AABB_1.scala 391:26]
    end
    if (reset) begin // @[Ray_AABB_1.scala 323:31]
      c1Min_temp_1 <= 32'h0; // @[Ray_AABB_1.scala 323:31]
    end else if (FCMP_11_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 399:42]
      c1Min_temp_1 <= cmpMin1_2; // @[Ray_AABB_1.scala 400:26]
    end else begin
      c1Min_temp_1 <= cmpMin1_1; // @[Ray_AABB_1.scala 402:26]
    end
    if (reset) begin // @[Ray_AABB_1.scala 324:31]
      c1Min_temp_2 <= 32'h0; // @[Ray_AABB_1.scala 324:31]
    end else if (FCMP_12_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 410:42]
      c1Min_temp_2 <= 32'h0; // @[Ray_AABB_1.scala 411:26]
    end else begin
      c1Min_temp_2 <= cmpMin1_3; // @[Ray_AABB_1.scala 413:26]
    end
    if (reset) begin // @[Ray_AABB_1.scala 325:31]
      c1Max_temp_1 <= 32'h0; // @[Ray_AABB_1.scala 325:31]
    end else if (FCMP_13_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 421:42]
      c1Max_temp_1 <= cmpMax1_1; // @[Ray_AABB_1.scala 422:26]
    end else begin
      c1Max_temp_1 <= cmpMax1_2; // @[Ray_AABB_1.scala 424:26]
    end
    if (reset) begin // @[Ray_AABB_1.scala 326:31]
      c1Max_temp_2 <= 32'h0; // @[Ray_AABB_1.scala 326:31]
    end else if (FCMP_14_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 432:42]
      c1Max_temp_2 <= cmpMax1_3; // @[Ray_AABB_1.scala 433:26]
    end else begin
      c1Max_temp_2 <= hitT_2; // @[Ray_AABB_1.scala 435:26]
    end
    if (reset) begin // @[Ray_AABB_1.scala 328:45]
      cidx_0_3 <= 32'sh0; // @[Ray_AABB_1.scala 328:45]
    end else begin
      cidx_0_3 <= cidx_0_2; // @[Ray_AABB_1.scala 336:38]
    end
    if (reset) begin // @[Ray_AABB_1.scala 329:45]
      cidx_1_3 <= 32'sh0; // @[Ray_AABB_1.scala 329:45]
    end else begin
      cidx_1_3 <= cidx_1_2; // @[Ray_AABB_1.scala 337:38]
    end
    if (reset) begin // @[Ray_AABB_1.scala 343:49]
      hitT_3 <= 32'h0; // @[Ray_AABB_1.scala 343:49]
    end else begin
      hitT_3 <= hitT_2; // @[Ray_AABB_1.scala 344:42]
    end
    if (reset) begin // @[Ray_AABB_1.scala 345:48]
      rayid_3 <= 32'h0; // @[Ray_AABB_1.scala 345:48]
    end else begin
      rayid_3 <= rayid_2; // @[Ray_AABB_1.scala 346:41]
    end
    if (reset) begin // @[Ray_AABB_1.scala 347:49]
      valid_3 <= 1'h0; // @[Ray_AABB_1.scala 347:49]
    end else begin
      valid_3 <= valid_2[0]; // @[Ray_AABB_1.scala 348:41]
    end
    if (reset) begin // @[Ray_AABB_1.scala 438:24]
      c0Min <= 32'h0; // @[Ray_AABB_1.scala 438:24]
    end else if (FCMP_15_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 470:42]
      c0Min <= c0Min_temp_2; // @[Ray_AABB_1.scala 471:19]
    end else begin
      c0Min <= c0Min_temp_1; // @[Ray_AABB_1.scala 473:19]
    end
    if (reset) begin // @[Ray_AABB_1.scala 439:24]
      c0Max <= 32'h0; // @[Ray_AABB_1.scala 439:24]
    end else if (FCMP_16_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 481:42]
      c0Max <= c0Max_temp_1; // @[Ray_AABB_1.scala 482:19]
    end else begin
      c0Max <= c0Max_temp_2; // @[Ray_AABB_1.scala 484:19]
    end
    if (reset) begin // @[Ray_AABB_1.scala 440:24]
      c1Min <= 32'h0; // @[Ray_AABB_1.scala 440:24]
    end else if (FCMP_17_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 492:42]
      c1Min <= c1Min_temp_2; // @[Ray_AABB_1.scala 493:19]
    end else begin
      c1Min <= c1Min_temp_1; // @[Ray_AABB_1.scala 495:19]
    end
    if (reset) begin // @[Ray_AABB_1.scala 441:24]
      c1Max <= 32'h0; // @[Ray_AABB_1.scala 441:24]
    end else if (FCMP_18_io_actual_out > 1'h0) begin // @[Ray_AABB_1.scala 503:42]
      c1Max <= c1Max_temp_1; // @[Ray_AABB_1.scala 504:19]
    end else begin
      c1Max <= c1Max_temp_2; // @[Ray_AABB_1.scala 506:19]
    end
    if (reset) begin // @[Ray_AABB_1.scala 443:45]
      cidx_0_4 <= 32'sh0; // @[Ray_AABB_1.scala 443:45]
    end else begin
      cidx_0_4 <= cidx_0_3; // @[Ray_AABB_1.scala 451:38]
    end
    if (reset) begin // @[Ray_AABB_1.scala 444:45]
      cidx_1_4 <= 32'sh0; // @[Ray_AABB_1.scala 444:45]
    end else begin
      cidx_1_4 <= cidx_1_3; // @[Ray_AABB_1.scala 452:38]
    end
    if (reset) begin // @[Ray_AABB_1.scala 458:49]
      hitT_4 <= 32'h0; // @[Ray_AABB_1.scala 458:49]
    end else begin
      hitT_4 <= hitT_3; // @[Ray_AABB_1.scala 459:43]
    end
    if (reset) begin // @[Ray_AABB_1.scala 460:48]
      rayid_4 <= 32'h0; // @[Ray_AABB_1.scala 460:48]
    end else begin
      rayid_4 <= rayid_3; // @[Ray_AABB_1.scala 461:42]
    end
    if (reset) begin // @[Ray_AABB_1.scala 462:49]
      valid_4 <= 1'h0; // @[Ray_AABB_1.scala 462:49]
    end else begin
      valid_4 <= valid_3; // @[Ray_AABB_1.scala 463:41]
    end
    if (reset) begin // @[Ray_AABB_1.scala 510:48]
      rayid_5 <= 32'h0; // @[Ray_AABB_1.scala 510:48]
    end else begin
      rayid_5 <= rayid_4; // @[Ray_AABB_1.scala 511:42]
    end
    if (reset) begin // @[Ray_AABB_1.scala 512:49]
      hitT_5 <= 32'h0; // @[Ray_AABB_1.scala 512:49]
    end else begin
      hitT_5 <= hitT_4; // @[Ray_AABB_1.scala 513:42]
    end
    if (reset) begin // @[Ray_AABB_1.scala 514:49]
      valid_5 <= 1'h0; // @[Ray_AABB_1.scala 514:49]
    end else begin
      valid_5 <= valid_4; // @[Ray_AABB_1.scala 515:41]
    end
    if (reset) begin // @[Ray_AABB_1.scala 519:45]
      cidx_0_5 <= 32'sh0; // @[Ray_AABB_1.scala 519:45]
    end else begin
      cidx_0_5 <= cidx_0_4; // @[Ray_AABB_1.scala 531:38]
    end
    if (reset) begin // @[Ray_AABB_1.scala 520:45]
      cidx_1_5 <= 32'sh0; // @[Ray_AABB_1.scala 520:45]
    end else begin
      cidx_1_5 <= cidx_1_4; // @[Ray_AABB_1.scala 532:38]
    end
    if (reset) begin // @[Ray_AABB_1.scala 526:49]
      swp <= 1'h0; // @[Ray_AABB_1.scala 526:49]
    end else begin
      swp <= _T_47;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  traverseChild0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  traverseChild1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  c0lox = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  c0hix = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  c0loy = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  c0hiy = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  c0loz = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  c0hiz = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  c1lox = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  c1hix = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  c1loy = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  c1hiy = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  c1loz = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  c1hiz = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  rayid_1 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  hitT_1 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  valid_1 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  cidx_0_1 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  cidx_1_1 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  rayid_temp = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  hitT_temp = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  valid_temp = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  cidx_0_temp = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  cidx_1_temp = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  cidx_0_2 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  cidx_1_2 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  rayid_2 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  hitT_2 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  valid_2 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  cmpMin0_1 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  cmpMin0_2 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  cmpMin0_3 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  cmpMax0_1 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  cmpMax0_2 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  cmpMax0_3 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  cmpMin1_1 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  cmpMin1_2 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  cmpMin1_3 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  cmpMax1_1 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  cmpMax1_2 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  cmpMax1_3 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  c0Min_temp_1 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  c0Min_temp_2 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  c0Max_temp_1 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  c0Max_temp_2 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  c1Min_temp_1 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  c1Min_temp_2 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  c1Max_temp_1 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  c1Max_temp_2 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  cidx_0_3 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  cidx_1_3 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  hitT_3 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  rayid_3 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  valid_3 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  c0Min = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  c0Max = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  c1Min = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  c1Max = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  cidx_0_4 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  cidx_1_4 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  hitT_4 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  rayid_4 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  valid_4 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  rayid_5 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  hitT_5 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  valid_5 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  cidx_0_5 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  cidx_1_5 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  swp = _RAND_68[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FIFO(
  input         clock,
  input         reset,
  input  [31:0] io_datain,
  output [31:0] io_dataout,
  input         io_wr,
  input         io_rd,
  output        io_empty
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] mem [0:34]; // @[FIFO.scala 23:16]
  wire [31:0] mem_MPORT_data; // @[FIFO.scala 23:16]
  wire [5:0] mem_MPORT_addr; // @[FIFO.scala 23:16]
  wire [31:0] mem_MPORT_3_data; // @[FIFO.scala 23:16]
  wire [5:0] mem_MPORT_3_addr; // @[FIFO.scala 23:16]
  wire [31:0] mem_MPORT_1_data; // @[FIFO.scala 23:16]
  wire [5:0] mem_MPORT_1_addr; // @[FIFO.scala 23:16]
  wire  mem_MPORT_1_mask; // @[FIFO.scala 23:16]
  wire  mem_MPORT_1_en; // @[FIFO.scala 23:16]
  wire [31:0] mem_MPORT_2_data; // @[FIFO.scala 23:16]
  wire [5:0] mem_MPORT_2_addr; // @[FIFO.scala 23:16]
  wire  mem_MPORT_2_mask; // @[FIFO.scala 23:16]
  wire  mem_MPORT_2_en; // @[FIFO.scala 23:16]
  reg [31:0] count; // @[FIFO.scala 22:22]
  reg [31:0] wPointer; // @[FIFO.scala 24:25]
  reg [31:0] rPointer; // @[FIFO.scala 25:25]
  reg [31:0] dataout; // @[FIFO.scala 26:24]
  wire  _T_2 = io_wr & io_rd; // @[FIFO.scala 34:25]
  wire [31:0] _T_7 = rPointer + 32'h1; // @[FIFO.scala 31:46]
  wire [31:0] _T_8 = rPointer == 32'h22 ? 32'h0 : _T_7; // @[FIFO.scala 31:10]
  wire [31:0] _T_12 = wPointer + 32'h1; // @[FIFO.scala 31:46]
  wire [31:0] _T_13 = wPointer == 32'h22 ? 32'h0 : _T_12; // @[FIFO.scala 31:10]
  wire  _GEN_4 = count == 32'h0 ? 1'h0 : 1'h1; // @[FIFO.scala 35:25 FIFO.scala 23:16 FIFO.scala 39:21]
  wire  _T_17 = count < 32'h23; // @[FIFO.scala 48:16]
  wire [31:0] _T_24 = count + 32'h1; // @[FIFO.scala 51:22]
  wire  _T_28 = count > 32'h0; // @[FIFO.scala 55:16]
  wire [31:0] _T_35 = count - 32'h1; // @[FIFO.scala 59:22]
  wire [31:0] _GEN_21 = count > 32'h0 ? $signed(mem_MPORT_3_data) : $signed(32'sh0); // @[FIFO.scala 55:23 FIFO.scala 56:15 FIFO.scala 61:15]
  wire [31:0] _GEN_22 = count > 32'h0 ? _T_8 : rPointer; // @[FIFO.scala 55:23 FIFO.scala 57:16 FIFO.scala 25:25]
  wire [31:0] _GEN_23 = count > 32'h0 ? _T_35 : count; // @[FIFO.scala 55:23 FIFO.scala 59:13 FIFO.scala 22:22]
  wire  _GEN_26 = ~io_wr & io_rd & _T_28; // @[FIFO.scala 54:55 FIFO.scala 23:16]
  wire  _GEN_31 = io_wr & ~io_rd ? 1'h0 : _GEN_26; // @[FIFO.scala 45:55]
  wire  _GEN_34 = io_wr & ~io_rd & _T_17; // @[FIFO.scala 45:55 FIFO.scala 23:16]
  assign mem_MPORT_addr = rPointer[5:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_data = mem[mem_MPORT_addr]; // @[FIFO.scala 23:16]
  `else
  assign mem_MPORT_data = mem_MPORT_addr >= 6'h23 ? _RAND_1[31:0] : mem[mem_MPORT_addr]; // @[FIFO.scala 23:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_3_addr = rPointer[5:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_3_data = mem[mem_MPORT_3_addr]; // @[FIFO.scala 23:16]
  `else
  assign mem_MPORT_3_data = mem_MPORT_3_addr >= 6'h23 ? _RAND_2[31:0] : mem[mem_MPORT_3_addr]; // @[FIFO.scala 23:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_1_data = io_datain;
  assign mem_MPORT_1_addr = wPointer[5:0];
  assign mem_MPORT_1_mask = 1'h1;
  assign mem_MPORT_1_en = _T_2 & _GEN_4;
  assign mem_MPORT_2_data = io_datain;
  assign mem_MPORT_2_addr = wPointer[5:0];
  assign mem_MPORT_2_mask = 1'h1;
  assign mem_MPORT_2_en = _T_2 ? 1'h0 : _GEN_34;
  assign io_dataout = dataout; // @[FIFO.scala 69:14]
  assign io_empty = count == 32'h0; // @[FIFO.scala 71:22]
  always @(posedge clock) begin
    if(mem_MPORT_1_en & mem_MPORT_1_mask) begin
      mem[mem_MPORT_1_addr] <= mem_MPORT_1_data; // @[FIFO.scala 23:16]
    end
    if(mem_MPORT_2_en & mem_MPORT_2_mask) begin
      mem[mem_MPORT_2_addr] <= mem_MPORT_2_data; // @[FIFO.scala 23:16]
    end
    if (reset) begin // @[FIFO.scala 22:22]
      count <= 32'h0; // @[FIFO.scala 22:22]
    end else if (!(io_wr & io_rd)) begin // @[FIFO.scala 34:46]
      if (io_wr & ~io_rd) begin // @[FIFO.scala 45:55]
        if (count < 32'h23) begin // @[FIFO.scala 48:26]
          count <= _T_24; // @[FIFO.scala 51:13]
        end
      end else if (~io_wr & io_rd) begin // @[FIFO.scala 54:55]
        count <= _GEN_23;
      end
    end
    if (reset) begin // @[FIFO.scala 24:25]
      wPointer <= 32'h0; // @[FIFO.scala 24:25]
    end else if (io_wr & io_rd) begin // @[FIFO.scala 34:46]
      if (!(count == 32'h0)) begin // @[FIFO.scala 35:25]
        wPointer <= _T_13; // @[FIFO.scala 43:16]
      end
    end else if (io_wr & ~io_rd) begin // @[FIFO.scala 45:55]
      if (count < 32'h23) begin // @[FIFO.scala 48:26]
        wPointer <= _T_13; // @[FIFO.scala 50:16]
      end
    end
    if (reset) begin // @[FIFO.scala 25:25]
      rPointer <= 32'h0; // @[FIFO.scala 25:25]
    end else if (io_wr & io_rd) begin // @[FIFO.scala 34:46]
      if (!(count == 32'h0)) begin // @[FIFO.scala 35:25]
        if (rPointer == 32'h22) begin // @[FIFO.scala 31:10]
          rPointer <= 32'h0;
        end else begin
          rPointer <= _T_7;
        end
      end
    end else if (!(io_wr & ~io_rd)) begin // @[FIFO.scala 45:55]
      if (~io_wr & io_rd) begin // @[FIFO.scala 54:55]
        rPointer <= _GEN_22;
      end
    end
    if (reset) begin // @[FIFO.scala 26:24]
      dataout <= 32'sh0; // @[FIFO.scala 26:24]
    end else if (io_wr & io_rd) begin // @[FIFO.scala 34:46]
      if (count == 32'h0) begin // @[FIFO.scala 35:25]
        dataout <= io_datain; // @[FIFO.scala 36:17]
      end else begin
        dataout <= mem_MPORT_data; // @[FIFO.scala 39:15]
      end
    end else if (io_wr & ~io_rd) begin // @[FIFO.scala 45:55]
      dataout <= 32'sh0; // @[FIFO.scala 46:13]
    end else if (~io_wr & io_rd) begin // @[FIFO.scala 54:55]
      dataout <= _GEN_21;
    end else begin
      dataout <= 32'sh0; // @[FIFO.scala 65:13]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {1{`RANDOM}};
  _RAND_2 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 35; initvar = initvar+1)
    mem[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  count = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  wPointer = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  rPointer = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  dataout = _RAND_6[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FIFO_0(
  input         clock,
  input         reset,
  input  [31:0] io_datain,
  output [31:0] io_dataout,
  input         io_wr,
  input         io_rd,
  output        io_empty
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] mem [0:34]; // @[FIFO_0.scala 23:16]
  wire [31:0] mem_MPORT_data; // @[FIFO_0.scala 23:16]
  wire [5:0] mem_MPORT_addr; // @[FIFO_0.scala 23:16]
  wire [31:0] mem_MPORT_3_data; // @[FIFO_0.scala 23:16]
  wire [5:0] mem_MPORT_3_addr; // @[FIFO_0.scala 23:16]
  wire [31:0] mem_MPORT_1_data; // @[FIFO_0.scala 23:16]
  wire [5:0] mem_MPORT_1_addr; // @[FIFO_0.scala 23:16]
  wire  mem_MPORT_1_mask; // @[FIFO_0.scala 23:16]
  wire  mem_MPORT_1_en; // @[FIFO_0.scala 23:16]
  wire [31:0] mem_MPORT_2_data; // @[FIFO_0.scala 23:16]
  wire [5:0] mem_MPORT_2_addr; // @[FIFO_0.scala 23:16]
  wire  mem_MPORT_2_mask; // @[FIFO_0.scala 23:16]
  wire  mem_MPORT_2_en; // @[FIFO_0.scala 23:16]
  reg [31:0] count; // @[FIFO_0.scala 22:22]
  reg [31:0] wPointer; // @[FIFO_0.scala 24:25]
  reg [31:0] rPointer; // @[FIFO_0.scala 25:25]
  reg [31:0] dataout; // @[FIFO_0.scala 26:24]
  wire  _T_2 = io_wr & io_rd; // @[FIFO_0.scala 33:25]
  wire [31:0] _T_7 = rPointer + 32'h1; // @[FIFO_0.scala 30:46]
  wire [31:0] _T_8 = rPointer == 32'h22 ? 32'h0 : _T_7; // @[FIFO_0.scala 30:10]
  wire [31:0] _T_12 = wPointer + 32'h1; // @[FIFO_0.scala 30:46]
  wire [31:0] _T_13 = wPointer == 32'h22 ? 32'h0 : _T_12; // @[FIFO_0.scala 30:10]
  wire  _GEN_4 = count == 32'h0 ? 1'h0 : 1'h1; // @[FIFO_0.scala 34:25 FIFO_0.scala 23:16 FIFO_0.scala 38:21]
  wire  _T_17 = count < 32'h23; // @[FIFO_0.scala 47:16]
  wire [31:0] _T_24 = count + 32'h1; // @[FIFO_0.scala 50:22]
  wire  _T_28 = count > 32'h0; // @[FIFO_0.scala 54:16]
  wire [31:0] _T_35 = count - 32'h1; // @[FIFO_0.scala 58:22]
  wire [31:0] _GEN_21 = count > 32'h0 ? mem_MPORT_3_data : 32'h0; // @[FIFO_0.scala 54:23 FIFO_0.scala 55:15 FIFO_0.scala 60:15]
  wire [31:0] _GEN_22 = count > 32'h0 ? _T_8 : rPointer; // @[FIFO_0.scala 54:23 FIFO_0.scala 56:16 FIFO_0.scala 25:25]
  wire [31:0] _GEN_23 = count > 32'h0 ? _T_35 : count; // @[FIFO_0.scala 54:23 FIFO_0.scala 58:13 FIFO_0.scala 22:22]
  wire  _GEN_26 = ~io_wr & io_rd & _T_28; // @[FIFO_0.scala 53:55 FIFO_0.scala 23:16]
  wire  _GEN_31 = io_wr & ~io_rd ? 1'h0 : _GEN_26; // @[FIFO_0.scala 44:55]
  wire  _GEN_34 = io_wr & ~io_rd & _T_17; // @[FIFO_0.scala 44:55 FIFO_0.scala 23:16]
  assign mem_MPORT_addr = rPointer[5:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_data = mem[mem_MPORT_addr]; // @[FIFO_0.scala 23:16]
  `else
  assign mem_MPORT_data = mem_MPORT_addr >= 6'h23 ? _RAND_1[31:0] : mem[mem_MPORT_addr]; // @[FIFO_0.scala 23:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_3_addr = rPointer[5:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_3_data = mem[mem_MPORT_3_addr]; // @[FIFO_0.scala 23:16]
  `else
  assign mem_MPORT_3_data = mem_MPORT_3_addr >= 6'h23 ? _RAND_2[31:0] : mem[mem_MPORT_3_addr]; // @[FIFO_0.scala 23:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_1_data = io_datain;
  assign mem_MPORT_1_addr = wPointer[5:0];
  assign mem_MPORT_1_mask = 1'h1;
  assign mem_MPORT_1_en = _T_2 & _GEN_4;
  assign mem_MPORT_2_data = io_datain;
  assign mem_MPORT_2_addr = wPointer[5:0];
  assign mem_MPORT_2_mask = 1'h1;
  assign mem_MPORT_2_en = _T_2 ? 1'h0 : _GEN_34;
  assign io_dataout = dataout; // @[FIFO_0.scala 68:14]
  assign io_empty = count == 32'h0; // @[FIFO_0.scala 70:22]
  always @(posedge clock) begin
    if(mem_MPORT_1_en & mem_MPORT_1_mask) begin
      mem[mem_MPORT_1_addr] <= mem_MPORT_1_data; // @[FIFO_0.scala 23:16]
    end
    if(mem_MPORT_2_en & mem_MPORT_2_mask) begin
      mem[mem_MPORT_2_addr] <= mem_MPORT_2_data; // @[FIFO_0.scala 23:16]
    end
    if (reset) begin // @[FIFO_0.scala 22:22]
      count <= 32'h0; // @[FIFO_0.scala 22:22]
    end else if (!(io_wr & io_rd)) begin // @[FIFO_0.scala 33:46]
      if (io_wr & ~io_rd) begin // @[FIFO_0.scala 44:55]
        if (count < 32'h23) begin // @[FIFO_0.scala 47:26]
          count <= _T_24; // @[FIFO_0.scala 50:13]
        end
      end else if (~io_wr & io_rd) begin // @[FIFO_0.scala 53:55]
        count <= _GEN_23;
      end
    end
    if (reset) begin // @[FIFO_0.scala 24:25]
      wPointer <= 32'h0; // @[FIFO_0.scala 24:25]
    end else if (io_wr & io_rd) begin // @[FIFO_0.scala 33:46]
      if (!(count == 32'h0)) begin // @[FIFO_0.scala 34:25]
        wPointer <= _T_13; // @[FIFO_0.scala 42:16]
      end
    end else if (io_wr & ~io_rd) begin // @[FIFO_0.scala 44:55]
      if (count < 32'h23) begin // @[FIFO_0.scala 47:26]
        wPointer <= _T_13; // @[FIFO_0.scala 49:16]
      end
    end
    if (reset) begin // @[FIFO_0.scala 25:25]
      rPointer <= 32'h0; // @[FIFO_0.scala 25:25]
    end else if (io_wr & io_rd) begin // @[FIFO_0.scala 33:46]
      if (!(count == 32'h0)) begin // @[FIFO_0.scala 34:25]
        if (rPointer == 32'h22) begin // @[FIFO_0.scala 30:10]
          rPointer <= 32'h0;
        end else begin
          rPointer <= _T_7;
        end
      end
    end else if (!(io_wr & ~io_rd)) begin // @[FIFO_0.scala 44:55]
      if (~io_wr & io_rd) begin // @[FIFO_0.scala 53:55]
        rPointer <= _GEN_22;
      end
    end
    if (reset) begin // @[FIFO_0.scala 26:24]
      dataout <= 32'h0; // @[FIFO_0.scala 26:24]
    end else if (io_wr & io_rd) begin // @[FIFO_0.scala 33:46]
      if (count == 32'h0) begin // @[FIFO_0.scala 34:25]
        dataout <= io_datain; // @[FIFO_0.scala 35:17]
      end else begin
        dataout <= mem_MPORT_data; // @[FIFO_0.scala 38:15]
      end
    end else if (io_wr & ~io_rd) begin // @[FIFO_0.scala 44:55]
      dataout <= 32'h0; // @[FIFO_0.scala 45:13]
    end else if (~io_wr & io_rd) begin // @[FIFO_0.scala 53:55]
      dataout <= _GEN_21;
    end else begin
      dataout <= 32'h0; // @[FIFO_0.scala 64:13]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {1{`RANDOM}};
  _RAND_2 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 35; initvar = initvar+1)
    mem[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  count = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  wPointer = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  rPointer = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  dataout = _RAND_6[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbitration_1(
  input         clock,
  input         reset,
  input  [31:0] io_node_id_0,
  input  [63:0] io_ray_id_0,
  input  [31:0] io_hit_0,
  input         io_valid_0,
  input  [31:0] io_node_id_1,
  input  [31:0] io_ray_id_1,
  input         io_valid_1,
  input  [31:0] io_ray_id_2,
  input         io_valid_2,
  output [31:0] io_node_id_out,
  output [31:0] io_ray_id_out,
  output [31:0] io_hit_out,
  output        io_valid_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  FIFO_A_1_0_node_clock; // @[Arbitration_1_1.scala 29:38]
  wire  FIFO_A_1_0_node_reset; // @[Arbitration_1_1.scala 29:38]
  wire [31:0] FIFO_A_1_0_node_io_datain; // @[Arbitration_1_1.scala 29:38]
  wire [31:0] FIFO_A_1_0_node_io_dataout; // @[Arbitration_1_1.scala 29:38]
  wire  FIFO_A_1_0_node_io_wr; // @[Arbitration_1_1.scala 29:38]
  wire  FIFO_A_1_0_node_io_rd; // @[Arbitration_1_1.scala 29:38]
  wire  FIFO_A_1_0_node_io_empty; // @[Arbitration_1_1.scala 29:38]
  wire  FIFO_A_1_0_ray_clock; // @[Arbitration_1_1.scala 30:41]
  wire  FIFO_A_1_0_ray_reset; // @[Arbitration_1_1.scala 30:41]
  wire [31:0] FIFO_A_1_0_ray_io_datain; // @[Arbitration_1_1.scala 30:41]
  wire [31:0] FIFO_A_1_0_ray_io_dataout; // @[Arbitration_1_1.scala 30:41]
  wire  FIFO_A_1_0_ray_io_wr; // @[Arbitration_1_1.scala 30:41]
  wire  FIFO_A_1_0_ray_io_rd; // @[Arbitration_1_1.scala 30:41]
  wire  FIFO_A_1_0_ray_io_empty; // @[Arbitration_1_1.scala 30:41]
  wire  FIFO_A_1_0_hit_clock; // @[Arbitration_1_1.scala 31:42]
  wire  FIFO_A_1_0_hit_reset; // @[Arbitration_1_1.scala 31:42]
  wire [31:0] FIFO_A_1_0_hit_io_datain; // @[Arbitration_1_1.scala 31:42]
  wire [31:0] FIFO_A_1_0_hit_io_dataout; // @[Arbitration_1_1.scala 31:42]
  wire  FIFO_A_1_0_hit_io_wr; // @[Arbitration_1_1.scala 31:42]
  wire  FIFO_A_1_0_hit_io_rd; // @[Arbitration_1_1.scala 31:42]
  wire  FIFO_A_1_0_hit_io_empty; // @[Arbitration_1_1.scala 31:42]
  wire  FIFO_A_1_1_node_clock; // @[Arbitration_1_1.scala 33:38]
  wire  FIFO_A_1_1_node_reset; // @[Arbitration_1_1.scala 33:38]
  wire [31:0] FIFO_A_1_1_node_io_datain; // @[Arbitration_1_1.scala 33:38]
  wire [31:0] FIFO_A_1_1_node_io_dataout; // @[Arbitration_1_1.scala 33:38]
  wire  FIFO_A_1_1_node_io_wr; // @[Arbitration_1_1.scala 33:38]
  wire  FIFO_A_1_1_node_io_rd; // @[Arbitration_1_1.scala 33:38]
  wire  FIFO_A_1_1_node_io_empty; // @[Arbitration_1_1.scala 33:38]
  wire  FIFO_A_1_1_ray_clock; // @[Arbitration_1_1.scala 34:41]
  wire  FIFO_A_1_1_ray_reset; // @[Arbitration_1_1.scala 34:41]
  wire [31:0] FIFO_A_1_1_ray_io_datain; // @[Arbitration_1_1.scala 34:41]
  wire [31:0] FIFO_A_1_1_ray_io_dataout; // @[Arbitration_1_1.scala 34:41]
  wire  FIFO_A_1_1_ray_io_wr; // @[Arbitration_1_1.scala 34:41]
  wire  FIFO_A_1_1_ray_io_rd; // @[Arbitration_1_1.scala 34:41]
  wire  FIFO_A_1_1_ray_io_empty; // @[Arbitration_1_1.scala 34:41]
  wire  FIFO_A_1_2_node_clock; // @[Arbitration_1_1.scala 36:38]
  wire  FIFO_A_1_2_node_reset; // @[Arbitration_1_1.scala 36:38]
  wire [31:0] FIFO_A_1_2_node_io_datain; // @[Arbitration_1_1.scala 36:38]
  wire [31:0] FIFO_A_1_2_node_io_dataout; // @[Arbitration_1_1.scala 36:38]
  wire  FIFO_A_1_2_node_io_wr; // @[Arbitration_1_1.scala 36:38]
  wire  FIFO_A_1_2_node_io_rd; // @[Arbitration_1_1.scala 36:38]
  wire  FIFO_A_1_2_node_io_empty; // @[Arbitration_1_1.scala 36:38]
  wire  FIFO_A_1_2_ray_clock; // @[Arbitration_1_1.scala 37:41]
  wire  FIFO_A_1_2_ray_reset; // @[Arbitration_1_1.scala 37:41]
  wire [31:0] FIFO_A_1_2_ray_io_datain; // @[Arbitration_1_1.scala 37:41]
  wire [31:0] FIFO_A_1_2_ray_io_dataout; // @[Arbitration_1_1.scala 37:41]
  wire  FIFO_A_1_2_ray_io_wr; // @[Arbitration_1_1.scala 37:41]
  wire  FIFO_A_1_2_ray_io_rd; // @[Arbitration_1_1.scala 37:41]
  wire  FIFO_A_1_2_ray_io_empty; // @[Arbitration_1_1.scala 37:41]
  reg  valid_out_temp; // @[Arbitration_1_1.scala 63:59]
  wire  _T_1 = FIFO_A_1_0_node_io_empty; // @[Arbitration_1_1.scala 78:45]
  wire  _T_3 = FIFO_A_1_0_node_io_empty & ~FIFO_A_1_1_node_io_empty; // @[Arbitration_1_1.scala 78:53]
  wire  _T_8 = _T_1 & FIFO_A_1_1_node_io_empty & ~FIFO_A_1_2_node_io_empty; // @[Arbitration_1_1.scala 91:88]
  wire  _GEN_4 = FIFO_A_1_0_node_io_empty & ~FIFO_A_1_1_node_io_empty ? 1'h0 : _T_8; // @[Arbitration_1_1.scala 78:89 Arbitration_1_1.scala 84:44]
  reg  FIFO_0_empty; // @[Arbitration_1_1.scala 116:58]
  reg  FIFO_1_empty; // @[Arbitration_1_1.scala 117:58]
  reg  FIFO_2_empty; // @[Arbitration_1_1.scala 118:58]
  wire [31:0] _GEN_8 = FIFO_0_empty & FIFO_1_empty & ~FIFO_2_empty ? $signed(FIFO_A_1_2_node_io_dataout) : $signed(32'sh0
    ); // @[Arbitration_1_1.scala 157:85 Arbitration_1_1.scala 158:45 Arbitration_1_1.scala 165:45]
  wire [31:0] _GEN_9 = FIFO_0_empty & FIFO_1_empty & ~FIFO_2_empty ? FIFO_A_1_2_ray_io_dataout : 32'h0; // @[Arbitration_1_1.scala 157:85 Arbitration_1_1.scala 159:48 Arbitration_1_1.scala 166:48]
  wire  _GEN_11 = FIFO_0_empty & FIFO_1_empty & ~FIFO_2_empty & valid_out_temp; // @[Arbitration_1_1.scala 157:85 Arbitration_1_1.scala 162:50 Arbitration_1_1.scala 168:50]
  wire [31:0] _GEN_12 = FIFO_0_empty & ~FIFO_1_empty ? $signed(FIFO_A_1_1_node_io_dataout) : $signed(_GEN_8); // @[Arbitration_1_1.scala 151:63 Arbitration_1_1.scala 152:46]
  wire [31:0] _GEN_13 = FIFO_0_empty & ~FIFO_1_empty ? FIFO_A_1_1_ray_io_dataout : _GEN_9; // @[Arbitration_1_1.scala 151:63 Arbitration_1_1.scala 153:49]
  wire  _GEN_15 = FIFO_0_empty & ~FIFO_1_empty ? valid_out_temp : _GEN_11; // @[Arbitration_1_1.scala 151:63 Arbitration_1_1.scala 155:50]
  FIFO FIFO_A_1_0_node ( // @[Arbitration_1_1.scala 29:38]
    .clock(FIFO_A_1_0_node_clock),
    .reset(FIFO_A_1_0_node_reset),
    .io_datain(FIFO_A_1_0_node_io_datain),
    .io_dataout(FIFO_A_1_0_node_io_dataout),
    .io_wr(FIFO_A_1_0_node_io_wr),
    .io_rd(FIFO_A_1_0_node_io_rd),
    .io_empty(FIFO_A_1_0_node_io_empty)
  );
  FIFO_0 FIFO_A_1_0_ray ( // @[Arbitration_1_1.scala 30:41]
    .clock(FIFO_A_1_0_ray_clock),
    .reset(FIFO_A_1_0_ray_reset),
    .io_datain(FIFO_A_1_0_ray_io_datain),
    .io_dataout(FIFO_A_1_0_ray_io_dataout),
    .io_wr(FIFO_A_1_0_ray_io_wr),
    .io_rd(FIFO_A_1_0_ray_io_rd),
    .io_empty(FIFO_A_1_0_ray_io_empty)
  );
  FIFO_0 FIFO_A_1_0_hit ( // @[Arbitration_1_1.scala 31:42]
    .clock(FIFO_A_1_0_hit_clock),
    .reset(FIFO_A_1_0_hit_reset),
    .io_datain(FIFO_A_1_0_hit_io_datain),
    .io_dataout(FIFO_A_1_0_hit_io_dataout),
    .io_wr(FIFO_A_1_0_hit_io_wr),
    .io_rd(FIFO_A_1_0_hit_io_rd),
    .io_empty(FIFO_A_1_0_hit_io_empty)
  );
  FIFO FIFO_A_1_1_node ( // @[Arbitration_1_1.scala 33:38]
    .clock(FIFO_A_1_1_node_clock),
    .reset(FIFO_A_1_1_node_reset),
    .io_datain(FIFO_A_1_1_node_io_datain),
    .io_dataout(FIFO_A_1_1_node_io_dataout),
    .io_wr(FIFO_A_1_1_node_io_wr),
    .io_rd(FIFO_A_1_1_node_io_rd),
    .io_empty(FIFO_A_1_1_node_io_empty)
  );
  FIFO_0 FIFO_A_1_1_ray ( // @[Arbitration_1_1.scala 34:41]
    .clock(FIFO_A_1_1_ray_clock),
    .reset(FIFO_A_1_1_ray_reset),
    .io_datain(FIFO_A_1_1_ray_io_datain),
    .io_dataout(FIFO_A_1_1_ray_io_dataout),
    .io_wr(FIFO_A_1_1_ray_io_wr),
    .io_rd(FIFO_A_1_1_ray_io_rd),
    .io_empty(FIFO_A_1_1_ray_io_empty)
  );
  FIFO FIFO_A_1_2_node ( // @[Arbitration_1_1.scala 36:38]
    .clock(FIFO_A_1_2_node_clock),
    .reset(FIFO_A_1_2_node_reset),
    .io_datain(FIFO_A_1_2_node_io_datain),
    .io_dataout(FIFO_A_1_2_node_io_dataout),
    .io_wr(FIFO_A_1_2_node_io_wr),
    .io_rd(FIFO_A_1_2_node_io_rd),
    .io_empty(FIFO_A_1_2_node_io_empty)
  );
  FIFO_0 FIFO_A_1_2_ray ( // @[Arbitration_1_1.scala 37:41]
    .clock(FIFO_A_1_2_ray_clock),
    .reset(FIFO_A_1_2_ray_reset),
    .io_datain(FIFO_A_1_2_ray_io_datain),
    .io_dataout(FIFO_A_1_2_ray_io_dataout),
    .io_wr(FIFO_A_1_2_ray_io_wr),
    .io_rd(FIFO_A_1_2_ray_io_rd),
    .io_empty(FIFO_A_1_2_ray_io_empty)
  );
  assign io_node_id_out = ~FIFO_0_empty ? $signed(FIFO_A_1_0_node_io_dataout) : $signed(_GEN_12); // @[Arbitration_1_1.scala 143:35 Arbitration_1_1.scala 144:45]
  assign io_ray_id_out = ~FIFO_0_empty ? FIFO_A_1_0_ray_io_dataout : _GEN_13; // @[Arbitration_1_1.scala 143:35 Arbitration_1_1.scala 145:46]
  assign io_hit_out = ~FIFO_0_empty ? FIFO_A_1_0_hit_io_dataout : 32'h0; // @[Arbitration_1_1.scala 143:35 Arbitration_1_1.scala 147:52]
  assign io_valid_out = ~FIFO_0_empty ? valid_out_temp : _GEN_15; // @[Arbitration_1_1.scala 143:35 Arbitration_1_1.scala 150:50]
  assign FIFO_A_1_0_node_clock = clock;
  assign FIFO_A_1_0_node_reset = reset;
  assign FIFO_A_1_0_node_io_datain = io_node_id_0; // @[Arbitration_1_1.scala 42:40]
  assign FIFO_A_1_0_node_io_wr = io_valid_0; // @[Arbitration_1_1.scala 39:44]
  assign FIFO_A_1_0_node_io_rd = ~FIFO_A_1_0_node_io_empty; // @[Arbitration_1_1.scala 65:39]
  assign FIFO_A_1_0_ray_clock = clock;
  assign FIFO_A_1_0_ray_reset = reset;
  assign FIFO_A_1_0_ray_io_datain = io_ray_id_0[31:0]; // @[Arbitration_1_1.scala 43:43]
  assign FIFO_A_1_0_ray_io_wr = io_valid_0; // @[Arbitration_1_1.scala 40:47]
  assign FIFO_A_1_0_ray_io_rd = ~FIFO_A_1_0_node_io_empty; // @[Arbitration_1_1.scala 65:39]
  assign FIFO_A_1_0_hit_clock = clock;
  assign FIFO_A_1_0_hit_reset = reset;
  assign FIFO_A_1_0_hit_io_datain = io_hit_0; // @[Arbitration_1_1.scala 44:44]
  assign FIFO_A_1_0_hit_io_wr = io_valid_0; // @[Arbitration_1_1.scala 41:48]
  assign FIFO_A_1_0_hit_io_rd = ~FIFO_A_1_0_node_io_empty; // @[Arbitration_1_1.scala 65:39]
  assign FIFO_A_1_1_node_clock = clock;
  assign FIFO_A_1_1_node_reset = reset;
  assign FIFO_A_1_1_node_io_datain = io_node_id_1; // @[Arbitration_1_1.scala 48:40]
  assign FIFO_A_1_1_node_io_wr = io_valid_1; // @[Arbitration_1_1.scala 46:44]
  assign FIFO_A_1_1_node_io_rd = ~FIFO_A_1_0_node_io_empty ? 1'h0 : _T_3; // @[Arbitration_1_1.scala 65:47 Arbitration_1_1.scala 69:44]
  assign FIFO_A_1_1_ray_clock = clock;
  assign FIFO_A_1_1_ray_reset = reset;
  assign FIFO_A_1_1_ray_io_datain = io_ray_id_1; // @[Arbitration_1_1.scala 49:43]
  assign FIFO_A_1_1_ray_io_wr = io_valid_1; // @[Arbitration_1_1.scala 47:47]
  assign FIFO_A_1_1_ray_io_rd = ~FIFO_A_1_0_node_io_empty ? 1'h0 : _T_3; // @[Arbitration_1_1.scala 65:47 Arbitration_1_1.scala 69:44]
  assign FIFO_A_1_2_node_clock = clock;
  assign FIFO_A_1_2_node_reset = reset;
  assign FIFO_A_1_2_node_io_datain = 32'sh0; // @[Arbitration_1_1.scala 53:40]
  assign FIFO_A_1_2_node_io_wr = io_valid_2; // @[Arbitration_1_1.scala 51:44]
  assign FIFO_A_1_2_node_io_rd = ~FIFO_A_1_0_node_io_empty ? 1'h0 : _GEN_4; // @[Arbitration_1_1.scala 65:47 Arbitration_1_1.scala 71:44]
  assign FIFO_A_1_2_ray_clock = clock;
  assign FIFO_A_1_2_ray_reset = reset;
  assign FIFO_A_1_2_ray_io_datain = io_ray_id_2; // @[Arbitration_1_1.scala 54:43]
  assign FIFO_A_1_2_ray_io_wr = io_valid_2; // @[Arbitration_1_1.scala 52:47]
  assign FIFO_A_1_2_ray_io_rd = ~FIFO_A_1_0_node_io_empty ? 1'h0 : _GEN_4; // @[Arbitration_1_1.scala 65:47 Arbitration_1_1.scala 71:44]
  always @(posedge clock) begin
    if (reset) begin // @[Arbitration_1_1.scala 63:59]
      valid_out_temp <= 1'h0; // @[Arbitration_1_1.scala 63:59]
    end else begin
      valid_out_temp <= FIFO_A_1_0_node_io_rd | FIFO_A_1_1_node_io_rd | FIFO_A_1_2_node_io_rd; // @[Arbitration_1_1.scala 139:51]
    end
    if (reset) begin // @[Arbitration_1_1.scala 116:58]
      FIFO_0_empty <= 1'h0; // @[Arbitration_1_1.scala 116:58]
    end else begin
      FIFO_0_empty <= FIFO_A_1_0_node_io_empty; // @[Arbitration_1_1.scala 120:52]
    end
    if (reset) begin // @[Arbitration_1_1.scala 117:58]
      FIFO_1_empty <= 1'h0; // @[Arbitration_1_1.scala 117:58]
    end else begin
      FIFO_1_empty <= FIFO_A_1_1_node_io_empty; // @[Arbitration_1_1.scala 121:52]
    end
    if (reset) begin // @[Arbitration_1_1.scala 118:58]
      FIFO_2_empty <= 1'h0; // @[Arbitration_1_1.scala 118:58]
    end else begin
      FIFO_2_empty <= FIFO_A_1_2_node_io_empty; // @[Arbitration_1_1.scala 122:52]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid_out_temp = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  FIFO_0_empty = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  FIFO_1_empty = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  FIFO_2_empty = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbitration_2_1(
  input         clock,
  input         reset,
  input  [31:0] io_ray_id_2_0,
  input  [31:0] io_hit_2_0,
  input         io_valid_2_0,
  input  [31:0] io_ray_id_2_1,
  input  [31:0] io_hit_2_1,
  input         io_valid_2_1,
  input  [31:0] io_ray_id_2_2,
  input  [31:0] io_hit_2_2,
  input         io_valid_2_2,
  input  [31:0] io_ray_id_2_3,
  input  [31:0] io_hit_2_3,
  input         io_valid_2_3,
  output [31:0] io_ray_id_out,
  output [31:0] io_hit_out,
  output        io_valid_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  FIFO_A_2_0_ray_clock; // @[Arbitration_2_1.scala 38:41]
  wire  FIFO_A_2_0_ray_reset; // @[Arbitration_2_1.scala 38:41]
  wire [31:0] FIFO_A_2_0_ray_io_datain; // @[Arbitration_2_1.scala 38:41]
  wire [31:0] FIFO_A_2_0_ray_io_dataout; // @[Arbitration_2_1.scala 38:41]
  wire  FIFO_A_2_0_ray_io_wr; // @[Arbitration_2_1.scala 38:41]
  wire  FIFO_A_2_0_ray_io_rd; // @[Arbitration_2_1.scala 38:41]
  wire  FIFO_A_2_0_ray_io_empty; // @[Arbitration_2_1.scala 38:41]
  wire  FIFO_A_2_0_hit_clock; // @[Arbitration_2_1.scala 39:42]
  wire  FIFO_A_2_0_hit_reset; // @[Arbitration_2_1.scala 39:42]
  wire [31:0] FIFO_A_2_0_hit_io_datain; // @[Arbitration_2_1.scala 39:42]
  wire [31:0] FIFO_A_2_0_hit_io_dataout; // @[Arbitration_2_1.scala 39:42]
  wire  FIFO_A_2_0_hit_io_wr; // @[Arbitration_2_1.scala 39:42]
  wire  FIFO_A_2_0_hit_io_rd; // @[Arbitration_2_1.scala 39:42]
  wire  FIFO_A_2_0_hit_io_empty; // @[Arbitration_2_1.scala 39:42]
  wire  FIFO_A_2_1_ray_clock; // @[Arbitration_2_1.scala 41:41]
  wire  FIFO_A_2_1_ray_reset; // @[Arbitration_2_1.scala 41:41]
  wire [31:0] FIFO_A_2_1_ray_io_datain; // @[Arbitration_2_1.scala 41:41]
  wire [31:0] FIFO_A_2_1_ray_io_dataout; // @[Arbitration_2_1.scala 41:41]
  wire  FIFO_A_2_1_ray_io_wr; // @[Arbitration_2_1.scala 41:41]
  wire  FIFO_A_2_1_ray_io_rd; // @[Arbitration_2_1.scala 41:41]
  wire  FIFO_A_2_1_ray_io_empty; // @[Arbitration_2_1.scala 41:41]
  wire  FIFO_A_2_1_hit_clock; // @[Arbitration_2_1.scala 42:42]
  wire  FIFO_A_2_1_hit_reset; // @[Arbitration_2_1.scala 42:42]
  wire [31:0] FIFO_A_2_1_hit_io_datain; // @[Arbitration_2_1.scala 42:42]
  wire [31:0] FIFO_A_2_1_hit_io_dataout; // @[Arbitration_2_1.scala 42:42]
  wire  FIFO_A_2_1_hit_io_wr; // @[Arbitration_2_1.scala 42:42]
  wire  FIFO_A_2_1_hit_io_rd; // @[Arbitration_2_1.scala 42:42]
  wire  FIFO_A_2_1_hit_io_empty; // @[Arbitration_2_1.scala 42:42]
  wire  FIFO_A_2_2_ray_clock; // @[Arbitration_2_1.scala 44:41]
  wire  FIFO_A_2_2_ray_reset; // @[Arbitration_2_1.scala 44:41]
  wire [31:0] FIFO_A_2_2_ray_io_datain; // @[Arbitration_2_1.scala 44:41]
  wire [31:0] FIFO_A_2_2_ray_io_dataout; // @[Arbitration_2_1.scala 44:41]
  wire  FIFO_A_2_2_ray_io_wr; // @[Arbitration_2_1.scala 44:41]
  wire  FIFO_A_2_2_ray_io_rd; // @[Arbitration_2_1.scala 44:41]
  wire  FIFO_A_2_2_ray_io_empty; // @[Arbitration_2_1.scala 44:41]
  wire  FIFO_A_2_2_hit_clock; // @[Arbitration_2_1.scala 45:42]
  wire  FIFO_A_2_2_hit_reset; // @[Arbitration_2_1.scala 45:42]
  wire [31:0] FIFO_A_2_2_hit_io_datain; // @[Arbitration_2_1.scala 45:42]
  wire [31:0] FIFO_A_2_2_hit_io_dataout; // @[Arbitration_2_1.scala 45:42]
  wire  FIFO_A_2_2_hit_io_wr; // @[Arbitration_2_1.scala 45:42]
  wire  FIFO_A_2_2_hit_io_rd; // @[Arbitration_2_1.scala 45:42]
  wire  FIFO_A_2_2_hit_io_empty; // @[Arbitration_2_1.scala 45:42]
  wire  FIFO_A_2_3_ray_clock; // @[Arbitration_2_1.scala 47:41]
  wire  FIFO_A_2_3_ray_reset; // @[Arbitration_2_1.scala 47:41]
  wire [31:0] FIFO_A_2_3_ray_io_datain; // @[Arbitration_2_1.scala 47:41]
  wire [31:0] FIFO_A_2_3_ray_io_dataout; // @[Arbitration_2_1.scala 47:41]
  wire  FIFO_A_2_3_ray_io_wr; // @[Arbitration_2_1.scala 47:41]
  wire  FIFO_A_2_3_ray_io_rd; // @[Arbitration_2_1.scala 47:41]
  wire  FIFO_A_2_3_ray_io_empty; // @[Arbitration_2_1.scala 47:41]
  wire  FIFO_A_2_3_hit_clock; // @[Arbitration_2_1.scala 48:42]
  wire  FIFO_A_2_3_hit_reset; // @[Arbitration_2_1.scala 48:42]
  wire [31:0] FIFO_A_2_3_hit_io_datain; // @[Arbitration_2_1.scala 48:42]
  wire [31:0] FIFO_A_2_3_hit_io_dataout; // @[Arbitration_2_1.scala 48:42]
  wire  FIFO_A_2_3_hit_io_wr; // @[Arbitration_2_1.scala 48:42]
  wire  FIFO_A_2_3_hit_io_rd; // @[Arbitration_2_1.scala 48:42]
  wire  FIFO_A_2_3_hit_io_empty; // @[Arbitration_2_1.scala 48:42]
  reg  valid_out_temp; // @[Arbitration_2_1.scala 73:59]
  wire  _T_1 = FIFO_A_2_0_ray_io_empty; // @[Arbitration_2_1.scala 84:44]
  wire  _T_3 = FIFO_A_2_0_ray_io_empty & ~FIFO_A_2_1_ray_io_empty; // @[Arbitration_2_1.scala 84:52]
  wire  _T_6 = _T_1 & FIFO_A_2_1_ray_io_empty; // @[Arbitration_2_1.scala 93:52]
  wire  _T_8 = _T_1 & FIFO_A_2_1_ray_io_empty & ~FIFO_A_2_2_ray_io_empty; // @[Arbitration_2_1.scala 93:86]
  wire  _T_15 = _T_6 & FIFO_A_2_2_ray_io_empty & ~FIFO_A_2_3_ray_io_empty; // @[Arbitration_2_1.scala 102:119]
  wire  _GEN_4 = _T_1 & FIFO_A_2_1_ray_io_empty & ~FIFO_A_2_2_ray_io_empty ? 1'h0 : _T_15; // @[Arbitration_2_1.scala 93:120 Arbitration_2_1.scala 100:47]
  wire  _GEN_7 = FIFO_A_2_0_ray_io_empty & ~FIFO_A_2_1_ray_io_empty ? 1'h0 : _T_8; // @[Arbitration_2_1.scala 84:87 Arbitration_2_1.scala 89:47]
  wire  _GEN_8 = FIFO_A_2_0_ray_io_empty & ~FIFO_A_2_1_ray_io_empty ? 1'h0 : _GEN_4; // @[Arbitration_2_1.scala 84:87 Arbitration_2_1.scala 91:47]
  reg  FIFO_0_empty; // @[Arbitration_2_1.scala 121:58]
  reg  FIFO_1_empty; // @[Arbitration_2_1.scala 122:58]
  reg  FIFO_2_empty; // @[Arbitration_2_1.scala 123:58]
  reg  FIFO_3_empty; // @[Arbitration_2_1.scala 124:58]
  wire  _T_26 = FIFO_0_empty & FIFO_1_empty; // @[Arbitration_2_1.scala 158:40]
  wire [31:0] _GEN_13 = _T_26 & FIFO_2_empty & ~FIFO_3_empty ? FIFO_A_2_3_ray_io_dataout : 32'h0; // @[Arbitration_2_1.scala 162:107 Arbitration_2_1.scala 166:56 Arbitration_2_1.scala 173:60]
  wire [31:0] _GEN_14 = _T_26 & FIFO_2_empty & ~FIFO_3_empty ? FIFO_A_2_3_hit_io_dataout : 32'h0; // @[Arbitration_2_1.scala 162:107 Arbitration_2_1.scala 167:61 Arbitration_2_1.scala 174:64]
  wire  _GEN_15 = _T_26 & FIFO_2_empty & ~FIFO_3_empty & valid_out_temp; // @[Arbitration_2_1.scala 162:107 Arbitration_2_1.scala 168:59 Arbitration_2_1.scala 175:62]
  wire [31:0] _GEN_16 = FIFO_0_empty & FIFO_1_empty & ~FIFO_2_empty ? FIFO_A_2_2_ray_io_dataout : _GEN_13; // @[Arbitration_2_1.scala 158:85 Arbitration_2_1.scala 159:56]
  wire [31:0] _GEN_17 = FIFO_0_empty & FIFO_1_empty & ~FIFO_2_empty ? FIFO_A_2_2_hit_io_dataout : _GEN_14; // @[Arbitration_2_1.scala 158:85 Arbitration_2_1.scala 160:61]
  wire  _GEN_18 = FIFO_0_empty & FIFO_1_empty & ~FIFO_2_empty ? valid_out_temp : _GEN_15; // @[Arbitration_2_1.scala 158:85 Arbitration_2_1.scala 161:59]
  wire [31:0] _GEN_19 = FIFO_0_empty & ~FIFO_1_empty ? FIFO_A_2_1_ray_io_dataout : _GEN_16; // @[Arbitration_2_1.scala 154:63 Arbitration_2_1.scala 155:56]
  wire [31:0] _GEN_20 = FIFO_0_empty & ~FIFO_1_empty ? FIFO_A_2_1_hit_io_dataout : _GEN_17; // @[Arbitration_2_1.scala 154:63 Arbitration_2_1.scala 156:61]
  wire  _GEN_21 = FIFO_0_empty & ~FIFO_1_empty ? valid_out_temp : _GEN_18; // @[Arbitration_2_1.scala 154:63 Arbitration_2_1.scala 157:59]
  FIFO_0 FIFO_A_2_0_ray ( // @[Arbitration_2_1.scala 38:41]
    .clock(FIFO_A_2_0_ray_clock),
    .reset(FIFO_A_2_0_ray_reset),
    .io_datain(FIFO_A_2_0_ray_io_datain),
    .io_dataout(FIFO_A_2_0_ray_io_dataout),
    .io_wr(FIFO_A_2_0_ray_io_wr),
    .io_rd(FIFO_A_2_0_ray_io_rd),
    .io_empty(FIFO_A_2_0_ray_io_empty)
  );
  FIFO_0 FIFO_A_2_0_hit ( // @[Arbitration_2_1.scala 39:42]
    .clock(FIFO_A_2_0_hit_clock),
    .reset(FIFO_A_2_0_hit_reset),
    .io_datain(FIFO_A_2_0_hit_io_datain),
    .io_dataout(FIFO_A_2_0_hit_io_dataout),
    .io_wr(FIFO_A_2_0_hit_io_wr),
    .io_rd(FIFO_A_2_0_hit_io_rd),
    .io_empty(FIFO_A_2_0_hit_io_empty)
  );
  FIFO_0 FIFO_A_2_1_ray ( // @[Arbitration_2_1.scala 41:41]
    .clock(FIFO_A_2_1_ray_clock),
    .reset(FIFO_A_2_1_ray_reset),
    .io_datain(FIFO_A_2_1_ray_io_datain),
    .io_dataout(FIFO_A_2_1_ray_io_dataout),
    .io_wr(FIFO_A_2_1_ray_io_wr),
    .io_rd(FIFO_A_2_1_ray_io_rd),
    .io_empty(FIFO_A_2_1_ray_io_empty)
  );
  FIFO_0 FIFO_A_2_1_hit ( // @[Arbitration_2_1.scala 42:42]
    .clock(FIFO_A_2_1_hit_clock),
    .reset(FIFO_A_2_1_hit_reset),
    .io_datain(FIFO_A_2_1_hit_io_datain),
    .io_dataout(FIFO_A_2_1_hit_io_dataout),
    .io_wr(FIFO_A_2_1_hit_io_wr),
    .io_rd(FIFO_A_2_1_hit_io_rd),
    .io_empty(FIFO_A_2_1_hit_io_empty)
  );
  FIFO_0 FIFO_A_2_2_ray ( // @[Arbitration_2_1.scala 44:41]
    .clock(FIFO_A_2_2_ray_clock),
    .reset(FIFO_A_2_2_ray_reset),
    .io_datain(FIFO_A_2_2_ray_io_datain),
    .io_dataout(FIFO_A_2_2_ray_io_dataout),
    .io_wr(FIFO_A_2_2_ray_io_wr),
    .io_rd(FIFO_A_2_2_ray_io_rd),
    .io_empty(FIFO_A_2_2_ray_io_empty)
  );
  FIFO_0 FIFO_A_2_2_hit ( // @[Arbitration_2_1.scala 45:42]
    .clock(FIFO_A_2_2_hit_clock),
    .reset(FIFO_A_2_2_hit_reset),
    .io_datain(FIFO_A_2_2_hit_io_datain),
    .io_dataout(FIFO_A_2_2_hit_io_dataout),
    .io_wr(FIFO_A_2_2_hit_io_wr),
    .io_rd(FIFO_A_2_2_hit_io_rd),
    .io_empty(FIFO_A_2_2_hit_io_empty)
  );
  FIFO_0 FIFO_A_2_3_ray ( // @[Arbitration_2_1.scala 47:41]
    .clock(FIFO_A_2_3_ray_clock),
    .reset(FIFO_A_2_3_ray_reset),
    .io_datain(FIFO_A_2_3_ray_io_datain),
    .io_dataout(FIFO_A_2_3_ray_io_dataout),
    .io_wr(FIFO_A_2_3_ray_io_wr),
    .io_rd(FIFO_A_2_3_ray_io_rd),
    .io_empty(FIFO_A_2_3_ray_io_empty)
  );
  FIFO_0 FIFO_A_2_3_hit ( // @[Arbitration_2_1.scala 48:42]
    .clock(FIFO_A_2_3_hit_clock),
    .reset(FIFO_A_2_3_hit_reset),
    .io_datain(FIFO_A_2_3_hit_io_datain),
    .io_dataout(FIFO_A_2_3_hit_io_dataout),
    .io_wr(FIFO_A_2_3_hit_io_wr),
    .io_rd(FIFO_A_2_3_hit_io_rd),
    .io_empty(FIFO_A_2_3_hit_io_empty)
  );
  assign io_ray_id_out = ~FIFO_0_empty ? FIFO_A_2_0_ray_io_dataout : _GEN_19; // @[Arbitration_2_1.scala 150:35 Arbitration_2_1.scala 151:55]
  assign io_hit_out = ~FIFO_0_empty ? FIFO_A_2_0_hit_io_dataout : _GEN_20; // @[Arbitration_2_1.scala 150:35 Arbitration_2_1.scala 152:59]
  assign io_valid_out = ~FIFO_0_empty ? valid_out_temp : _GEN_21; // @[Arbitration_2_1.scala 150:35 Arbitration_2_1.scala 153:57]
  assign FIFO_A_2_0_ray_clock = clock;
  assign FIFO_A_2_0_ray_reset = reset;
  assign FIFO_A_2_0_ray_io_datain = io_ray_id_2_0; // @[Arbitration_2_1.scala 52:43]
  assign FIFO_A_2_0_ray_io_wr = io_valid_2_0; // @[Arbitration_2_1.scala 50:47]
  assign FIFO_A_2_0_ray_io_rd = ~FIFO_A_2_0_ray_io_empty; // @[Arbitration_2_1.scala 75:38]
  assign FIFO_A_2_0_hit_clock = clock;
  assign FIFO_A_2_0_hit_reset = reset;
  assign FIFO_A_2_0_hit_io_datain = io_hit_2_0; // @[Arbitration_2_1.scala 53:44]
  assign FIFO_A_2_0_hit_io_wr = io_valid_2_0; // @[Arbitration_2_1.scala 51:48]
  assign FIFO_A_2_0_hit_io_rd = ~FIFO_A_2_0_ray_io_empty; // @[Arbitration_2_1.scala 75:38]
  assign FIFO_A_2_1_ray_clock = clock;
  assign FIFO_A_2_1_ray_reset = reset;
  assign FIFO_A_2_1_ray_io_datain = io_ray_id_2_1; // @[Arbitration_2_1.scala 57:43]
  assign FIFO_A_2_1_ray_io_wr = io_valid_2_1; // @[Arbitration_2_1.scala 55:47]
  assign FIFO_A_2_1_ray_io_rd = ~FIFO_A_2_0_ray_io_empty ? 1'h0 : _T_3; // @[Arbitration_2_1.scala 75:46 Arbitration_2_1.scala 78:47]
  assign FIFO_A_2_1_hit_clock = clock;
  assign FIFO_A_2_1_hit_reset = reset;
  assign FIFO_A_2_1_hit_io_datain = io_hit_2_1; // @[Arbitration_2_1.scala 58:44]
  assign FIFO_A_2_1_hit_io_wr = io_valid_2_1; // @[Arbitration_2_1.scala 56:48]
  assign FIFO_A_2_1_hit_io_rd = ~FIFO_A_2_0_ray_io_empty ? 1'h0 : _T_3; // @[Arbitration_2_1.scala 75:46 Arbitration_2_1.scala 78:47]
  assign FIFO_A_2_2_ray_clock = clock;
  assign FIFO_A_2_2_ray_reset = reset;
  assign FIFO_A_2_2_ray_io_datain = io_ray_id_2_2; // @[Arbitration_2_1.scala 62:43]
  assign FIFO_A_2_2_ray_io_wr = io_valid_2_2; // @[Arbitration_2_1.scala 60:47]
  assign FIFO_A_2_2_ray_io_rd = ~FIFO_A_2_0_ray_io_empty ? 1'h0 : _GEN_7; // @[Arbitration_2_1.scala 75:46 Arbitration_2_1.scala 80:47]
  assign FIFO_A_2_2_hit_clock = clock;
  assign FIFO_A_2_2_hit_reset = reset;
  assign FIFO_A_2_2_hit_io_datain = io_hit_2_2; // @[Arbitration_2_1.scala 63:44]
  assign FIFO_A_2_2_hit_io_wr = io_valid_2_2; // @[Arbitration_2_1.scala 61:48]
  assign FIFO_A_2_2_hit_io_rd = ~FIFO_A_2_0_ray_io_empty ? 1'h0 : _GEN_7; // @[Arbitration_2_1.scala 75:46 Arbitration_2_1.scala 80:47]
  assign FIFO_A_2_3_ray_clock = clock;
  assign FIFO_A_2_3_ray_reset = reset;
  assign FIFO_A_2_3_ray_io_datain = io_ray_id_2_3; // @[Arbitration_2_1.scala 67:43]
  assign FIFO_A_2_3_ray_io_wr = io_valid_2_3; // @[Arbitration_2_1.scala 65:47]
  assign FIFO_A_2_3_ray_io_rd = ~FIFO_A_2_0_ray_io_empty ? 1'h0 : _GEN_8; // @[Arbitration_2_1.scala 75:46 Arbitration_2_1.scala 82:47]
  assign FIFO_A_2_3_hit_clock = clock;
  assign FIFO_A_2_3_hit_reset = reset;
  assign FIFO_A_2_3_hit_io_datain = io_hit_2_3; // @[Arbitration_2_1.scala 68:44]
  assign FIFO_A_2_3_hit_io_wr = io_valid_2_3; // @[Arbitration_2_1.scala 66:48]
  assign FIFO_A_2_3_hit_io_rd = ~FIFO_A_2_0_ray_io_empty ? 1'h0 : _GEN_8; // @[Arbitration_2_1.scala 75:46 Arbitration_2_1.scala 82:47]
  always @(posedge clock) begin
    if (reset) begin // @[Arbitration_2_1.scala 73:59]
      valid_out_temp <= 1'h0; // @[Arbitration_2_1.scala 73:59]
    end else begin
      valid_out_temp <= FIFO_A_2_0_ray_io_rd | FIFO_A_2_1_ray_io_rd | FIFO_A_2_2_ray_io_rd | FIFO_A_2_3_ray_io_rd; // @[Arbitration_2_1.scala 149:51]
    end
    if (reset) begin // @[Arbitration_2_1.scala 121:58]
      FIFO_0_empty <= 1'h0; // @[Arbitration_2_1.scala 121:58]
    end else begin
      FIFO_0_empty <= FIFO_A_2_0_ray_io_empty; // @[Arbitration_2_1.scala 126:52]
    end
    if (reset) begin // @[Arbitration_2_1.scala 122:58]
      FIFO_1_empty <= 1'h0; // @[Arbitration_2_1.scala 122:58]
    end else begin
      FIFO_1_empty <= FIFO_A_2_1_ray_io_empty; // @[Arbitration_2_1.scala 127:52]
    end
    if (reset) begin // @[Arbitration_2_1.scala 123:58]
      FIFO_2_empty <= 1'h0; // @[Arbitration_2_1.scala 123:58]
    end else begin
      FIFO_2_empty <= FIFO_A_2_2_ray_io_empty; // @[Arbitration_2_1.scala 128:52]
    end
    if (reset) begin // @[Arbitration_2_1.scala 124:58]
      FIFO_3_empty <= 1'h0; // @[Arbitration_2_1.scala 124:58]
    end else begin
      FIFO_3_empty <= FIFO_A_2_3_ray_io_empty; // @[Arbitration_2_1.scala 129:52]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid_out_temp = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  FIFO_0_empty = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  FIFO_1_empty = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  FIFO_2_empty = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  FIFO_3_empty = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbitration_3(
  input         clock,
  input         reset,
  input  [31:0] io_node_id_3_0,
  input  [31:0] io_ray_id_3_0,
  input  [31:0] io_hit_3_0,
  input         io_valid_3_0,
  input  [31:0] io_node_id_3_1,
  input  [31:0] io_ray_id_3_1,
  input  [31:0] io_hit_3_1,
  input         io_valid_3_1,
  input  [31:0] io_node_id_3_2,
  input  [31:0] io_ray_id_3_2,
  input  [31:0] io_hit_3_2,
  input         io_valid_3_2,
  input  [31:0] io_node_id_3_3,
  input  [31:0] io_ray_id_3_3,
  input  [31:0] io_hit_3_3,
  input         io_valid_3_3,
  input  [31:0] io_node_id_3_4,
  input  [31:0] io_ray_id_3_4,
  input  [31:0] io_hit_3_4,
  input         io_valid_3_4,
  output [31:0] io_node_id_out,
  output [31:0] io_ray_id_out,
  output [31:0] io_hit_out,
  output        io_valid_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire  FIFO_A_3_0_node_clock; // @[Arbitration_3.scala 42:38]
  wire  FIFO_A_3_0_node_reset; // @[Arbitration_3.scala 42:38]
  wire [31:0] FIFO_A_3_0_node_io_datain; // @[Arbitration_3.scala 42:38]
  wire [31:0] FIFO_A_3_0_node_io_dataout; // @[Arbitration_3.scala 42:38]
  wire  FIFO_A_3_0_node_io_wr; // @[Arbitration_3.scala 42:38]
  wire  FIFO_A_3_0_node_io_rd; // @[Arbitration_3.scala 42:38]
  wire  FIFO_A_3_0_node_io_empty; // @[Arbitration_3.scala 42:38]
  wire  FIFO_A_3_0_ray_clock; // @[Arbitration_3.scala 43:41]
  wire  FIFO_A_3_0_ray_reset; // @[Arbitration_3.scala 43:41]
  wire [31:0] FIFO_A_3_0_ray_io_datain; // @[Arbitration_3.scala 43:41]
  wire [31:0] FIFO_A_3_0_ray_io_dataout; // @[Arbitration_3.scala 43:41]
  wire  FIFO_A_3_0_ray_io_wr; // @[Arbitration_3.scala 43:41]
  wire  FIFO_A_3_0_ray_io_rd; // @[Arbitration_3.scala 43:41]
  wire  FIFO_A_3_0_ray_io_empty; // @[Arbitration_3.scala 43:41]
  wire  FIFO_A_3_0_hit_clock; // @[Arbitration_3.scala 44:42]
  wire  FIFO_A_3_0_hit_reset; // @[Arbitration_3.scala 44:42]
  wire [31:0] FIFO_A_3_0_hit_io_datain; // @[Arbitration_3.scala 44:42]
  wire [31:0] FIFO_A_3_0_hit_io_dataout; // @[Arbitration_3.scala 44:42]
  wire  FIFO_A_3_0_hit_io_wr; // @[Arbitration_3.scala 44:42]
  wire  FIFO_A_3_0_hit_io_rd; // @[Arbitration_3.scala 44:42]
  wire  FIFO_A_3_0_hit_io_empty; // @[Arbitration_3.scala 44:42]
  wire  FIFO_A_3_1_node_clock; // @[Arbitration_3.scala 46:38]
  wire  FIFO_A_3_1_node_reset; // @[Arbitration_3.scala 46:38]
  wire [31:0] FIFO_A_3_1_node_io_datain; // @[Arbitration_3.scala 46:38]
  wire [31:0] FIFO_A_3_1_node_io_dataout; // @[Arbitration_3.scala 46:38]
  wire  FIFO_A_3_1_node_io_wr; // @[Arbitration_3.scala 46:38]
  wire  FIFO_A_3_1_node_io_rd; // @[Arbitration_3.scala 46:38]
  wire  FIFO_A_3_1_node_io_empty; // @[Arbitration_3.scala 46:38]
  wire  FIFO_A_3_1_ray_clock; // @[Arbitration_3.scala 47:41]
  wire  FIFO_A_3_1_ray_reset; // @[Arbitration_3.scala 47:41]
  wire [31:0] FIFO_A_3_1_ray_io_datain; // @[Arbitration_3.scala 47:41]
  wire [31:0] FIFO_A_3_1_ray_io_dataout; // @[Arbitration_3.scala 47:41]
  wire  FIFO_A_3_1_ray_io_wr; // @[Arbitration_3.scala 47:41]
  wire  FIFO_A_3_1_ray_io_rd; // @[Arbitration_3.scala 47:41]
  wire  FIFO_A_3_1_ray_io_empty; // @[Arbitration_3.scala 47:41]
  wire  FIFO_A_3_1_hit_clock; // @[Arbitration_3.scala 48:42]
  wire  FIFO_A_3_1_hit_reset; // @[Arbitration_3.scala 48:42]
  wire [31:0] FIFO_A_3_1_hit_io_datain; // @[Arbitration_3.scala 48:42]
  wire [31:0] FIFO_A_3_1_hit_io_dataout; // @[Arbitration_3.scala 48:42]
  wire  FIFO_A_3_1_hit_io_wr; // @[Arbitration_3.scala 48:42]
  wire  FIFO_A_3_1_hit_io_rd; // @[Arbitration_3.scala 48:42]
  wire  FIFO_A_3_1_hit_io_empty; // @[Arbitration_3.scala 48:42]
  wire  FIFO_A_3_2_node_clock; // @[Arbitration_3.scala 50:38]
  wire  FIFO_A_3_2_node_reset; // @[Arbitration_3.scala 50:38]
  wire [31:0] FIFO_A_3_2_node_io_datain; // @[Arbitration_3.scala 50:38]
  wire [31:0] FIFO_A_3_2_node_io_dataout; // @[Arbitration_3.scala 50:38]
  wire  FIFO_A_3_2_node_io_wr; // @[Arbitration_3.scala 50:38]
  wire  FIFO_A_3_2_node_io_rd; // @[Arbitration_3.scala 50:38]
  wire  FIFO_A_3_2_node_io_empty; // @[Arbitration_3.scala 50:38]
  wire  FIFO_A_3_2_ray_clock; // @[Arbitration_3.scala 51:41]
  wire  FIFO_A_3_2_ray_reset; // @[Arbitration_3.scala 51:41]
  wire [31:0] FIFO_A_3_2_ray_io_datain; // @[Arbitration_3.scala 51:41]
  wire [31:0] FIFO_A_3_2_ray_io_dataout; // @[Arbitration_3.scala 51:41]
  wire  FIFO_A_3_2_ray_io_wr; // @[Arbitration_3.scala 51:41]
  wire  FIFO_A_3_2_ray_io_rd; // @[Arbitration_3.scala 51:41]
  wire  FIFO_A_3_2_ray_io_empty; // @[Arbitration_3.scala 51:41]
  wire  FIFO_A_3_2_hit_clock; // @[Arbitration_3.scala 52:42]
  wire  FIFO_A_3_2_hit_reset; // @[Arbitration_3.scala 52:42]
  wire [31:0] FIFO_A_3_2_hit_io_datain; // @[Arbitration_3.scala 52:42]
  wire [31:0] FIFO_A_3_2_hit_io_dataout; // @[Arbitration_3.scala 52:42]
  wire  FIFO_A_3_2_hit_io_wr; // @[Arbitration_3.scala 52:42]
  wire  FIFO_A_3_2_hit_io_rd; // @[Arbitration_3.scala 52:42]
  wire  FIFO_A_3_2_hit_io_empty; // @[Arbitration_3.scala 52:42]
  wire  FIFO_A_3_3_node_clock; // @[Arbitration_3.scala 54:38]
  wire  FIFO_A_3_3_node_reset; // @[Arbitration_3.scala 54:38]
  wire [31:0] FIFO_A_3_3_node_io_datain; // @[Arbitration_3.scala 54:38]
  wire [31:0] FIFO_A_3_3_node_io_dataout; // @[Arbitration_3.scala 54:38]
  wire  FIFO_A_3_3_node_io_wr; // @[Arbitration_3.scala 54:38]
  wire  FIFO_A_3_3_node_io_rd; // @[Arbitration_3.scala 54:38]
  wire  FIFO_A_3_3_node_io_empty; // @[Arbitration_3.scala 54:38]
  wire  FIFO_A_3_3_ray_clock; // @[Arbitration_3.scala 55:41]
  wire  FIFO_A_3_3_ray_reset; // @[Arbitration_3.scala 55:41]
  wire [31:0] FIFO_A_3_3_ray_io_datain; // @[Arbitration_3.scala 55:41]
  wire [31:0] FIFO_A_3_3_ray_io_dataout; // @[Arbitration_3.scala 55:41]
  wire  FIFO_A_3_3_ray_io_wr; // @[Arbitration_3.scala 55:41]
  wire  FIFO_A_3_3_ray_io_rd; // @[Arbitration_3.scala 55:41]
  wire  FIFO_A_3_3_ray_io_empty; // @[Arbitration_3.scala 55:41]
  wire  FIFO_A_3_3_hit_clock; // @[Arbitration_3.scala 56:42]
  wire  FIFO_A_3_3_hit_reset; // @[Arbitration_3.scala 56:42]
  wire [31:0] FIFO_A_3_3_hit_io_datain; // @[Arbitration_3.scala 56:42]
  wire [31:0] FIFO_A_3_3_hit_io_dataout; // @[Arbitration_3.scala 56:42]
  wire  FIFO_A_3_3_hit_io_wr; // @[Arbitration_3.scala 56:42]
  wire  FIFO_A_3_3_hit_io_rd; // @[Arbitration_3.scala 56:42]
  wire  FIFO_A_3_3_hit_io_empty; // @[Arbitration_3.scala 56:42]
  wire  FIFO_A_3_4_node_clock; // @[Arbitration_3.scala 58:38]
  wire  FIFO_A_3_4_node_reset; // @[Arbitration_3.scala 58:38]
  wire [31:0] FIFO_A_3_4_node_io_datain; // @[Arbitration_3.scala 58:38]
  wire [31:0] FIFO_A_3_4_node_io_dataout; // @[Arbitration_3.scala 58:38]
  wire  FIFO_A_3_4_node_io_wr; // @[Arbitration_3.scala 58:38]
  wire  FIFO_A_3_4_node_io_rd; // @[Arbitration_3.scala 58:38]
  wire  FIFO_A_3_4_node_io_empty; // @[Arbitration_3.scala 58:38]
  wire  FIFO_A_3_4_ray_clock; // @[Arbitration_3.scala 59:41]
  wire  FIFO_A_3_4_ray_reset; // @[Arbitration_3.scala 59:41]
  wire [31:0] FIFO_A_3_4_ray_io_datain; // @[Arbitration_3.scala 59:41]
  wire [31:0] FIFO_A_3_4_ray_io_dataout; // @[Arbitration_3.scala 59:41]
  wire  FIFO_A_3_4_ray_io_wr; // @[Arbitration_3.scala 59:41]
  wire  FIFO_A_3_4_ray_io_rd; // @[Arbitration_3.scala 59:41]
  wire  FIFO_A_3_4_ray_io_empty; // @[Arbitration_3.scala 59:41]
  wire  FIFO_A_3_4_hit_clock; // @[Arbitration_3.scala 60:42]
  wire  FIFO_A_3_4_hit_reset; // @[Arbitration_3.scala 60:42]
  wire [31:0] FIFO_A_3_4_hit_io_datain; // @[Arbitration_3.scala 60:42]
  wire [31:0] FIFO_A_3_4_hit_io_dataout; // @[Arbitration_3.scala 60:42]
  wire  FIFO_A_3_4_hit_io_wr; // @[Arbitration_3.scala 60:42]
  wire  FIFO_A_3_4_hit_io_rd; // @[Arbitration_3.scala 60:42]
  wire  FIFO_A_3_4_hit_io_empty; // @[Arbitration_3.scala 60:42]
  reg  valid_out_temp; // @[Arbitration_3.scala 101:59]
  wire  _T_1 = FIFO_A_3_0_node_io_empty; // @[Arbitration_3.scala 119:45]
  wire  _T_3 = FIFO_A_3_0_node_io_empty & ~FIFO_A_3_1_node_io_empty; // @[Arbitration_3.scala 119:53]
  wire  _T_6 = _T_1 & FIFO_A_3_1_node_io_empty; // @[Arbitration_3.scala 135:53]
  wire  _T_8 = _T_1 & FIFO_A_3_1_node_io_empty & ~FIFO_A_3_2_node_io_empty; // @[Arbitration_3.scala 135:88]
  wire  _T_13 = _T_6 & FIFO_A_3_2_node_io_empty; // @[Arbitration_3.scala 151:88]
  wire  _T_15 = _T_6 & FIFO_A_3_2_node_io_empty & ~FIFO_A_3_3_node_io_empty; // @[Arbitration_3.scala 151:123]
  wire  _T_24 = _T_13 & FIFO_A_3_3_node_io_empty & ~FIFO_A_3_4_node_io_empty; // @[Arbitration_3.scala 167:157]
  wire  _GEN_4 = _T_6 & FIFO_A_3_2_node_io_empty & ~FIFO_A_3_3_node_io_empty ? 1'h0 : _T_24; // @[Arbitration_3.scala 151:158 Arbitration_3.scala 164:44]
  wire  _GEN_7 = _T_1 & FIFO_A_3_1_node_io_empty & ~FIFO_A_3_2_node_io_empty ? 1'h0 : _T_15; // @[Arbitration_3.scala 135:124 Arbitration_3.scala 145:44]
  wire  _GEN_8 = _T_1 & FIFO_A_3_1_node_io_empty & ~FIFO_A_3_2_node_io_empty ? 1'h0 : _GEN_4; // @[Arbitration_3.scala 135:124 Arbitration_3.scala 148:44]
  wire  _GEN_11 = FIFO_A_3_0_node_io_empty & ~FIFO_A_3_1_node_io_empty ? 1'h0 : _T_8; // @[Arbitration_3.scala 119:89 Arbitration_3.scala 126:44]
  wire  _GEN_12 = FIFO_A_3_0_node_io_empty & ~FIFO_A_3_1_node_io_empty ? 1'h0 : _GEN_7; // @[Arbitration_3.scala 119:89 Arbitration_3.scala 129:44]
  wire  _GEN_13 = FIFO_A_3_0_node_io_empty & ~FIFO_A_3_1_node_io_empty ? 1'h0 : _GEN_8; // @[Arbitration_3.scala 119:89 Arbitration_3.scala 132:44]
  reg  FIFO_0_empty; // @[Arbitration_3.scala 200:58]
  reg  FIFO_1_empty; // @[Arbitration_3.scala 201:58]
  reg  FIFO_2_empty; // @[Arbitration_3.scala 202:58]
  reg  FIFO_3_empty; // @[Arbitration_3.scala 203:58]
  reg  FIFO_4_empty; // @[Arbitration_3.scala 204:58]
  wire  _T_36 = FIFO_0_empty & FIFO_1_empty; // @[Arbitration_3.scala 237:40]
  wire  _T_43 = _T_36 & FIFO_2_empty; // @[Arbitration_3.scala 242:62]
  wire [31:0] _GEN_19 = _T_43 & FIFO_3_empty & ~FIFO_4_empty ? $signed(FIFO_A_3_4_node_io_dataout) : $signed(32'sh0); // @[Arbitration_3.scala 247:129 Arbitration_3.scala 248:46 Arbitration_3.scala 253:46]
  wire [31:0] _GEN_20 = _T_43 & FIFO_3_empty & ~FIFO_4_empty ? FIFO_A_3_4_ray_io_dataout : 32'h0; // @[Arbitration_3.scala 247:129 Arbitration_3.scala 249:48 Arbitration_3.scala 254:48]
  wire [31:0] _GEN_21 = _T_43 & FIFO_3_empty & ~FIFO_4_empty ? FIFO_A_3_4_hit_io_dataout : 32'h0; // @[Arbitration_3.scala 247:129 Arbitration_3.scala 250:52 Arbitration_3.scala 255:53]
  wire  _GEN_22 = _T_43 & FIFO_3_empty & ~FIFO_4_empty & valid_out_temp; // @[Arbitration_3.scala 247:129 Arbitration_3.scala 251:50 Arbitration_3.scala 256:50]
  wire [31:0] _GEN_23 = _T_36 & FIFO_2_empty & ~FIFO_3_empty ? $signed(FIFO_A_3_3_node_io_dataout) : $signed(_GEN_19); // @[Arbitration_3.scala 242:107 Arbitration_3.scala 243:46]
  wire [31:0] _GEN_24 = _T_36 & FIFO_2_empty & ~FIFO_3_empty ? FIFO_A_3_3_ray_io_dataout : _GEN_20; // @[Arbitration_3.scala 242:107 Arbitration_3.scala 244:47]
  wire [31:0] _GEN_25 = _T_36 & FIFO_2_empty & ~FIFO_3_empty ? FIFO_A_3_3_hit_io_dataout : _GEN_21; // @[Arbitration_3.scala 242:107 Arbitration_3.scala 245:53]
  wire  _GEN_26 = _T_36 & FIFO_2_empty & ~FIFO_3_empty ? valid_out_temp : _GEN_22; // @[Arbitration_3.scala 242:107 Arbitration_3.scala 246:50]
  wire [31:0] _GEN_27 = FIFO_0_empty & FIFO_1_empty & ~FIFO_2_empty ? $signed(FIFO_A_3_2_node_io_dataout) : $signed(
    _GEN_23); // @[Arbitration_3.scala 237:85 Arbitration_3.scala 238:46]
  wire [31:0] _GEN_28 = FIFO_0_empty & FIFO_1_empty & ~FIFO_2_empty ? FIFO_A_3_2_ray_io_dataout : _GEN_24; // @[Arbitration_3.scala 237:85 Arbitration_3.scala 239:48]
  wire [31:0] _GEN_29 = FIFO_0_empty & FIFO_1_empty & ~FIFO_2_empty ? FIFO_A_3_2_hit_io_dataout : _GEN_25; // @[Arbitration_3.scala 237:85 Arbitration_3.scala 240:53]
  wire  _GEN_30 = FIFO_0_empty & FIFO_1_empty & ~FIFO_2_empty ? valid_out_temp : _GEN_26; // @[Arbitration_3.scala 237:85 Arbitration_3.scala 241:50]
  wire [31:0] _GEN_31 = FIFO_0_empty & ~FIFO_1_empty ? $signed(FIFO_A_3_1_node_io_dataout) : $signed(_GEN_27); // @[Arbitration_3.scala 232:63 Arbitration_3.scala 233:45]
  wire [31:0] _GEN_32 = FIFO_0_empty & ~FIFO_1_empty ? FIFO_A_3_1_ray_io_dataout : _GEN_28; // @[Arbitration_3.scala 232:63 Arbitration_3.scala 234:48]
  wire [31:0] _GEN_33 = FIFO_0_empty & ~FIFO_1_empty ? FIFO_A_3_1_hit_io_dataout : _GEN_29; // @[Arbitration_3.scala 232:63 Arbitration_3.scala 235:53]
  wire  _GEN_34 = FIFO_0_empty & ~FIFO_1_empty ? valid_out_temp : _GEN_30; // @[Arbitration_3.scala 232:63 Arbitration_3.scala 236:50]
  FIFO FIFO_A_3_0_node ( // @[Arbitration_3.scala 42:38]
    .clock(FIFO_A_3_0_node_clock),
    .reset(FIFO_A_3_0_node_reset),
    .io_datain(FIFO_A_3_0_node_io_datain),
    .io_dataout(FIFO_A_3_0_node_io_dataout),
    .io_wr(FIFO_A_3_0_node_io_wr),
    .io_rd(FIFO_A_3_0_node_io_rd),
    .io_empty(FIFO_A_3_0_node_io_empty)
  );
  FIFO_0 FIFO_A_3_0_ray ( // @[Arbitration_3.scala 43:41]
    .clock(FIFO_A_3_0_ray_clock),
    .reset(FIFO_A_3_0_ray_reset),
    .io_datain(FIFO_A_3_0_ray_io_datain),
    .io_dataout(FIFO_A_3_0_ray_io_dataout),
    .io_wr(FIFO_A_3_0_ray_io_wr),
    .io_rd(FIFO_A_3_0_ray_io_rd),
    .io_empty(FIFO_A_3_0_ray_io_empty)
  );
  FIFO_0 FIFO_A_3_0_hit ( // @[Arbitration_3.scala 44:42]
    .clock(FIFO_A_3_0_hit_clock),
    .reset(FIFO_A_3_0_hit_reset),
    .io_datain(FIFO_A_3_0_hit_io_datain),
    .io_dataout(FIFO_A_3_0_hit_io_dataout),
    .io_wr(FIFO_A_3_0_hit_io_wr),
    .io_rd(FIFO_A_3_0_hit_io_rd),
    .io_empty(FIFO_A_3_0_hit_io_empty)
  );
  FIFO FIFO_A_3_1_node ( // @[Arbitration_3.scala 46:38]
    .clock(FIFO_A_3_1_node_clock),
    .reset(FIFO_A_3_1_node_reset),
    .io_datain(FIFO_A_3_1_node_io_datain),
    .io_dataout(FIFO_A_3_1_node_io_dataout),
    .io_wr(FIFO_A_3_1_node_io_wr),
    .io_rd(FIFO_A_3_1_node_io_rd),
    .io_empty(FIFO_A_3_1_node_io_empty)
  );
  FIFO_0 FIFO_A_3_1_ray ( // @[Arbitration_3.scala 47:41]
    .clock(FIFO_A_3_1_ray_clock),
    .reset(FIFO_A_3_1_ray_reset),
    .io_datain(FIFO_A_3_1_ray_io_datain),
    .io_dataout(FIFO_A_3_1_ray_io_dataout),
    .io_wr(FIFO_A_3_1_ray_io_wr),
    .io_rd(FIFO_A_3_1_ray_io_rd),
    .io_empty(FIFO_A_3_1_ray_io_empty)
  );
  FIFO_0 FIFO_A_3_1_hit ( // @[Arbitration_3.scala 48:42]
    .clock(FIFO_A_3_1_hit_clock),
    .reset(FIFO_A_3_1_hit_reset),
    .io_datain(FIFO_A_3_1_hit_io_datain),
    .io_dataout(FIFO_A_3_1_hit_io_dataout),
    .io_wr(FIFO_A_3_1_hit_io_wr),
    .io_rd(FIFO_A_3_1_hit_io_rd),
    .io_empty(FIFO_A_3_1_hit_io_empty)
  );
  FIFO FIFO_A_3_2_node ( // @[Arbitration_3.scala 50:38]
    .clock(FIFO_A_3_2_node_clock),
    .reset(FIFO_A_3_2_node_reset),
    .io_datain(FIFO_A_3_2_node_io_datain),
    .io_dataout(FIFO_A_3_2_node_io_dataout),
    .io_wr(FIFO_A_3_2_node_io_wr),
    .io_rd(FIFO_A_3_2_node_io_rd),
    .io_empty(FIFO_A_3_2_node_io_empty)
  );
  FIFO_0 FIFO_A_3_2_ray ( // @[Arbitration_3.scala 51:41]
    .clock(FIFO_A_3_2_ray_clock),
    .reset(FIFO_A_3_2_ray_reset),
    .io_datain(FIFO_A_3_2_ray_io_datain),
    .io_dataout(FIFO_A_3_2_ray_io_dataout),
    .io_wr(FIFO_A_3_2_ray_io_wr),
    .io_rd(FIFO_A_3_2_ray_io_rd),
    .io_empty(FIFO_A_3_2_ray_io_empty)
  );
  FIFO_0 FIFO_A_3_2_hit ( // @[Arbitration_3.scala 52:42]
    .clock(FIFO_A_3_2_hit_clock),
    .reset(FIFO_A_3_2_hit_reset),
    .io_datain(FIFO_A_3_2_hit_io_datain),
    .io_dataout(FIFO_A_3_2_hit_io_dataout),
    .io_wr(FIFO_A_3_2_hit_io_wr),
    .io_rd(FIFO_A_3_2_hit_io_rd),
    .io_empty(FIFO_A_3_2_hit_io_empty)
  );
  FIFO FIFO_A_3_3_node ( // @[Arbitration_3.scala 54:38]
    .clock(FIFO_A_3_3_node_clock),
    .reset(FIFO_A_3_3_node_reset),
    .io_datain(FIFO_A_3_3_node_io_datain),
    .io_dataout(FIFO_A_3_3_node_io_dataout),
    .io_wr(FIFO_A_3_3_node_io_wr),
    .io_rd(FIFO_A_3_3_node_io_rd),
    .io_empty(FIFO_A_3_3_node_io_empty)
  );
  FIFO_0 FIFO_A_3_3_ray ( // @[Arbitration_3.scala 55:41]
    .clock(FIFO_A_3_3_ray_clock),
    .reset(FIFO_A_3_3_ray_reset),
    .io_datain(FIFO_A_3_3_ray_io_datain),
    .io_dataout(FIFO_A_3_3_ray_io_dataout),
    .io_wr(FIFO_A_3_3_ray_io_wr),
    .io_rd(FIFO_A_3_3_ray_io_rd),
    .io_empty(FIFO_A_3_3_ray_io_empty)
  );
  FIFO_0 FIFO_A_3_3_hit ( // @[Arbitration_3.scala 56:42]
    .clock(FIFO_A_3_3_hit_clock),
    .reset(FIFO_A_3_3_hit_reset),
    .io_datain(FIFO_A_3_3_hit_io_datain),
    .io_dataout(FIFO_A_3_3_hit_io_dataout),
    .io_wr(FIFO_A_3_3_hit_io_wr),
    .io_rd(FIFO_A_3_3_hit_io_rd),
    .io_empty(FIFO_A_3_3_hit_io_empty)
  );
  FIFO FIFO_A_3_4_node ( // @[Arbitration_3.scala 58:38]
    .clock(FIFO_A_3_4_node_clock),
    .reset(FIFO_A_3_4_node_reset),
    .io_datain(FIFO_A_3_4_node_io_datain),
    .io_dataout(FIFO_A_3_4_node_io_dataout),
    .io_wr(FIFO_A_3_4_node_io_wr),
    .io_rd(FIFO_A_3_4_node_io_rd),
    .io_empty(FIFO_A_3_4_node_io_empty)
  );
  FIFO_0 FIFO_A_3_4_ray ( // @[Arbitration_3.scala 59:41]
    .clock(FIFO_A_3_4_ray_clock),
    .reset(FIFO_A_3_4_ray_reset),
    .io_datain(FIFO_A_3_4_ray_io_datain),
    .io_dataout(FIFO_A_3_4_ray_io_dataout),
    .io_wr(FIFO_A_3_4_ray_io_wr),
    .io_rd(FIFO_A_3_4_ray_io_rd),
    .io_empty(FIFO_A_3_4_ray_io_empty)
  );
  FIFO_0 FIFO_A_3_4_hit ( // @[Arbitration_3.scala 60:42]
    .clock(FIFO_A_3_4_hit_clock),
    .reset(FIFO_A_3_4_hit_reset),
    .io_datain(FIFO_A_3_4_hit_io_datain),
    .io_dataout(FIFO_A_3_4_hit_io_dataout),
    .io_wr(FIFO_A_3_4_hit_io_wr),
    .io_rd(FIFO_A_3_4_hit_io_rd),
    .io_empty(FIFO_A_3_4_hit_io_empty)
  );
  assign io_node_id_out = ~FIFO_0_empty ? $signed(FIFO_A_3_0_node_io_dataout) : $signed(_GEN_31); // @[Arbitration_3.scala 227:35 Arbitration_3.scala 228:46]
  assign io_ray_id_out = ~FIFO_0_empty ? FIFO_A_3_0_ray_io_dataout : _GEN_32; // @[Arbitration_3.scala 227:35 Arbitration_3.scala 229:48]
  assign io_hit_out = ~FIFO_0_empty ? FIFO_A_3_0_hit_io_dataout : _GEN_33; // @[Arbitration_3.scala 227:35 Arbitration_3.scala 230:53]
  assign io_valid_out = ~FIFO_0_empty ? valid_out_temp : _GEN_34; // @[Arbitration_3.scala 227:35 Arbitration_3.scala 231:50]
  assign FIFO_A_3_0_node_clock = clock;
  assign FIFO_A_3_0_node_reset = reset;
  assign FIFO_A_3_0_node_io_datain = io_node_id_3_0; // @[Arbitration_3.scala 66:40]
  assign FIFO_A_3_0_node_io_wr = io_valid_3_0; // @[Arbitration_3.scala 63:44]
  assign FIFO_A_3_0_node_io_rd = ~FIFO_A_3_0_node_io_empty; // @[Arbitration_3.scala 103:39]
  assign FIFO_A_3_0_ray_clock = clock;
  assign FIFO_A_3_0_ray_reset = reset;
  assign FIFO_A_3_0_ray_io_datain = io_ray_id_3_0; // @[Arbitration_3.scala 67:43]
  assign FIFO_A_3_0_ray_io_wr = io_valid_3_0; // @[Arbitration_3.scala 64:47]
  assign FIFO_A_3_0_ray_io_rd = ~FIFO_A_3_0_node_io_empty; // @[Arbitration_3.scala 103:39]
  assign FIFO_A_3_0_hit_clock = clock;
  assign FIFO_A_3_0_hit_reset = reset;
  assign FIFO_A_3_0_hit_io_datain = io_hit_3_0; // @[Arbitration_3.scala 68:44]
  assign FIFO_A_3_0_hit_io_wr = io_valid_3_0; // @[Arbitration_3.scala 65:48]
  assign FIFO_A_3_0_hit_io_rd = ~FIFO_A_3_0_node_io_empty; // @[Arbitration_3.scala 103:39]
  assign FIFO_A_3_1_node_clock = clock;
  assign FIFO_A_3_1_node_reset = reset;
  assign FIFO_A_3_1_node_io_datain = io_node_id_3_1; // @[Arbitration_3.scala 73:40]
  assign FIFO_A_3_1_node_io_wr = io_valid_3_1; // @[Arbitration_3.scala 70:44]
  assign FIFO_A_3_1_node_io_rd = ~FIFO_A_3_0_node_io_empty ? 1'h0 : _T_3; // @[Arbitration_3.scala 103:47 Arbitration_3.scala 107:44]
  assign FIFO_A_3_1_ray_clock = clock;
  assign FIFO_A_3_1_ray_reset = reset;
  assign FIFO_A_3_1_ray_io_datain = io_ray_id_3_1; // @[Arbitration_3.scala 74:43]
  assign FIFO_A_3_1_ray_io_wr = io_valid_3_1; // @[Arbitration_3.scala 71:47]
  assign FIFO_A_3_1_ray_io_rd = ~FIFO_A_3_0_node_io_empty ? 1'h0 : _T_3; // @[Arbitration_3.scala 103:47 Arbitration_3.scala 107:44]
  assign FIFO_A_3_1_hit_clock = clock;
  assign FIFO_A_3_1_hit_reset = reset;
  assign FIFO_A_3_1_hit_io_datain = io_hit_3_1; // @[Arbitration_3.scala 75:44]
  assign FIFO_A_3_1_hit_io_wr = io_valid_3_1; // @[Arbitration_3.scala 72:48]
  assign FIFO_A_3_1_hit_io_rd = ~FIFO_A_3_0_node_io_empty ? 1'h0 : _T_3; // @[Arbitration_3.scala 103:47 Arbitration_3.scala 107:44]
  assign FIFO_A_3_2_node_clock = clock;
  assign FIFO_A_3_2_node_reset = reset;
  assign FIFO_A_3_2_node_io_datain = io_node_id_3_2; // @[Arbitration_3.scala 80:40]
  assign FIFO_A_3_2_node_io_wr = io_valid_3_2; // @[Arbitration_3.scala 77:44]
  assign FIFO_A_3_2_node_io_rd = ~FIFO_A_3_0_node_io_empty ? 1'h0 : _GEN_11; // @[Arbitration_3.scala 103:47 Arbitration_3.scala 110:44]
  assign FIFO_A_3_2_ray_clock = clock;
  assign FIFO_A_3_2_ray_reset = reset;
  assign FIFO_A_3_2_ray_io_datain = io_ray_id_3_2; // @[Arbitration_3.scala 81:43]
  assign FIFO_A_3_2_ray_io_wr = io_valid_3_2; // @[Arbitration_3.scala 78:47]
  assign FIFO_A_3_2_ray_io_rd = ~FIFO_A_3_0_node_io_empty ? 1'h0 : _GEN_11; // @[Arbitration_3.scala 103:47 Arbitration_3.scala 110:44]
  assign FIFO_A_3_2_hit_clock = clock;
  assign FIFO_A_3_2_hit_reset = reset;
  assign FIFO_A_3_2_hit_io_datain = io_hit_3_2; // @[Arbitration_3.scala 82:44]
  assign FIFO_A_3_2_hit_io_wr = io_valid_3_2; // @[Arbitration_3.scala 79:48]
  assign FIFO_A_3_2_hit_io_rd = ~FIFO_A_3_0_node_io_empty ? 1'h0 : _GEN_11; // @[Arbitration_3.scala 103:47 Arbitration_3.scala 110:44]
  assign FIFO_A_3_3_node_clock = clock;
  assign FIFO_A_3_3_node_reset = reset;
  assign FIFO_A_3_3_node_io_datain = io_node_id_3_3; // @[Arbitration_3.scala 87:40]
  assign FIFO_A_3_3_node_io_wr = io_valid_3_3; // @[Arbitration_3.scala 84:44]
  assign FIFO_A_3_3_node_io_rd = ~FIFO_A_3_0_node_io_empty ? 1'h0 : _GEN_12; // @[Arbitration_3.scala 103:47 Arbitration_3.scala 113:44]
  assign FIFO_A_3_3_ray_clock = clock;
  assign FIFO_A_3_3_ray_reset = reset;
  assign FIFO_A_3_3_ray_io_datain = io_ray_id_3_3; // @[Arbitration_3.scala 88:43]
  assign FIFO_A_3_3_ray_io_wr = io_valid_3_3; // @[Arbitration_3.scala 85:47]
  assign FIFO_A_3_3_ray_io_rd = ~FIFO_A_3_0_node_io_empty ? 1'h0 : _GEN_12; // @[Arbitration_3.scala 103:47 Arbitration_3.scala 113:44]
  assign FIFO_A_3_3_hit_clock = clock;
  assign FIFO_A_3_3_hit_reset = reset;
  assign FIFO_A_3_3_hit_io_datain = io_hit_3_3; // @[Arbitration_3.scala 89:44]
  assign FIFO_A_3_3_hit_io_wr = io_valid_3_3; // @[Arbitration_3.scala 86:48]
  assign FIFO_A_3_3_hit_io_rd = ~FIFO_A_3_0_node_io_empty ? 1'h0 : _GEN_12; // @[Arbitration_3.scala 103:47 Arbitration_3.scala 113:44]
  assign FIFO_A_3_4_node_clock = clock;
  assign FIFO_A_3_4_node_reset = reset;
  assign FIFO_A_3_4_node_io_datain = io_node_id_3_4; // @[Arbitration_3.scala 94:40]
  assign FIFO_A_3_4_node_io_wr = io_valid_3_4; // @[Arbitration_3.scala 91:44]
  assign FIFO_A_3_4_node_io_rd = ~FIFO_A_3_0_node_io_empty ? 1'h0 : _GEN_13; // @[Arbitration_3.scala 103:47 Arbitration_3.scala 116:44]
  assign FIFO_A_3_4_ray_clock = clock;
  assign FIFO_A_3_4_ray_reset = reset;
  assign FIFO_A_3_4_ray_io_datain = io_ray_id_3_4; // @[Arbitration_3.scala 95:43]
  assign FIFO_A_3_4_ray_io_wr = io_valid_3_4; // @[Arbitration_3.scala 92:47]
  assign FIFO_A_3_4_ray_io_rd = ~FIFO_A_3_0_node_io_empty ? 1'h0 : _GEN_13; // @[Arbitration_3.scala 103:47 Arbitration_3.scala 116:44]
  assign FIFO_A_3_4_hit_clock = clock;
  assign FIFO_A_3_4_hit_reset = reset;
  assign FIFO_A_3_4_hit_io_datain = io_hit_3_4; // @[Arbitration_3.scala 96:44]
  assign FIFO_A_3_4_hit_io_wr = io_valid_3_4; // @[Arbitration_3.scala 93:48]
  assign FIFO_A_3_4_hit_io_rd = ~FIFO_A_3_0_node_io_empty ? 1'h0 : _GEN_13; // @[Arbitration_3.scala 103:47 Arbitration_3.scala 116:44]
  always @(posedge clock) begin
    if (reset) begin // @[Arbitration_3.scala 101:59]
      valid_out_temp <= 1'h0; // @[Arbitration_3.scala 101:59]
    end else begin
      valid_out_temp <= FIFO_A_3_0_node_io_rd | FIFO_A_3_1_node_io_rd | FIFO_A_3_2_node_io_rd | FIFO_A_3_3_node_io_rd |
        FIFO_A_3_4_node_io_rd; // @[Arbitration_3.scala 225:51]
    end
    if (reset) begin // @[Arbitration_3.scala 200:58]
      FIFO_0_empty <= 1'h0; // @[Arbitration_3.scala 200:58]
    end else begin
      FIFO_0_empty <= FIFO_A_3_0_node_io_empty; // @[Arbitration_3.scala 206:52]
    end
    if (reset) begin // @[Arbitration_3.scala 201:58]
      FIFO_1_empty <= 1'h0; // @[Arbitration_3.scala 201:58]
    end else begin
      FIFO_1_empty <= FIFO_A_3_1_node_io_empty; // @[Arbitration_3.scala 207:52]
    end
    if (reset) begin // @[Arbitration_3.scala 202:58]
      FIFO_2_empty <= 1'h0; // @[Arbitration_3.scala 202:58]
    end else begin
      FIFO_2_empty <= FIFO_A_3_2_node_io_empty; // @[Arbitration_3.scala 208:52]
    end
    if (reset) begin // @[Arbitration_3.scala 203:58]
      FIFO_3_empty <= 1'h0; // @[Arbitration_3.scala 203:58]
    end else begin
      FIFO_3_empty <= FIFO_A_3_3_node_io_empty; // @[Arbitration_3.scala 209:52]
    end
    if (reset) begin // @[Arbitration_3.scala 204:58]
      FIFO_4_empty <= 1'h0; // @[Arbitration_3.scala 204:58]
    end else begin
      FIFO_4_empty <= FIFO_A_3_4_node_io_empty; // @[Arbitration_3.scala 210:52]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid_out_temp = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  FIFO_0_empty = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  FIFO_1_empty = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  FIFO_2_empty = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  FIFO_3_empty = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  FIFO_4_empty = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FSM_1(
  input   clock,
  input   reset,
  input   io_request_0,
  input   io_request_1,
  output  io_grant_0,
  output  io_grant_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] grant; // @[FSM.scala 18:26]
  reg [1:0] stateReg; // @[FSM.scala 19:23]
  wire  _T = 2'h0 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_4 = ~io_request_1; // @[FSM.scala 29:44]
  wire [1:0] _GEN_2 = ~io_request_0 & io_request_1 ? 2'h2 : 2'h0; // @[FSM.scala 26:56 FSM.scala 27:27]
  wire [1:0] _GEN_4 = io_request_0 ? 2'h1 : _GEN_2; // @[FSM.scala 23:31 FSM.scala 24:27]
  wire  _T_6 = 2'h1 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_8 = _T_4 & io_request_0; // @[FSM.scala 41:39]
  wire  _T_12 = 2'h2 == stateReg; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_16 = io_request_0 ? 2'h1 : 2'h2; // @[FSM.scala 53:31 FSM.scala 54:27]
  assign io_grant_0 = grant == 2'h1; // @[FSM.scala 90:38]
  assign io_grant_1 = grant == 2'h2; // @[FSM.scala 91:38]
  always @(posedge clock) begin
    if (reset) begin // @[FSM.scala 18:26]
      grant <= 2'h0; // @[FSM.scala 18:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      grant <= _GEN_4;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      if (io_request_1) begin // @[FSM.scala 38:31]
        grant <= 2'h2; // @[FSM.scala 40:31]
      end else begin
        grant <= {{1'd0}, _T_8};
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      grant <= _GEN_4;
    end
    if (reset) begin // @[FSM.scala 19:23]
      stateReg <= 2'h0; // @[FSM.scala 19:23]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_request_0) begin // @[FSM.scala 23:31]
        stateReg <= 2'h1; // @[FSM.scala 24:27]
      end else if (~io_request_0 & io_request_1) begin // @[FSM.scala 26:56]
        stateReg <= 2'h2; // @[FSM.scala 27:27]
      end else begin
        stateReg <= 2'h0;
      end
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      if (io_request_1) begin // @[FSM.scala 38:31]
        stateReg <= 2'h2; // @[FSM.scala 39:27]
      end else begin
        stateReg <= 2'h1;
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      stateReg <= _GEN_16;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  grant = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  stateReg = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbitration_4(
  input         clock,
  input         reset,
  input  [31:0] io_node_id_4_0,
  input  [31:0] io_ray_id_4_0,
  input  [31:0] io_hit_4_0,
  input         io_valid_4_0,
  input  [31:0] io_node_id_4_1,
  input  [31:0] io_ray_id_4_1,
  input  [31:0] io_hit_4_1,
  input         io_valid_4_1,
  output [31:0] io_node_id_out,
  output [31:0] io_ray_id_out,
  output [31:0] io_hit_out,
  output        io_RAY_AABB_out,
  output        io_RAY_AABB_2_out,
  output        io_valid_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  FSM_clock; // @[Arbitration_4.scala 31:55]
  wire  FSM_reset; // @[Arbitration_4.scala 31:55]
  wire  FSM_io_request_0; // @[Arbitration_4.scala 31:55]
  wire  FSM_io_request_1; // @[Arbitration_4.scala 31:55]
  wire  FSM_io_grant_0; // @[Arbitration_4.scala 31:55]
  wire  FSM_io_grant_1; // @[Arbitration_4.scala 31:55]
  wire  FIFO_A_4_0_node_clock; // @[Arbitration_4.scala 33:38]
  wire  FIFO_A_4_0_node_reset; // @[Arbitration_4.scala 33:38]
  wire [31:0] FIFO_A_4_0_node_io_datain; // @[Arbitration_4.scala 33:38]
  wire [31:0] FIFO_A_4_0_node_io_dataout; // @[Arbitration_4.scala 33:38]
  wire  FIFO_A_4_0_node_io_wr; // @[Arbitration_4.scala 33:38]
  wire  FIFO_A_4_0_node_io_rd; // @[Arbitration_4.scala 33:38]
  wire  FIFO_A_4_0_node_io_empty; // @[Arbitration_4.scala 33:38]
  wire  FIFO_A_4_0_ray_clock; // @[Arbitration_4.scala 34:41]
  wire  FIFO_A_4_0_ray_reset; // @[Arbitration_4.scala 34:41]
  wire [31:0] FIFO_A_4_0_ray_io_datain; // @[Arbitration_4.scala 34:41]
  wire [31:0] FIFO_A_4_0_ray_io_dataout; // @[Arbitration_4.scala 34:41]
  wire  FIFO_A_4_0_ray_io_wr; // @[Arbitration_4.scala 34:41]
  wire  FIFO_A_4_0_ray_io_rd; // @[Arbitration_4.scala 34:41]
  wire  FIFO_A_4_0_ray_io_empty; // @[Arbitration_4.scala 34:41]
  wire  FIFO_A_4_0_hit_clock; // @[Arbitration_4.scala 35:42]
  wire  FIFO_A_4_0_hit_reset; // @[Arbitration_4.scala 35:42]
  wire [31:0] FIFO_A_4_0_hit_io_datain; // @[Arbitration_4.scala 35:42]
  wire [31:0] FIFO_A_4_0_hit_io_dataout; // @[Arbitration_4.scala 35:42]
  wire  FIFO_A_4_0_hit_io_wr; // @[Arbitration_4.scala 35:42]
  wire  FIFO_A_4_0_hit_io_rd; // @[Arbitration_4.scala 35:42]
  wire  FIFO_A_4_0_hit_io_empty; // @[Arbitration_4.scala 35:42]
  wire  FIFO_A_4_1_node_clock; // @[Arbitration_4.scala 37:38]
  wire  FIFO_A_4_1_node_reset; // @[Arbitration_4.scala 37:38]
  wire [31:0] FIFO_A_4_1_node_io_datain; // @[Arbitration_4.scala 37:38]
  wire [31:0] FIFO_A_4_1_node_io_dataout; // @[Arbitration_4.scala 37:38]
  wire  FIFO_A_4_1_node_io_wr; // @[Arbitration_4.scala 37:38]
  wire  FIFO_A_4_1_node_io_rd; // @[Arbitration_4.scala 37:38]
  wire  FIFO_A_4_1_node_io_empty; // @[Arbitration_4.scala 37:38]
  wire  FIFO_A_4_1_ray_clock; // @[Arbitration_4.scala 38:41]
  wire  FIFO_A_4_1_ray_reset; // @[Arbitration_4.scala 38:41]
  wire [31:0] FIFO_A_4_1_ray_io_datain; // @[Arbitration_4.scala 38:41]
  wire [31:0] FIFO_A_4_1_ray_io_dataout; // @[Arbitration_4.scala 38:41]
  wire  FIFO_A_4_1_ray_io_wr; // @[Arbitration_4.scala 38:41]
  wire  FIFO_A_4_1_ray_io_rd; // @[Arbitration_4.scala 38:41]
  wire  FIFO_A_4_1_ray_io_empty; // @[Arbitration_4.scala 38:41]
  wire  FIFO_A_4_1_hit_clock; // @[Arbitration_4.scala 39:42]
  wire  FIFO_A_4_1_hit_reset; // @[Arbitration_4.scala 39:42]
  wire [31:0] FIFO_A_4_1_hit_io_datain; // @[Arbitration_4.scala 39:42]
  wire [31:0] FIFO_A_4_1_hit_io_dataout; // @[Arbitration_4.scala 39:42]
  wire  FIFO_A_4_1_hit_io_wr; // @[Arbitration_4.scala 39:42]
  wire  FIFO_A_4_1_hit_io_rd; // @[Arbitration_4.scala 39:42]
  wire  FIFO_A_4_1_hit_io_empty; // @[Arbitration_4.scala 39:42]
  wire  _T = ~FIFO_A_4_0_ray_io_empty; // @[Arbitration_4.scala 59:76]
  wire  _T_1 = ~FIFO_A_4_1_ray_io_empty; // @[Arbitration_4.scala 60:76]
  reg  valid_0; // @[Arbitration_4.scala 61:66]
  reg  valid_1; // @[Arbitration_4.scala 62:66]
  wire  _T_3 = FSM_io_grant_0 & _T; // @[Arbitration_4.scala 63:28]
  wire  _T_5 = FSM_io_grant_1 & _T_1; // @[Arbitration_4.scala 72:35]
  wire [31:0] _GEN_4 = valid_1 ? $signed(FIFO_A_4_1_node_io_dataout) : $signed(32'sh0); // @[Arbitration_4.scala 134:34 Arbitration_4.scala 135:45 Arbitration_4.scala 151:46]
  wire [31:0] _GEN_5 = valid_1 ? FIFO_A_4_1_ray_io_dataout : 32'h0; // @[Arbitration_4.scala 134:34 Arbitration_4.scala 136:48 Arbitration_4.scala 152:48]
  wire [31:0] _GEN_6 = valid_1 ? FIFO_A_4_1_hit_io_dataout : 32'h0; // @[Arbitration_4.scala 134:34 Arbitration_4.scala 137:53 Arbitration_4.scala 153:53]
  FSM_1 FSM ( // @[Arbitration_4.scala 31:55]
    .clock(FSM_clock),
    .reset(FSM_reset),
    .io_request_0(FSM_io_request_0),
    .io_request_1(FSM_io_request_1),
    .io_grant_0(FSM_io_grant_0),
    .io_grant_1(FSM_io_grant_1)
  );
  FIFO FIFO_A_4_0_node ( // @[Arbitration_4.scala 33:38]
    .clock(FIFO_A_4_0_node_clock),
    .reset(FIFO_A_4_0_node_reset),
    .io_datain(FIFO_A_4_0_node_io_datain),
    .io_dataout(FIFO_A_4_0_node_io_dataout),
    .io_wr(FIFO_A_4_0_node_io_wr),
    .io_rd(FIFO_A_4_0_node_io_rd),
    .io_empty(FIFO_A_4_0_node_io_empty)
  );
  FIFO_0 FIFO_A_4_0_ray ( // @[Arbitration_4.scala 34:41]
    .clock(FIFO_A_4_0_ray_clock),
    .reset(FIFO_A_4_0_ray_reset),
    .io_datain(FIFO_A_4_0_ray_io_datain),
    .io_dataout(FIFO_A_4_0_ray_io_dataout),
    .io_wr(FIFO_A_4_0_ray_io_wr),
    .io_rd(FIFO_A_4_0_ray_io_rd),
    .io_empty(FIFO_A_4_0_ray_io_empty)
  );
  FIFO_0 FIFO_A_4_0_hit ( // @[Arbitration_4.scala 35:42]
    .clock(FIFO_A_4_0_hit_clock),
    .reset(FIFO_A_4_0_hit_reset),
    .io_datain(FIFO_A_4_0_hit_io_datain),
    .io_dataout(FIFO_A_4_0_hit_io_dataout),
    .io_wr(FIFO_A_4_0_hit_io_wr),
    .io_rd(FIFO_A_4_0_hit_io_rd),
    .io_empty(FIFO_A_4_0_hit_io_empty)
  );
  FIFO FIFO_A_4_1_node ( // @[Arbitration_4.scala 37:38]
    .clock(FIFO_A_4_1_node_clock),
    .reset(FIFO_A_4_1_node_reset),
    .io_datain(FIFO_A_4_1_node_io_datain),
    .io_dataout(FIFO_A_4_1_node_io_dataout),
    .io_wr(FIFO_A_4_1_node_io_wr),
    .io_rd(FIFO_A_4_1_node_io_rd),
    .io_empty(FIFO_A_4_1_node_io_empty)
  );
  FIFO_0 FIFO_A_4_1_ray ( // @[Arbitration_4.scala 38:41]
    .clock(FIFO_A_4_1_ray_clock),
    .reset(FIFO_A_4_1_ray_reset),
    .io_datain(FIFO_A_4_1_ray_io_datain),
    .io_dataout(FIFO_A_4_1_ray_io_dataout),
    .io_wr(FIFO_A_4_1_ray_io_wr),
    .io_rd(FIFO_A_4_1_ray_io_rd),
    .io_empty(FIFO_A_4_1_ray_io_empty)
  );
  FIFO_0 FIFO_A_4_1_hit ( // @[Arbitration_4.scala 39:42]
    .clock(FIFO_A_4_1_hit_clock),
    .reset(FIFO_A_4_1_hit_reset),
    .io_datain(FIFO_A_4_1_hit_io_datain),
    .io_dataout(FIFO_A_4_1_hit_io_dataout),
    .io_wr(FIFO_A_4_1_hit_io_wr),
    .io_rd(FIFO_A_4_1_hit_io_rd),
    .io_empty(FIFO_A_4_1_hit_io_empty)
  );
  assign io_node_id_out = valid_0 ? $signed(FIFO_A_4_0_node_io_dataout) : $signed(_GEN_4); // @[Arbitration_4.scala 126:29 Arbitration_4.scala 127:46]
  assign io_ray_id_out = valid_0 ? FIFO_A_4_0_ray_io_dataout : _GEN_5; // @[Arbitration_4.scala 126:29 Arbitration_4.scala 128:48]
  assign io_hit_out = valid_0 ? FIFO_A_4_0_hit_io_dataout : _GEN_6; // @[Arbitration_4.scala 126:29 Arbitration_4.scala 129:53]
  assign io_RAY_AABB_out = valid_0; // @[Arbitration_4.scala 126:29 Arbitration_4.scala 131:41]
  assign io_RAY_AABB_2_out = valid_0 ? 1'h0 : valid_1; // @[Arbitration_4.scala 126:29 Arbitration_4.scala 132:38]
  assign io_valid_out = valid_0 | valid_1; // @[Arbitration_4.scala 126:29 Arbitration_4.scala 130:50]
  assign FSM_clock = clock;
  assign FSM_reset = reset;
  assign FSM_io_request_0 = ~FIFO_A_4_0_ray_io_empty; // @[Arbitration_4.scala 59:76]
  assign FSM_io_request_1 = ~FIFO_A_4_1_ray_io_empty; // @[Arbitration_4.scala 60:76]
  assign FIFO_A_4_0_node_clock = clock;
  assign FIFO_A_4_0_node_reset = reset;
  assign FIFO_A_4_0_node_io_datain = io_node_id_4_0; // @[Arbitration_4.scala 44:40]
  assign FIFO_A_4_0_node_io_wr = io_valid_4_0; // @[Arbitration_4.scala 41:44]
  assign FIFO_A_4_0_node_io_rd = FSM_io_grant_0 & _T; // @[Arbitration_4.scala 63:28]
  assign FIFO_A_4_0_ray_clock = clock;
  assign FIFO_A_4_0_ray_reset = reset;
  assign FIFO_A_4_0_ray_io_datain = io_ray_id_4_0; // @[Arbitration_4.scala 45:43]
  assign FIFO_A_4_0_ray_io_wr = io_valid_4_0; // @[Arbitration_4.scala 42:47]
  assign FIFO_A_4_0_ray_io_rd = FSM_io_grant_0 & _T; // @[Arbitration_4.scala 63:28]
  assign FIFO_A_4_0_hit_clock = clock;
  assign FIFO_A_4_0_hit_reset = reset;
  assign FIFO_A_4_0_hit_io_datain = io_hit_4_0; // @[Arbitration_4.scala 46:44]
  assign FIFO_A_4_0_hit_io_wr = io_valid_4_0; // @[Arbitration_4.scala 43:48]
  assign FIFO_A_4_0_hit_io_rd = FSM_io_grant_0 & _T; // @[Arbitration_4.scala 63:28]
  assign FIFO_A_4_1_node_clock = clock;
  assign FIFO_A_4_1_node_reset = reset;
  assign FIFO_A_4_1_node_io_datain = io_node_id_4_1; // @[Arbitration_4.scala 51:40]
  assign FIFO_A_4_1_node_io_wr = io_valid_4_1; // @[Arbitration_4.scala 48:44]
  assign FIFO_A_4_1_node_io_rd = FSM_io_grant_0 & _T ? 1'h0 : _T_5; // @[Arbitration_4.scala 63:57 Arbitration_4.scala 67:44]
  assign FIFO_A_4_1_ray_clock = clock;
  assign FIFO_A_4_1_ray_reset = reset;
  assign FIFO_A_4_1_ray_io_datain = io_ray_id_4_1; // @[Arbitration_4.scala 52:43]
  assign FIFO_A_4_1_ray_io_wr = io_valid_4_1; // @[Arbitration_4.scala 49:47]
  assign FIFO_A_4_1_ray_io_rd = FSM_io_grant_0 & _T ? 1'h0 : _T_5; // @[Arbitration_4.scala 63:57 Arbitration_4.scala 67:44]
  assign FIFO_A_4_1_hit_clock = clock;
  assign FIFO_A_4_1_hit_reset = reset;
  assign FIFO_A_4_1_hit_io_datain = io_hit_4_1; // @[Arbitration_4.scala 53:44]
  assign FIFO_A_4_1_hit_io_wr = io_valid_4_1; // @[Arbitration_4.scala 50:48]
  assign FIFO_A_4_1_hit_io_rd = FSM_io_grant_0 & _T ? 1'h0 : _T_5; // @[Arbitration_4.scala 63:57 Arbitration_4.scala 67:44]
  always @(posedge clock) begin
    if (reset) begin // @[Arbitration_4.scala 61:66]
      valid_0 <= 1'h0; // @[Arbitration_4.scala 61:66]
    end else begin
      valid_0 <= _T_3;
    end
    if (reset) begin // @[Arbitration_4.scala 62:66]
      valid_1 <= 1'h0; // @[Arbitration_4.scala 62:66]
    end else if (FSM_io_grant_0 & _T) begin // @[Arbitration_4.scala 63:57]
      valid_1 <= 1'h0; // @[Arbitration_4.scala 67:44]
    end else begin
      valid_1 <= _T_5;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  valid_1 = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LUT(
  input         clock,
  input         reset,
  input         io_push,
  input         io_push_valid,
  input         io_pop,
  input         io_pop_valid,
  input         io_empty_0,
  input         io_empty_1,
  input         io_empty_2,
  input         io_empty_3,
  input         io_empty_4,
  input         io_empty_5,
  input         io_empty_6,
  input         io_empty_7,
  input         io_empty_8,
  input         io_empty_9,
  input         io_empty_10,
  input         io_empty_11,
  input         io_empty_12,
  input         io_empty_13,
  input         io_empty_14,
  input         io_empty_15,
  input         io_empty_16,
  input         io_empty_17,
  input         io_empty_18,
  input         io_empty_19,
  input         io_empty_20,
  input         io_empty_21,
  input         io_empty_22,
  input         io_empty_23,
  input         io_empty_24,
  input         io_empty_25,
  input         io_empty_26,
  input         io_empty_27,
  input         io_empty_28,
  input         io_empty_29,
  input         io_empty_30,
  input         io_empty_31,
  input         io_empty_32,
  input         io_empty_33,
  input         io_empty_34,
  input         io_dispatch_0,
  input         io_dispatch_1,
  input         io_dispatch_2,
  input         io_dispatch_3,
  input         io_dispatch_4,
  input         io_dispatch_5,
  input         io_dispatch_6,
  input         io_dispatch_7,
  input         io_dispatch_8,
  input         io_dispatch_9,
  input         io_dispatch_10,
  input         io_dispatch_11,
  input         io_dispatch_12,
  input         io_dispatch_13,
  input         io_dispatch_14,
  input         io_dispatch_15,
  input         io_dispatch_16,
  input         io_dispatch_17,
  input         io_dispatch_18,
  input         io_dispatch_19,
  input         io_dispatch_20,
  input         io_dispatch_21,
  input         io_dispatch_22,
  input         io_dispatch_23,
  input         io_dispatch_24,
  input         io_dispatch_25,
  input         io_dispatch_26,
  input         io_dispatch_27,
  input         io_dispatch_28,
  input         io_dispatch_29,
  input         io_dispatch_30,
  input         io_dispatch_31,
  input         io_dispatch_32,
  input         io_dispatch_33,
  input         io_dispatch_34,
  input  [31:0] io_ray_id_push,
  input  [31:0] io_ray_id_pop,
  input  [31:0] io_node_id_push_in,
  input  [31:0] io_hitT_in,
  output [31:0] io_ray_id_pop_out,
  output [31:0] io_hitT_out,
  output        io_pop_0,
  output        io_pop_1,
  output        io_pop_2,
  output        io_pop_3,
  output        io_pop_4,
  output        io_pop_5,
  output        io_pop_6,
  output        io_pop_7,
  output        io_pop_8,
  output        io_pop_9,
  output        io_pop_10,
  output        io_pop_11,
  output        io_pop_12,
  output        io_pop_13,
  output        io_pop_14,
  output        io_pop_15,
  output        io_pop_16,
  output        io_pop_17,
  output        io_pop_18,
  output        io_pop_19,
  output        io_pop_20,
  output        io_pop_21,
  output        io_pop_22,
  output        io_pop_23,
  output        io_pop_24,
  output        io_pop_25,
  output        io_pop_26,
  output        io_pop_27,
  output        io_pop_28,
  output        io_pop_29,
  output        io_pop_30,
  output        io_pop_31,
  output        io_pop_32,
  output        io_pop_33,
  output        io_pop_34,
  output        io_pop_en,
  output        io_push_0,
  output        io_push_1,
  output        io_push_2,
  output        io_push_3,
  output        io_push_4,
  output        io_push_5,
  output        io_push_6,
  output        io_push_7,
  output        io_push_8,
  output        io_push_9,
  output        io_push_10,
  output        io_push_11,
  output        io_push_12,
  output        io_push_13,
  output        io_push_14,
  output        io_push_15,
  output        io_push_16,
  output        io_push_17,
  output        io_push_18,
  output        io_push_19,
  output        io_push_20,
  output        io_push_21,
  output        io_push_22,
  output        io_push_23,
  output        io_push_24,
  output        io_push_25,
  output        io_push_26,
  output        io_push_27,
  output        io_push_28,
  output        io_push_29,
  output        io_push_30,
  output        io_push_31,
  output        io_push_32,
  output        io_push_33,
  output        io_push_34,
  output        io_push_en,
  output        io_no_match
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [63:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [63:0] _RAND_62;
  reg [63:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [63:0] _RAND_65;
  reg [63:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [63:0] _RAND_68;
  reg [63:0] _RAND_69;
  reg [63:0] _RAND_70;
  reg [63:0] _RAND_71;
  reg [63:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [63:0] _RAND_74;
  reg [63:0] _RAND_75;
  reg [63:0] _RAND_76;
  reg [63:0] _RAND_77;
  reg [63:0] _RAND_78;
  reg [63:0] _RAND_79;
  reg [63:0] _RAND_80;
  reg [63:0] _RAND_81;
  reg [63:0] _RAND_82;
  reg [63:0] _RAND_83;
  reg [63:0] _RAND_84;
  reg [63:0] _RAND_85;
  reg [63:0] _RAND_86;
  reg [63:0] _RAND_87;
  reg [63:0] _RAND_88;
  reg [63:0] _RAND_89;
  reg [63:0] _RAND_90;
  reg [63:0] _RAND_91;
  reg [63:0] _RAND_92;
  reg [63:0] _RAND_93;
  reg [63:0] _RAND_94;
  reg [63:0] _RAND_95;
  reg [63:0] _RAND_96;
  reg [63:0] _RAND_97;
  reg [63:0] _RAND_98;
  reg [63:0] _RAND_99;
  reg [63:0] _RAND_100;
  reg [63:0] _RAND_101;
  reg [63:0] _RAND_102;
  reg [63:0] _RAND_103;
  reg [63:0] _RAND_104;
  reg [63:0] _RAND_105;
  reg [63:0] _RAND_106;
  reg [63:0] _RAND_107;
  reg [63:0] _RAND_108;
  reg [63:0] _RAND_109;
  reg [63:0] _RAND_110;
  reg [63:0] _RAND_111;
  reg [63:0] _RAND_112;
  reg [63:0] _RAND_113;
  reg [63:0] _RAND_114;
  reg [63:0] _RAND_115;
  reg [63:0] _RAND_116;
  reg [63:0] _RAND_117;
  reg [63:0] _RAND_118;
  reg [63:0] _RAND_119;
  reg [63:0] _RAND_120;
  reg [63:0] _RAND_121;
  reg [63:0] _RAND_122;
  reg [63:0] _RAND_123;
  reg [63:0] _RAND_124;
  reg [63:0] _RAND_125;
  reg [63:0] _RAND_126;
  reg [63:0] _RAND_127;
  reg [63:0] _RAND_128;
  reg [63:0] _RAND_129;
  reg [63:0] _RAND_130;
  reg [63:0] _RAND_131;
  reg [63:0] _RAND_132;
  reg [63:0] _RAND_133;
  reg [63:0] _RAND_134;
  reg [63:0] _RAND_135;
  reg [63:0] _RAND_136;
  reg [63:0] _RAND_137;
  reg [63:0] _RAND_138;
  reg [63:0] _RAND_139;
  reg [63:0] _RAND_140;
  reg [63:0] _RAND_141;
  reg [63:0] _RAND_142;
  reg [63:0] _RAND_143;
  reg [63:0] _RAND_144;
  reg [63:0] _RAND_145;
  reg [63:0] _RAND_146;
  reg [63:0] _RAND_147;
  reg [63:0] _RAND_148;
  reg [63:0] _RAND_149;
  reg [63:0] _RAND_150;
  reg [63:0] _RAND_151;
  reg [63:0] _RAND_152;
  reg [63:0] _RAND_153;
  reg [63:0] _RAND_154;
  reg [63:0] _RAND_155;
  reg [63:0] _RAND_156;
  reg [63:0] _RAND_157;
  reg [63:0] _RAND_158;
  reg [63:0] _RAND_159;
  reg [63:0] _RAND_160;
  reg [63:0] _RAND_161;
  reg [63:0] _RAND_162;
  reg [63:0] _RAND_163;
  reg [63:0] _RAND_164;
  reg [63:0] _RAND_165;
  reg [63:0] _RAND_166;
  reg [63:0] _RAND_167;
  reg [63:0] _RAND_168;
  reg [63:0] _RAND_169;
  reg [63:0] _RAND_170;
  reg [63:0] _RAND_171;
  reg [63:0] _RAND_172;
  reg [63:0] _RAND_173;
  reg [63:0] _RAND_174;
  reg [63:0] _RAND_175;
  reg [63:0] _RAND_176;
  reg [63:0] _RAND_177;
  reg [63:0] _RAND_178;
  reg [63:0] _RAND_179;
  reg [63:0] _RAND_180;
  reg [63:0] _RAND_181;
  reg [63:0] _RAND_182;
  reg [63:0] _RAND_183;
  reg [63:0] _RAND_184;
  reg [63:0] _RAND_185;
  reg [63:0] _RAND_186;
  reg [63:0] _RAND_187;
  reg [63:0] _RAND_188;
  reg [63:0] _RAND_189;
  reg [63:0] _RAND_190;
  reg [63:0] _RAND_191;
  reg [63:0] _RAND_192;
  reg [63:0] _RAND_193;
  reg [63:0] _RAND_194;
  reg [63:0] _RAND_195;
  reg [63:0] _RAND_196;
  reg [63:0] _RAND_197;
  reg [63:0] _RAND_198;
  reg [63:0] _RAND_199;
  reg [63:0] _RAND_200;
  reg [63:0] _RAND_201;
  reg [63:0] _RAND_202;
  reg [63:0] _RAND_203;
  reg [63:0] _RAND_204;
  reg [63:0] _RAND_205;
  reg [63:0] _RAND_206;
  reg [63:0] _RAND_207;
  reg [63:0] _RAND_208;
  reg [63:0] _RAND_209;
  reg [63:0] _RAND_210;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
`endif // RANDOMIZE_REG_INIT
  reg [32:0] LUT_mem [0:34]; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_1_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_1_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_3_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_3_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_5_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_5_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_7_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_7_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_9_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_9_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_11_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_11_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_13_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_13_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_15_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_15_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_17_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_17_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_19_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_19_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_21_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_21_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_23_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_23_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_25_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_25_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_27_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_27_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_29_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_29_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_31_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_31_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_33_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_33_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_35_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_35_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_37_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_37_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_39_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_39_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_41_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_41_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_43_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_43_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_45_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_45_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_47_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_47_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_49_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_49_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_51_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_51_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_53_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_53_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_55_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_55_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_57_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_57_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_59_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_59_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_61_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_61_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_63_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_63_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_65_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_65_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_67_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_67_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_69_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_69_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_71_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_71_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_73_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_73_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_75_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_75_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_77_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_77_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_79_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_79_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_81_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_81_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_83_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_83_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_85_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_85_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_87_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_87_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_89_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_89_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_91_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_91_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_93_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_93_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_95_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_95_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_97_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_97_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_99_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_99_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_101_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_101_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_103_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_103_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_105_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_105_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_107_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_107_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_109_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_109_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_111_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_111_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_113_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_113_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_115_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_115_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_117_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_117_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_119_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_119_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_121_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_121_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_123_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_123_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_125_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_125_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_127_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_127_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_129_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_129_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_131_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_131_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_133_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_133_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_135_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_135_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_137_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_137_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_139_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_139_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_140_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_140_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_141_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_141_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_142_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_142_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_143_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_143_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_144_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_144_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_145_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_145_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_146_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_146_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_147_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_147_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_148_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_148_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_149_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_149_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_150_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_150_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_151_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_151_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_152_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_152_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_153_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_153_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_154_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_154_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_155_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_155_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_156_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_156_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_157_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_157_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_158_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_158_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_159_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_159_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_160_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_160_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_161_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_161_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_162_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_162_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_163_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_163_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_164_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_164_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_165_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_165_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_166_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_166_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_167_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_167_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_168_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_168_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_169_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_169_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_170_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_170_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_171_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_171_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_172_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_172_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_173_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_173_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_174_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_174_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_175_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_175_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_176_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_176_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_177_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_177_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_178_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_178_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_179_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_179_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_180_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_180_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_181_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_181_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_182_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_182_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_183_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_183_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_184_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_184_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_185_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_185_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_186_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_186_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_187_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_187_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_188_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_188_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_189_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_189_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_190_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_190_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_191_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_191_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_192_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_192_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_193_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_193_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_194_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_194_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_195_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_195_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_196_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_196_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_197_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_197_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_198_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_198_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_199_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_199_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_200_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_200_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_201_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_201_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_202_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_202_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_203_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_203_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_204_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_204_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_205_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_205_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_206_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_206_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_207_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_207_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_208_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_208_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_209_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_209_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_210_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_210_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_212_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_212_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_214_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_214_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_216_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_216_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_218_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_218_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_220_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_220_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_222_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_222_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_224_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_224_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_226_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_226_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_228_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_228_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_230_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_230_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_232_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_232_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_234_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_234_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_236_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_236_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_238_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_238_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_240_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_240_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_242_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_242_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_244_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_244_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_246_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_246_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_248_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_248_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_250_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_250_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_252_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_252_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_254_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_254_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_256_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_256_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_258_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_258_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_260_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_260_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_262_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_262_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_264_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_264_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_266_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_266_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_268_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_268_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_270_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_270_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_272_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_272_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_274_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_274_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_276_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_276_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_278_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_278_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_280_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_280_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_281_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_281_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_282_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_282_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_283_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_283_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_284_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_284_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_285_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_285_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_286_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_286_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_287_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_287_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_288_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_288_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_289_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_289_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_290_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_290_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_291_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_291_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_292_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_292_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_293_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_293_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_294_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_294_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_295_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_295_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_296_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_296_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_297_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_297_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_298_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_298_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_299_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_299_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_300_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_300_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_301_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_301_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_302_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_302_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_303_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_303_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_304_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_304_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_305_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_305_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_306_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_306_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_307_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_307_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_308_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_308_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_309_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_309_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_310_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_310_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_311_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_311_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_312_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_312_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_313_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_313_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_314_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_314_addr; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_2_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_2_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_2_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_2_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_4_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_4_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_4_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_4_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_6_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_6_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_6_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_6_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_8_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_8_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_8_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_8_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_10_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_10_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_10_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_10_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_12_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_12_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_12_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_12_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_14_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_14_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_14_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_14_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_16_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_16_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_16_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_16_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_18_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_18_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_18_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_18_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_20_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_20_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_20_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_20_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_22_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_22_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_22_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_22_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_24_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_24_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_24_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_24_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_26_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_26_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_26_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_26_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_28_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_28_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_28_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_28_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_30_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_30_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_30_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_30_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_32_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_32_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_32_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_32_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_34_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_34_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_34_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_34_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_36_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_36_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_36_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_36_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_38_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_38_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_38_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_38_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_40_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_40_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_40_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_40_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_42_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_42_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_42_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_42_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_44_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_44_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_44_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_44_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_46_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_46_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_46_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_46_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_48_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_48_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_48_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_48_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_50_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_50_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_50_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_50_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_52_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_52_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_52_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_52_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_54_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_54_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_54_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_54_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_56_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_56_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_56_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_56_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_58_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_58_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_58_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_58_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_60_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_60_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_60_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_60_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_62_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_62_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_62_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_62_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_64_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_64_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_64_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_64_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_66_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_66_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_66_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_66_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_68_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_68_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_68_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_68_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_70_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_70_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_70_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_70_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_72_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_72_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_72_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_72_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_74_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_74_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_74_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_74_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_76_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_76_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_76_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_76_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_78_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_78_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_78_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_78_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_80_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_80_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_80_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_80_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_82_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_82_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_82_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_82_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_84_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_84_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_84_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_84_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_86_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_86_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_86_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_86_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_88_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_88_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_88_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_88_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_90_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_90_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_90_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_90_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_92_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_92_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_92_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_92_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_94_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_94_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_94_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_94_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_96_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_96_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_96_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_96_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_98_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_98_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_98_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_98_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_100_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_100_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_100_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_100_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_102_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_102_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_102_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_102_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_104_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_104_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_104_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_104_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_106_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_106_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_106_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_106_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_108_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_108_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_108_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_108_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_110_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_110_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_110_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_110_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_112_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_112_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_112_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_112_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_114_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_114_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_114_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_114_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_116_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_116_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_116_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_116_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_118_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_118_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_118_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_118_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_120_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_120_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_120_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_120_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_122_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_122_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_122_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_122_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_124_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_124_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_124_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_124_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_126_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_126_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_126_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_126_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_128_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_128_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_128_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_128_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_130_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_130_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_130_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_130_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_132_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_132_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_132_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_132_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_134_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_134_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_134_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_134_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_136_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_136_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_136_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_136_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_138_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_138_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_138_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_138_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_211_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_211_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_211_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_211_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_213_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_213_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_213_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_213_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_215_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_215_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_215_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_215_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_217_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_217_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_217_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_217_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_219_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_219_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_219_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_219_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_221_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_221_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_221_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_221_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_223_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_223_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_223_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_223_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_225_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_225_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_225_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_225_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_227_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_227_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_227_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_227_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_229_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_229_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_229_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_229_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_231_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_231_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_231_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_231_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_233_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_233_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_233_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_233_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_235_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_235_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_235_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_235_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_237_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_237_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_237_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_237_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_239_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_239_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_239_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_239_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_241_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_241_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_241_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_241_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_243_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_243_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_243_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_243_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_245_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_245_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_245_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_245_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_247_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_247_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_247_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_247_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_249_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_249_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_249_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_249_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_251_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_251_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_251_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_251_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_253_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_253_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_253_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_253_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_255_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_255_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_255_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_255_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_257_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_257_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_257_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_257_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_259_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_259_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_259_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_259_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_261_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_261_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_261_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_261_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_263_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_263_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_263_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_263_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_265_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_265_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_265_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_265_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_267_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_267_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_267_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_267_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_269_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_269_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_269_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_269_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_271_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_271_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_271_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_271_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_273_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_273_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_273_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_273_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_275_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_275_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_275_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_275_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_277_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_277_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_277_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_277_en; // @[lut_35.scala 177:26]
  wire [32:0] LUT_mem_MPORT_279_data; // @[lut_35.scala 177:26]
  wire [5:0] LUT_mem_MPORT_279_addr; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_279_mask; // @[lut_35.scala 177:26]
  wire  LUT_mem_MPORT_279_en; // @[lut_35.scala 177:26]
  reg [31:0] read_stack0; // @[lut_35.scala 178:30]
  reg [31:0] read_stack1; // @[lut_35.scala 179:30]
  reg [31:0] read_stack2; // @[lut_35.scala 180:30]
  reg [31:0] read_stack3; // @[lut_35.scala 181:30]
  reg [31:0] read_stack4; // @[lut_35.scala 182:30]
  reg [31:0] read_stack5; // @[lut_35.scala 183:30]
  reg [31:0] read_stack6; // @[lut_35.scala 184:30]
  reg [31:0] read_stack7; // @[lut_35.scala 185:30]
  reg [31:0] read_stack8; // @[lut_35.scala 186:30]
  reg [31:0] read_stack9; // @[lut_35.scala 187:30]
  reg [31:0] read_stack10; // @[lut_35.scala 188:31]
  reg [31:0] read_stack11; // @[lut_35.scala 189:31]
  reg [31:0] read_stack12; // @[lut_35.scala 190:31]
  reg [31:0] read_stack13; // @[lut_35.scala 191:31]
  reg [31:0] read_stack14; // @[lut_35.scala 192:31]
  reg [31:0] read_stack15; // @[lut_35.scala 193:31]
  reg [31:0] read_stack16; // @[lut_35.scala 194:31]
  reg [31:0] read_stack17; // @[lut_35.scala 195:31]
  reg [31:0] read_stack18; // @[lut_35.scala 196:31]
  reg [31:0] read_stack19; // @[lut_35.scala 197:31]
  reg [31:0] read_stack20; // @[lut_35.scala 198:31]
  reg [31:0] read_stack21; // @[lut_35.scala 199:31]
  reg [31:0] read_stack22; // @[lut_35.scala 200:31]
  reg [31:0] read_stack23; // @[lut_35.scala 201:31]
  reg [31:0] read_stack24; // @[lut_35.scala 202:31]
  reg [31:0] read_stack25; // @[lut_35.scala 203:31]
  reg [31:0] read_stack26; // @[lut_35.scala 204:31]
  reg [31:0] read_stack27; // @[lut_35.scala 205:31]
  reg [31:0] read_stack28; // @[lut_35.scala 206:31]
  reg [31:0] read_stack29; // @[lut_35.scala 207:31]
  reg [31:0] read_stack30; // @[lut_35.scala 208:31]
  reg [31:0] read_stack31; // @[lut_35.scala 209:31]
  reg [31:0] read_stack32; // @[lut_35.scala 210:31]
  reg [31:0] read_stack33; // @[lut_35.scala 211:31]
  reg [31:0] read_stack34; // @[lut_35.scala 212:31]
  reg  push_0_1; // @[lut_35.scala 214:31]
  reg  push_1_1; // @[lut_35.scala 215:31]
  reg  push_2_1; // @[lut_35.scala 216:31]
  reg  push_3_1; // @[lut_35.scala 217:31]
  reg  push_4_1; // @[lut_35.scala 218:31]
  reg  push_5_1; // @[lut_35.scala 219:31]
  reg  push_6_1; // @[lut_35.scala 220:31]
  reg  push_7_1; // @[lut_35.scala 221:31]
  reg  push_8_1; // @[lut_35.scala 222:31]
  reg  push_9_1; // @[lut_35.scala 223:31]
  reg  push_10_1; // @[lut_35.scala 224:32]
  reg  push_11_1; // @[lut_35.scala 225:32]
  reg  push_12_1; // @[lut_35.scala 226:32]
  reg  push_13_1; // @[lut_35.scala 227:32]
  reg  push_14_1; // @[lut_35.scala 228:32]
  reg  push_15_1; // @[lut_35.scala 229:32]
  reg  push_16_1; // @[lut_35.scala 230:32]
  reg  push_17_1; // @[lut_35.scala 231:32]
  reg  push_18_1; // @[lut_35.scala 232:32]
  reg  push_19_1; // @[lut_35.scala 233:32]
  reg  push_20_1; // @[lut_35.scala 234:32]
  reg  push_21_1; // @[lut_35.scala 235:32]
  reg  push_22_1; // @[lut_35.scala 236:32]
  reg  push_23_1; // @[lut_35.scala 237:32]
  reg  push_24_1; // @[lut_35.scala 238:32]
  reg  push_25_1; // @[lut_35.scala 239:32]
  reg  push_26_1; // @[lut_35.scala 240:32]
  reg  push_27_1; // @[lut_35.scala 241:32]
  reg  push_28_1; // @[lut_35.scala 242:32]
  reg  push_29_1; // @[lut_35.scala 243:32]
  reg  push_30_1; // @[lut_35.scala 244:32]
  reg  push_31_1; // @[lut_35.scala 245:32]
  reg  push_32_1; // @[lut_35.scala 246:32]
  reg  push_33_1; // @[lut_35.scala 247:32]
  reg  push_34_1; // @[lut_35.scala 248:32]
  reg  push_1; // @[lut_35.scala 252:40]
  reg  push_valid; // @[lut_35.scala 253:41]
  reg [31:0] push_ray_id; // @[lut_35.scala 255:41]
  reg  push_valid_2; // @[lut_35.scala 295:41]
  wire [31:0] lo = LUT_mem_MPORT_1_data[31:0]; // @[lut_35.scala 301:42]
  wire [31:0] lo_1 = LUT_mem_MPORT_5_data[31:0]; // @[lut_35.scala 307:42]
  wire [31:0] lo_2 = LUT_mem_MPORT_9_data[31:0]; // @[lut_35.scala 313:42]
  wire [31:0] lo_3 = LUT_mem_MPORT_13_data[31:0]; // @[lut_35.scala 319:42]
  wire [31:0] lo_4 = LUT_mem_MPORT_17_data[31:0]; // @[lut_35.scala 325:42]
  wire [31:0] lo_5 = LUT_mem_MPORT_21_data[31:0]; // @[lut_35.scala 331:42]
  wire [31:0] lo_6 = LUT_mem_MPORT_25_data[31:0]; // @[lut_35.scala 337:42]
  wire [31:0] lo_7 = LUT_mem_MPORT_29_data[31:0]; // @[lut_35.scala 343:42]
  wire [31:0] lo_8 = LUT_mem_MPORT_33_data[31:0]; // @[lut_35.scala 349:42]
  wire [31:0] lo_9 = LUT_mem_MPORT_37_data[31:0]; // @[lut_35.scala 355:42]
  wire [31:0] lo_10 = LUT_mem_MPORT_41_data[31:0]; // @[lut_35.scala 361:44]
  wire [31:0] lo_11 = LUT_mem_MPORT_45_data[31:0]; // @[lut_35.scala 367:44]
  wire [31:0] lo_12 = LUT_mem_MPORT_49_data[31:0]; // @[lut_35.scala 373:44]
  wire [31:0] lo_13 = LUT_mem_MPORT_53_data[31:0]; // @[lut_35.scala 379:44]
  wire [31:0] lo_14 = LUT_mem_MPORT_57_data[31:0]; // @[lut_35.scala 385:44]
  wire [31:0] lo_15 = LUT_mem_MPORT_61_data[31:0]; // @[lut_35.scala 391:44]
  wire [31:0] lo_16 = LUT_mem_MPORT_65_data[31:0]; // @[lut_35.scala 397:44]
  wire [31:0] lo_17 = LUT_mem_MPORT_69_data[31:0]; // @[lut_35.scala 403:44]
  wire [31:0] lo_18 = LUT_mem_MPORT_73_data[31:0]; // @[lut_35.scala 409:44]
  wire [31:0] lo_19 = LUT_mem_MPORT_77_data[31:0]; // @[lut_35.scala 415:44]
  wire [31:0] lo_20 = LUT_mem_MPORT_81_data[31:0]; // @[lut_35.scala 421:44]
  wire [31:0] lo_21 = LUT_mem_MPORT_85_data[31:0]; // @[lut_35.scala 427:44]
  wire [31:0] lo_22 = LUT_mem_MPORT_89_data[31:0]; // @[lut_35.scala 433:44]
  wire [31:0] lo_23 = LUT_mem_MPORT_93_data[31:0]; // @[lut_35.scala 439:44]
  wire [31:0] lo_24 = LUT_mem_MPORT_97_data[31:0]; // @[lut_35.scala 445:44]
  wire [31:0] lo_25 = LUT_mem_MPORT_101_data[31:0]; // @[lut_35.scala 451:44]
  wire [31:0] lo_26 = LUT_mem_MPORT_105_data[31:0]; // @[lut_35.scala 457:44]
  wire [31:0] lo_27 = LUT_mem_MPORT_109_data[31:0]; // @[lut_35.scala 463:44]
  wire [31:0] lo_28 = LUT_mem_MPORT_113_data[31:0]; // @[lut_35.scala 469:44]
  wire [31:0] lo_29 = LUT_mem_MPORT_117_data[31:0]; // @[lut_35.scala 475:44]
  wire [31:0] lo_30 = LUT_mem_MPORT_121_data[31:0]; // @[lut_35.scala 481:44]
  wire [31:0] lo_31 = LUT_mem_MPORT_125_data[31:0]; // @[lut_35.scala 487:44]
  wire [31:0] lo_32 = LUT_mem_MPORT_129_data[31:0]; // @[lut_35.scala 493:44]
  wire [31:0] lo_33 = LUT_mem_MPORT_133_data[31:0]; // @[lut_35.scala 499:44]
  wire [31:0] lo_34 = LUT_mem_MPORT_137_data[31:0]; // @[lut_35.scala 505:44]
  wire  _T_106 = io_push & io_push_valid; // @[lut_35.scala 596:29]
  wire  _GEN_351 = io_push & io_push_valid & io_push_valid; // @[lut_35.scala 596:46 lut_35.scala 601:28 lut_35.scala 603:28]
  wire  _T_109 = push_1 & push_valid; // @[lut_35.scala 617:24]
  wire  _T_266 = read_stack0 != push_ray_id & read_stack1 != push_ray_id & read_stack2 != push_ray_id & read_stack3 !=
    push_ray_id & read_stack4 != push_ray_id & read_stack5 != push_ray_id & read_stack6 != push_ray_id & read_stack7 !=
    push_ray_id & read_stack8 != push_ray_id; // @[lut_35.scala 1948:264]
  wire  _T_280 = _T_266 & read_stack9 != push_ray_id & read_stack10 != push_ray_id & read_stack11 != push_ray_id &
    read_stack12 != push_ray_id & read_stack13 != push_ray_id & read_stack14 != push_ray_id & read_stack15 !=
    push_ray_id; // @[lut_35.scala 1949:194]
  wire  _T_292 = _T_280 & read_stack16 != push_ray_id & read_stack17 != push_ray_id & read_stack18 != push_ray_id &
    read_stack19 != push_ray_id & read_stack20 != push_ray_id & read_stack21 != push_ray_id; // @[lut_35.scala 1950:164]
  wire  _T_304 = _T_292 & read_stack22 != push_ray_id & read_stack23 != push_ray_id & read_stack24 != push_ray_id &
    read_stack25 != push_ray_id & read_stack26 != push_ray_id & read_stack27 != push_ray_id; // @[lut_35.scala 1951:165]
  wire  _T_312 = _T_304 & read_stack28 != push_ray_id & read_stack29 != push_ray_id & read_stack30 != push_ray_id &
    read_stack31 != push_ray_id; // @[lut_35.scala 1952:102]
  wire  _T_320 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid; // @[lut_35.scala 1953:102]
  wire  _T_328 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32]; // @[lut_35.scala 1954:78]
  wire  _T_337 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32]; // @[lut_35.scala 1994:78]
  wire  _T_346 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32]; // @[lut_35.scala 2034:78]
  wire  _T_355 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32]; // @[lut_35.scala 2074:78]
  wire  _T_364 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32]; // @[lut_35.scala 2114:78]
  wire  _T_373 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32]; // @[lut_35.scala 2154:78]
  wire  _T_382 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32]; // @[lut_35.scala 2194:78]
  wire  _T_391 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32]; // @[lut_35.scala 2234:78]
  wire  _T_400 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32]; // @[lut_35.scala 2274:78]
  wire  _T_409 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32]; // @[lut_35.scala 2314:78]
  wire  _T_418 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32]; // @[lut_35.scala 2354:80]
  wire  _T_427 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32]; // @[lut_35.scala 2394:80]
  wire  _T_436 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32]; // @[lut_35.scala 2434:80]
  wire  _T_445 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32]; // @[lut_35.scala 2474:80]
  wire  _T_454 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_238_data[32]; // @[lut_35.scala 2514:80]
  wire  _T_463 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_240_data[32]; // @[lut_35.scala 2554:80]
  wire  _T_472 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_242_data[32]; // @[lut_35.scala 2594:80]
  wire  _T_481 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_244_data[32]; // @[lut_35.scala 2634:80]
  wire  _T_490 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_246_data[32]; // @[lut_35.scala 2674:80]
  wire  _T_499 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_248_data[32]; // @[lut_35.scala 2714:80]
  wire  _T_508 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_250_data[32]; // @[lut_35.scala 2754:80]
  wire  _T_517 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_252_data[32]; // @[lut_35.scala 2794:80]
  wire  _T_526 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_254_data[32]; // @[lut_35.scala 2834:80]
  wire  _T_535 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_256_data[32]; // @[lut_35.scala 2874:80]
  wire  _T_544 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_258_data[32]; // @[lut_35.scala 2915:80]
  wire  _T_553 = io_empty_25 & push_valid & ~push_25_1 & ~LUT_mem_MPORT_260_data[32]; // @[lut_35.scala 2955:82]
  wire  _T_562 = io_empty_26 & push_valid & ~push_26_1 & ~LUT_mem_MPORT_262_data[32]; // @[lut_35.scala 2995:82]
  wire  _T_571 = io_empty_27 & push_valid & ~push_27_1 & ~LUT_mem_MPORT_264_data[32]; // @[lut_35.scala 3035:81]
  wire  _T_580 = io_empty_28 & push_valid & ~push_28_1 & ~LUT_mem_MPORT_266_data[32]; // @[lut_35.scala 3075:81]
  wire  _T_589 = io_empty_29 & push_valid & ~push_29_1 & ~LUT_mem_MPORT_268_data[32]; // @[lut_35.scala 3115:81]
  wire  _T_598 = io_empty_30 & push_valid & ~push_30_1 & ~LUT_mem_MPORT_270_data[32]; // @[lut_35.scala 3155:81]
  wire  _T_607 = io_empty_31 & push_valid & ~push_31_1 & ~LUT_mem_MPORT_272_data[32]; // @[lut_35.scala 3195:81]
  wire  _T_616 = io_empty_32 & push_valid & ~push_32_1 & ~LUT_mem_MPORT_274_data[32]; // @[lut_35.scala 3235:81]
  wire  _T_625 = io_empty_33 & push_valid & ~push_33_1 & ~LUT_mem_MPORT_276_data[32]; // @[lut_35.scala 3275:80]
  wire  _T_634 = io_empty_34 & push_valid & ~push_34_1 & ~LUT_mem_MPORT_278_data[32]; // @[lut_35.scala 3315:80]
  wire  _GEN_366 = io_empty_33 & push_valid & ~push_33_1 & ~LUT_mem_MPORT_276_data[32] ? 1'h0 : _T_634; // @[lut_35.scala 3275:105 lut_35.scala 3312:43]
  wire  _GEN_367 = io_empty_33 & push_valid & ~push_33_1 & ~LUT_mem_MPORT_276_data[32] | _T_634; // @[lut_35.scala 3275:105 lut_35.scala 3313:38]
  wire  _GEN_371 = io_empty_33 & push_valid & ~push_33_1 & ~LUT_mem_MPORT_276_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 3275:105 lut_35.scala 177:26 lut_35.scala 3315:89]
  wire  _GEN_383 = io_empty_32 & push_valid & ~push_32_1 & ~LUT_mem_MPORT_274_data[32] ? 1'h0 : _T_625; // @[lut_35.scala 3235:106 lut_35.scala 3271:43]
  wire  _GEN_384 = io_empty_32 & push_valid & ~push_32_1 & ~LUT_mem_MPORT_274_data[32] ? 1'h0 : _GEN_366; // @[lut_35.scala 3235:106 lut_35.scala 3272:43]
  wire  _GEN_385 = io_empty_32 & push_valid & ~push_32_1 & ~LUT_mem_MPORT_274_data[32] | _GEN_367; // @[lut_35.scala 3235:106 lut_35.scala 3273:38]
  wire  _GEN_389 = io_empty_32 & push_valid & ~push_32_1 & ~LUT_mem_MPORT_274_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 3235:106 lut_35.scala 177:26 lut_35.scala 3275:89]
  wire  _GEN_397 = io_empty_32 & push_valid & ~push_32_1 & ~LUT_mem_MPORT_274_data[32] ? 1'h0 : _GEN_371; // @[lut_35.scala 3235:106 lut_35.scala 177:26]
  wire  _GEN_409 = io_empty_31 & push_valid & ~push_31_1 & ~LUT_mem_MPORT_272_data[32] ? 1'h0 : _T_616; // @[lut_35.scala 3195:106 lut_35.scala 3230:43]
  wire  _GEN_410 = io_empty_31 & push_valid & ~push_31_1 & ~LUT_mem_MPORT_272_data[32] ? 1'h0 : _GEN_383; // @[lut_35.scala 3195:106 lut_35.scala 3231:43]
  wire  _GEN_411 = io_empty_31 & push_valid & ~push_31_1 & ~LUT_mem_MPORT_272_data[32] ? 1'h0 : _GEN_384; // @[lut_35.scala 3195:106 lut_35.scala 3232:43]
  wire  _GEN_412 = io_empty_31 & push_valid & ~push_31_1 & ~LUT_mem_MPORT_272_data[32] | _GEN_385; // @[lut_35.scala 3195:106 lut_35.scala 3233:38]
  wire  _GEN_416 = io_empty_31 & push_valid & ~push_31_1 & ~LUT_mem_MPORT_272_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 3195:106 lut_35.scala 177:26 lut_35.scala 3235:90]
  wire  _GEN_424 = io_empty_31 & push_valid & ~push_31_1 & ~LUT_mem_MPORT_272_data[32] ? 1'h0 : _GEN_389; // @[lut_35.scala 3195:106 lut_35.scala 177:26]
  wire  _GEN_432 = io_empty_31 & push_valid & ~push_31_1 & ~LUT_mem_MPORT_272_data[32] ? 1'h0 : _GEN_397; // @[lut_35.scala 3195:106 lut_35.scala 177:26]
  wire  _GEN_444 = io_empty_30 & push_valid & ~push_30_1 & ~LUT_mem_MPORT_270_data[32] ? 1'h0 : _T_607; // @[lut_35.scala 3155:106 lut_35.scala 3189:43]
  wire  _GEN_445 = io_empty_30 & push_valid & ~push_30_1 & ~LUT_mem_MPORT_270_data[32] ? 1'h0 : _GEN_409; // @[lut_35.scala 3155:106 lut_35.scala 3190:43]
  wire  _GEN_446 = io_empty_30 & push_valid & ~push_30_1 & ~LUT_mem_MPORT_270_data[32] ? 1'h0 : _GEN_410; // @[lut_35.scala 3155:106 lut_35.scala 3191:43]
  wire  _GEN_447 = io_empty_30 & push_valid & ~push_30_1 & ~LUT_mem_MPORT_270_data[32] ? 1'h0 : _GEN_411; // @[lut_35.scala 3155:106 lut_35.scala 3192:43]
  wire  _GEN_448 = io_empty_30 & push_valid & ~push_30_1 & ~LUT_mem_MPORT_270_data[32] | _GEN_412; // @[lut_35.scala 3155:106 lut_35.scala 3193:38]
  wire  _GEN_452 = io_empty_30 & push_valid & ~push_30_1 & ~LUT_mem_MPORT_270_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 3155:106 lut_35.scala 177:26 lut_35.scala 3195:90]
  wire  _GEN_460 = io_empty_30 & push_valid & ~push_30_1 & ~LUT_mem_MPORT_270_data[32] ? 1'h0 : _GEN_416; // @[lut_35.scala 3155:106 lut_35.scala 177:26]
  wire  _GEN_468 = io_empty_30 & push_valid & ~push_30_1 & ~LUT_mem_MPORT_270_data[32] ? 1'h0 : _GEN_424; // @[lut_35.scala 3155:106 lut_35.scala 177:26]
  wire  _GEN_476 = io_empty_30 & push_valid & ~push_30_1 & ~LUT_mem_MPORT_270_data[32] ? 1'h0 : _GEN_432; // @[lut_35.scala 3155:106 lut_35.scala 177:26]
  wire  _GEN_488 = io_empty_29 & push_valid & ~push_29_1 & ~LUT_mem_MPORT_268_data[32] ? 1'h0 : _T_598; // @[lut_35.scala 3115:106 lut_35.scala 3148:43]
  wire  _GEN_489 = io_empty_29 & push_valid & ~push_29_1 & ~LUT_mem_MPORT_268_data[32] ? 1'h0 : _GEN_444; // @[lut_35.scala 3115:106 lut_35.scala 3149:43]
  wire  _GEN_490 = io_empty_29 & push_valid & ~push_29_1 & ~LUT_mem_MPORT_268_data[32] ? 1'h0 : _GEN_445; // @[lut_35.scala 3115:106 lut_35.scala 3150:43]
  wire  _GEN_491 = io_empty_29 & push_valid & ~push_29_1 & ~LUT_mem_MPORT_268_data[32] ? 1'h0 : _GEN_446; // @[lut_35.scala 3115:106 lut_35.scala 3151:43]
  wire  _GEN_492 = io_empty_29 & push_valid & ~push_29_1 & ~LUT_mem_MPORT_268_data[32] ? 1'h0 : _GEN_447; // @[lut_35.scala 3115:106 lut_35.scala 3152:43]
  wire  _GEN_493 = io_empty_29 & push_valid & ~push_29_1 & ~LUT_mem_MPORT_268_data[32] | _GEN_448; // @[lut_35.scala 3115:106 lut_35.scala 3153:38]
  wire  _GEN_497 = io_empty_29 & push_valid & ~push_29_1 & ~LUT_mem_MPORT_268_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 3115:106 lut_35.scala 177:26 lut_35.scala 3155:90]
  wire  _GEN_505 = io_empty_29 & push_valid & ~push_29_1 & ~LUT_mem_MPORT_268_data[32] ? 1'h0 : _GEN_452; // @[lut_35.scala 3115:106 lut_35.scala 177:26]
  wire  _GEN_513 = io_empty_29 & push_valid & ~push_29_1 & ~LUT_mem_MPORT_268_data[32] ? 1'h0 : _GEN_460; // @[lut_35.scala 3115:106 lut_35.scala 177:26]
  wire  _GEN_521 = io_empty_29 & push_valid & ~push_29_1 & ~LUT_mem_MPORT_268_data[32] ? 1'h0 : _GEN_468; // @[lut_35.scala 3115:106 lut_35.scala 177:26]
  wire  _GEN_529 = io_empty_29 & push_valid & ~push_29_1 & ~LUT_mem_MPORT_268_data[32] ? 1'h0 : _GEN_476; // @[lut_35.scala 3115:106 lut_35.scala 177:26]
  wire  _GEN_541 = io_empty_28 & push_valid & ~push_28_1 & ~LUT_mem_MPORT_266_data[32] ? 1'h0 : _T_589; // @[lut_35.scala 3075:106 lut_35.scala 3107:43]
  wire  _GEN_542 = io_empty_28 & push_valid & ~push_28_1 & ~LUT_mem_MPORT_266_data[32] ? 1'h0 : _GEN_488; // @[lut_35.scala 3075:106 lut_35.scala 3108:43]
  wire  _GEN_543 = io_empty_28 & push_valid & ~push_28_1 & ~LUT_mem_MPORT_266_data[32] ? 1'h0 : _GEN_489; // @[lut_35.scala 3075:106 lut_35.scala 3109:43]
  wire  _GEN_544 = io_empty_28 & push_valid & ~push_28_1 & ~LUT_mem_MPORT_266_data[32] ? 1'h0 : _GEN_490; // @[lut_35.scala 3075:106 lut_35.scala 3110:43]
  wire  _GEN_545 = io_empty_28 & push_valid & ~push_28_1 & ~LUT_mem_MPORT_266_data[32] ? 1'h0 : _GEN_491; // @[lut_35.scala 3075:106 lut_35.scala 3111:43]
  wire  _GEN_546 = io_empty_28 & push_valid & ~push_28_1 & ~LUT_mem_MPORT_266_data[32] ? 1'h0 : _GEN_492; // @[lut_35.scala 3075:106 lut_35.scala 3112:43]
  wire  _GEN_547 = io_empty_28 & push_valid & ~push_28_1 & ~LUT_mem_MPORT_266_data[32] | _GEN_493; // @[lut_35.scala 3075:106 lut_35.scala 3113:38]
  wire  _GEN_551 = io_empty_28 & push_valid & ~push_28_1 & ~LUT_mem_MPORT_266_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 3075:106 lut_35.scala 177:26 lut_35.scala 3115:90]
  wire  _GEN_559 = io_empty_28 & push_valid & ~push_28_1 & ~LUT_mem_MPORT_266_data[32] ? 1'h0 : _GEN_497; // @[lut_35.scala 3075:106 lut_35.scala 177:26]
  wire  _GEN_567 = io_empty_28 & push_valid & ~push_28_1 & ~LUT_mem_MPORT_266_data[32] ? 1'h0 : _GEN_505; // @[lut_35.scala 3075:106 lut_35.scala 177:26]
  wire  _GEN_575 = io_empty_28 & push_valid & ~push_28_1 & ~LUT_mem_MPORT_266_data[32] ? 1'h0 : _GEN_513; // @[lut_35.scala 3075:106 lut_35.scala 177:26]
  wire  _GEN_583 = io_empty_28 & push_valid & ~push_28_1 & ~LUT_mem_MPORT_266_data[32] ? 1'h0 : _GEN_521; // @[lut_35.scala 3075:106 lut_35.scala 177:26]
  wire  _GEN_591 = io_empty_28 & push_valid & ~push_28_1 & ~LUT_mem_MPORT_266_data[32] ? 1'h0 : _GEN_529; // @[lut_35.scala 3075:106 lut_35.scala 177:26]
  wire  _GEN_603 = io_empty_27 & push_valid & ~push_27_1 & ~LUT_mem_MPORT_264_data[32] ? 1'h0 : _T_580; // @[lut_35.scala 3035:106 lut_35.scala 3066:43]
  wire  _GEN_604 = io_empty_27 & push_valid & ~push_27_1 & ~LUT_mem_MPORT_264_data[32] ? 1'h0 : _GEN_541; // @[lut_35.scala 3035:106 lut_35.scala 3067:43]
  wire  _GEN_605 = io_empty_27 & push_valid & ~push_27_1 & ~LUT_mem_MPORT_264_data[32] ? 1'h0 : _GEN_542; // @[lut_35.scala 3035:106 lut_35.scala 3068:43]
  wire  _GEN_606 = io_empty_27 & push_valid & ~push_27_1 & ~LUT_mem_MPORT_264_data[32] ? 1'h0 : _GEN_543; // @[lut_35.scala 3035:106 lut_35.scala 3069:43]
  wire  _GEN_607 = io_empty_27 & push_valid & ~push_27_1 & ~LUT_mem_MPORT_264_data[32] ? 1'h0 : _GEN_544; // @[lut_35.scala 3035:106 lut_35.scala 3070:43]
  wire  _GEN_608 = io_empty_27 & push_valid & ~push_27_1 & ~LUT_mem_MPORT_264_data[32] ? 1'h0 : _GEN_545; // @[lut_35.scala 3035:106 lut_35.scala 3071:43]
  wire  _GEN_609 = io_empty_27 & push_valid & ~push_27_1 & ~LUT_mem_MPORT_264_data[32] ? 1'h0 : _GEN_546; // @[lut_35.scala 3035:106 lut_35.scala 3072:43]
  wire  _GEN_610 = io_empty_27 & push_valid & ~push_27_1 & ~LUT_mem_MPORT_264_data[32] | _GEN_547; // @[lut_35.scala 3035:106 lut_35.scala 3073:38]
  wire  _GEN_614 = io_empty_27 & push_valid & ~push_27_1 & ~LUT_mem_MPORT_264_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 3035:106 lut_35.scala 177:26 lut_35.scala 3075:90]
  wire  _GEN_622 = io_empty_27 & push_valid & ~push_27_1 & ~LUT_mem_MPORT_264_data[32] ? 1'h0 : _GEN_551; // @[lut_35.scala 3035:106 lut_35.scala 177:26]
  wire  _GEN_630 = io_empty_27 & push_valid & ~push_27_1 & ~LUT_mem_MPORT_264_data[32] ? 1'h0 : _GEN_559; // @[lut_35.scala 3035:106 lut_35.scala 177:26]
  wire  _GEN_638 = io_empty_27 & push_valid & ~push_27_1 & ~LUT_mem_MPORT_264_data[32] ? 1'h0 : _GEN_567; // @[lut_35.scala 3035:106 lut_35.scala 177:26]
  wire  _GEN_646 = io_empty_27 & push_valid & ~push_27_1 & ~LUT_mem_MPORT_264_data[32] ? 1'h0 : _GEN_575; // @[lut_35.scala 3035:106 lut_35.scala 177:26]
  wire  _GEN_654 = io_empty_27 & push_valid & ~push_27_1 & ~LUT_mem_MPORT_264_data[32] ? 1'h0 : _GEN_583; // @[lut_35.scala 3035:106 lut_35.scala 177:26]
  wire  _GEN_662 = io_empty_27 & push_valid & ~push_27_1 & ~LUT_mem_MPORT_264_data[32] ? 1'h0 : _GEN_591; // @[lut_35.scala 3035:106 lut_35.scala 177:26]
  wire  _GEN_674 = io_empty_26 & push_valid & ~push_26_1 & ~LUT_mem_MPORT_262_data[32] ? 1'h0 : _T_571; // @[lut_35.scala 2995:107 lut_35.scala 3025:43]
  wire  _GEN_675 = io_empty_26 & push_valid & ~push_26_1 & ~LUT_mem_MPORT_262_data[32] ? 1'h0 : _GEN_603; // @[lut_35.scala 2995:107 lut_35.scala 3026:43]
  wire  _GEN_676 = io_empty_26 & push_valid & ~push_26_1 & ~LUT_mem_MPORT_262_data[32] ? 1'h0 : _GEN_604; // @[lut_35.scala 2995:107 lut_35.scala 3027:43]
  wire  _GEN_677 = io_empty_26 & push_valid & ~push_26_1 & ~LUT_mem_MPORT_262_data[32] ? 1'h0 : _GEN_605; // @[lut_35.scala 2995:107 lut_35.scala 3028:43]
  wire  _GEN_678 = io_empty_26 & push_valid & ~push_26_1 & ~LUT_mem_MPORT_262_data[32] ? 1'h0 : _GEN_606; // @[lut_35.scala 2995:107 lut_35.scala 3029:43]
  wire  _GEN_679 = io_empty_26 & push_valid & ~push_26_1 & ~LUT_mem_MPORT_262_data[32] ? 1'h0 : _GEN_607; // @[lut_35.scala 2995:107 lut_35.scala 3030:43]
  wire  _GEN_680 = io_empty_26 & push_valid & ~push_26_1 & ~LUT_mem_MPORT_262_data[32] ? 1'h0 : _GEN_608; // @[lut_35.scala 2995:107 lut_35.scala 3031:43]
  wire  _GEN_681 = io_empty_26 & push_valid & ~push_26_1 & ~LUT_mem_MPORT_262_data[32] ? 1'h0 : _GEN_609; // @[lut_35.scala 2995:107 lut_35.scala 3032:43]
  wire  _GEN_682 = io_empty_26 & push_valid & ~push_26_1 & ~LUT_mem_MPORT_262_data[32] | _GEN_610; // @[lut_35.scala 2995:107 lut_35.scala 3033:38]
  wire  _GEN_686 = io_empty_26 & push_valid & ~push_26_1 & ~LUT_mem_MPORT_262_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2995:107 lut_35.scala 177:26 lut_35.scala 3035:90]
  wire  _GEN_694 = io_empty_26 & push_valid & ~push_26_1 & ~LUT_mem_MPORT_262_data[32] ? 1'h0 : _GEN_614; // @[lut_35.scala 2995:107 lut_35.scala 177:26]
  wire  _GEN_702 = io_empty_26 & push_valid & ~push_26_1 & ~LUT_mem_MPORT_262_data[32] ? 1'h0 : _GEN_622; // @[lut_35.scala 2995:107 lut_35.scala 177:26]
  wire  _GEN_710 = io_empty_26 & push_valid & ~push_26_1 & ~LUT_mem_MPORT_262_data[32] ? 1'h0 : _GEN_630; // @[lut_35.scala 2995:107 lut_35.scala 177:26]
  wire  _GEN_718 = io_empty_26 & push_valid & ~push_26_1 & ~LUT_mem_MPORT_262_data[32] ? 1'h0 : _GEN_638; // @[lut_35.scala 2995:107 lut_35.scala 177:26]
  wire  _GEN_726 = io_empty_26 & push_valid & ~push_26_1 & ~LUT_mem_MPORT_262_data[32] ? 1'h0 : _GEN_646; // @[lut_35.scala 2995:107 lut_35.scala 177:26]
  wire  _GEN_734 = io_empty_26 & push_valid & ~push_26_1 & ~LUT_mem_MPORT_262_data[32] ? 1'h0 : _GEN_654; // @[lut_35.scala 2995:107 lut_35.scala 177:26]
  wire  _GEN_742 = io_empty_26 & push_valid & ~push_26_1 & ~LUT_mem_MPORT_262_data[32] ? 1'h0 : _GEN_662; // @[lut_35.scala 2995:107 lut_35.scala 177:26]
  wire  _GEN_754 = io_empty_25 & push_valid & ~push_25_1 & ~LUT_mem_MPORT_260_data[32] ? 1'h0 : _T_562; // @[lut_35.scala 2955:107 lut_35.scala 2984:43]
  wire  _GEN_755 = io_empty_25 & push_valid & ~push_25_1 & ~LUT_mem_MPORT_260_data[32] ? 1'h0 : _GEN_674; // @[lut_35.scala 2955:107 lut_35.scala 2985:43]
  wire  _GEN_756 = io_empty_25 & push_valid & ~push_25_1 & ~LUT_mem_MPORT_260_data[32] ? 1'h0 : _GEN_675; // @[lut_35.scala 2955:107 lut_35.scala 2986:43]
  wire  _GEN_757 = io_empty_25 & push_valid & ~push_25_1 & ~LUT_mem_MPORT_260_data[32] ? 1'h0 : _GEN_676; // @[lut_35.scala 2955:107 lut_35.scala 2987:43]
  wire  _GEN_758 = io_empty_25 & push_valid & ~push_25_1 & ~LUT_mem_MPORT_260_data[32] ? 1'h0 : _GEN_677; // @[lut_35.scala 2955:107 lut_35.scala 2988:43]
  wire  _GEN_759 = io_empty_25 & push_valid & ~push_25_1 & ~LUT_mem_MPORT_260_data[32] ? 1'h0 : _GEN_678; // @[lut_35.scala 2955:107 lut_35.scala 2989:43]
  wire  _GEN_760 = io_empty_25 & push_valid & ~push_25_1 & ~LUT_mem_MPORT_260_data[32] ? 1'h0 : _GEN_679; // @[lut_35.scala 2955:107 lut_35.scala 2990:43]
  wire  _GEN_761 = io_empty_25 & push_valid & ~push_25_1 & ~LUT_mem_MPORT_260_data[32] ? 1'h0 : _GEN_680; // @[lut_35.scala 2955:107 lut_35.scala 2991:43]
  wire  _GEN_762 = io_empty_25 & push_valid & ~push_25_1 & ~LUT_mem_MPORT_260_data[32] ? 1'h0 : _GEN_681; // @[lut_35.scala 2955:107 lut_35.scala 2992:43]
  wire  _GEN_763 = io_empty_25 & push_valid & ~push_25_1 & ~LUT_mem_MPORT_260_data[32] | _GEN_682; // @[lut_35.scala 2955:107 lut_35.scala 2993:38]
  wire  _GEN_767 = io_empty_25 & push_valid & ~push_25_1 & ~LUT_mem_MPORT_260_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2955:107 lut_35.scala 177:26 lut_35.scala 2995:91]
  wire  _GEN_775 = io_empty_25 & push_valid & ~push_25_1 & ~LUT_mem_MPORT_260_data[32] ? 1'h0 : _GEN_686; // @[lut_35.scala 2955:107 lut_35.scala 177:26]
  wire  _GEN_783 = io_empty_25 & push_valid & ~push_25_1 & ~LUT_mem_MPORT_260_data[32] ? 1'h0 : _GEN_694; // @[lut_35.scala 2955:107 lut_35.scala 177:26]
  wire  _GEN_791 = io_empty_25 & push_valid & ~push_25_1 & ~LUT_mem_MPORT_260_data[32] ? 1'h0 : _GEN_702; // @[lut_35.scala 2955:107 lut_35.scala 177:26]
  wire  _GEN_799 = io_empty_25 & push_valid & ~push_25_1 & ~LUT_mem_MPORT_260_data[32] ? 1'h0 : _GEN_710; // @[lut_35.scala 2955:107 lut_35.scala 177:26]
  wire  _GEN_807 = io_empty_25 & push_valid & ~push_25_1 & ~LUT_mem_MPORT_260_data[32] ? 1'h0 : _GEN_718; // @[lut_35.scala 2955:107 lut_35.scala 177:26]
  wire  _GEN_815 = io_empty_25 & push_valid & ~push_25_1 & ~LUT_mem_MPORT_260_data[32] ? 1'h0 : _GEN_726; // @[lut_35.scala 2955:107 lut_35.scala 177:26]
  wire  _GEN_823 = io_empty_25 & push_valid & ~push_25_1 & ~LUT_mem_MPORT_260_data[32] ? 1'h0 : _GEN_734; // @[lut_35.scala 2955:107 lut_35.scala 177:26]
  wire  _GEN_831 = io_empty_25 & push_valid & ~push_25_1 & ~LUT_mem_MPORT_260_data[32] ? 1'h0 : _GEN_742; // @[lut_35.scala 2955:107 lut_35.scala 177:26]
  wire  _GEN_843 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_258_data[32] ? 1'h0 : _T_553; // @[lut_35.scala 2915:105 lut_35.scala 2943:43]
  wire  _GEN_844 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_258_data[32] ? 1'h0 : _GEN_754; // @[lut_35.scala 2915:105 lut_35.scala 2944:43]
  wire  _GEN_845 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_258_data[32] ? 1'h0 : _GEN_755; // @[lut_35.scala 2915:105 lut_35.scala 2945:43]
  wire  _GEN_846 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_258_data[32] ? 1'h0 : _GEN_756; // @[lut_35.scala 2915:105 lut_35.scala 2946:43]
  wire  _GEN_847 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_258_data[32] ? 1'h0 : _GEN_757; // @[lut_35.scala 2915:105 lut_35.scala 2947:43]
  wire  _GEN_848 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_258_data[32] ? 1'h0 : _GEN_758; // @[lut_35.scala 2915:105 lut_35.scala 2948:43]
  wire  _GEN_849 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_258_data[32] ? 1'h0 : _GEN_759; // @[lut_35.scala 2915:105 lut_35.scala 2949:43]
  wire  _GEN_850 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_258_data[32] ? 1'h0 : _GEN_760; // @[lut_35.scala 2915:105 lut_35.scala 2950:43]
  wire  _GEN_851 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_258_data[32] ? 1'h0 : _GEN_761; // @[lut_35.scala 2915:105 lut_35.scala 2951:43]
  wire  _GEN_852 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_258_data[32] ? 1'h0 : _GEN_762; // @[lut_35.scala 2915:105 lut_35.scala 2952:43]
  wire  _GEN_853 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_258_data[32] | _GEN_763; // @[lut_35.scala 2915:105 lut_35.scala 2953:38]
  wire  _GEN_857 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_258_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2915:105 lut_35.scala 177:26 lut_35.scala 2955:91]
  wire  _GEN_865 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_258_data[32] ? 1'h0 : _GEN_767; // @[lut_35.scala 2915:105 lut_35.scala 177:26]
  wire  _GEN_873 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_258_data[32] ? 1'h0 : _GEN_775; // @[lut_35.scala 2915:105 lut_35.scala 177:26]
  wire  _GEN_881 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_258_data[32] ? 1'h0 : _GEN_783; // @[lut_35.scala 2915:105 lut_35.scala 177:26]
  wire  _GEN_889 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_258_data[32] ? 1'h0 : _GEN_791; // @[lut_35.scala 2915:105 lut_35.scala 177:26]
  wire  _GEN_897 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_258_data[32] ? 1'h0 : _GEN_799; // @[lut_35.scala 2915:105 lut_35.scala 177:26]
  wire  _GEN_905 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_258_data[32] ? 1'h0 : _GEN_807; // @[lut_35.scala 2915:105 lut_35.scala 177:26]
  wire  _GEN_913 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_258_data[32] ? 1'h0 : _GEN_815; // @[lut_35.scala 2915:105 lut_35.scala 177:26]
  wire  _GEN_921 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_258_data[32] ? 1'h0 : _GEN_823; // @[lut_35.scala 2915:105 lut_35.scala 177:26]
  wire  _GEN_929 = io_empty_24 & push_valid & ~push_24_1 & ~LUT_mem_MPORT_258_data[32] ? 1'h0 : _GEN_831; // @[lut_35.scala 2915:105 lut_35.scala 177:26]
  wire  _GEN_941 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_256_data[32] ? 1'h0 : _T_544; // @[lut_35.scala 2874:105 lut_35.scala 2901:43]
  wire  _GEN_942 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_256_data[32] ? 1'h0 : _GEN_843; // @[lut_35.scala 2874:105 lut_35.scala 2902:43]
  wire  _GEN_943 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_256_data[32] ? 1'h0 : _GEN_844; // @[lut_35.scala 2874:105 lut_35.scala 2903:43]
  wire  _GEN_944 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_256_data[32] ? 1'h0 : _GEN_845; // @[lut_35.scala 2874:105 lut_35.scala 2904:43]
  wire  _GEN_945 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_256_data[32] ? 1'h0 : _GEN_846; // @[lut_35.scala 2874:105 lut_35.scala 2905:43]
  wire  _GEN_946 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_256_data[32] ? 1'h0 : _GEN_847; // @[lut_35.scala 2874:105 lut_35.scala 2906:43]
  wire  _GEN_947 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_256_data[32] ? 1'h0 : _GEN_848; // @[lut_35.scala 2874:105 lut_35.scala 2907:43]
  wire  _GEN_948 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_256_data[32] ? 1'h0 : _GEN_849; // @[lut_35.scala 2874:105 lut_35.scala 2908:43]
  wire  _GEN_949 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_256_data[32] ? 1'h0 : _GEN_850; // @[lut_35.scala 2874:105 lut_35.scala 2909:43]
  wire  _GEN_950 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_256_data[32] ? 1'h0 : _GEN_851; // @[lut_35.scala 2874:105 lut_35.scala 2910:43]
  wire  _GEN_951 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_256_data[32] ? 1'h0 : _GEN_852; // @[lut_35.scala 2874:105 lut_35.scala 2911:43]
  wire  _GEN_952 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_256_data[32] | _GEN_853; // @[lut_35.scala 2874:105 lut_35.scala 2912:38]
  wire  _GEN_956 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_256_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2874:105 lut_35.scala 177:26 lut_35.scala 2915:89]
  wire  _GEN_964 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_256_data[32] ? 1'h0 : _GEN_857; // @[lut_35.scala 2874:105 lut_35.scala 177:26]
  wire  _GEN_972 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_256_data[32] ? 1'h0 : _GEN_865; // @[lut_35.scala 2874:105 lut_35.scala 177:26]
  wire  _GEN_980 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_256_data[32] ? 1'h0 : _GEN_873; // @[lut_35.scala 2874:105 lut_35.scala 177:26]
  wire  _GEN_988 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_256_data[32] ? 1'h0 : _GEN_881; // @[lut_35.scala 2874:105 lut_35.scala 177:26]
  wire  _GEN_996 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_256_data[32] ? 1'h0 : _GEN_889; // @[lut_35.scala 2874:105 lut_35.scala 177:26]
  wire  _GEN_1004 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_256_data[32] ? 1'h0 : _GEN_897; // @[lut_35.scala 2874:105 lut_35.scala 177:26]
  wire  _GEN_1012 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_256_data[32] ? 1'h0 : _GEN_905; // @[lut_35.scala 2874:105 lut_35.scala 177:26]
  wire  _GEN_1020 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_256_data[32] ? 1'h0 : _GEN_913; // @[lut_35.scala 2874:105 lut_35.scala 177:26]
  wire  _GEN_1028 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_256_data[32] ? 1'h0 : _GEN_921; // @[lut_35.scala 2874:105 lut_35.scala 177:26]
  wire  _GEN_1036 = io_empty_23 & push_valid & ~push_23_1 & ~LUT_mem_MPORT_256_data[32] ? 1'h0 : _GEN_929; // @[lut_35.scala 2874:105 lut_35.scala 177:26]
  wire  _GEN_1048 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_254_data[32] ? 1'h0 : _T_535; // @[lut_35.scala 2834:105 lut_35.scala 2860:43]
  wire  _GEN_1049 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_254_data[32] ? 1'h0 : _GEN_941; // @[lut_35.scala 2834:105 lut_35.scala 2861:43]
  wire  _GEN_1050 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_254_data[32] ? 1'h0 : _GEN_942; // @[lut_35.scala 2834:105 lut_35.scala 2862:43]
  wire  _GEN_1051 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_254_data[32] ? 1'h0 : _GEN_943; // @[lut_35.scala 2834:105 lut_35.scala 2863:43]
  wire  _GEN_1052 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_254_data[32] ? 1'h0 : _GEN_944; // @[lut_35.scala 2834:105 lut_35.scala 2864:43]
  wire  _GEN_1053 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_254_data[32] ? 1'h0 : _GEN_945; // @[lut_35.scala 2834:105 lut_35.scala 2865:43]
  wire  _GEN_1054 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_254_data[32] ? 1'h0 : _GEN_946; // @[lut_35.scala 2834:105 lut_35.scala 2866:43]
  wire  _GEN_1055 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_254_data[32] ? 1'h0 : _GEN_947; // @[lut_35.scala 2834:105 lut_35.scala 2867:43]
  wire  _GEN_1056 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_254_data[32] ? 1'h0 : _GEN_948; // @[lut_35.scala 2834:105 lut_35.scala 2868:43]
  wire  _GEN_1057 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_254_data[32] ? 1'h0 : _GEN_949; // @[lut_35.scala 2834:105 lut_35.scala 2869:43]
  wire  _GEN_1058 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_254_data[32] ? 1'h0 : _GEN_950; // @[lut_35.scala 2834:105 lut_35.scala 2870:43]
  wire  _GEN_1059 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_254_data[32] ? 1'h0 : _GEN_951; // @[lut_35.scala 2834:105 lut_35.scala 2871:43]
  wire  _GEN_1060 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_254_data[32] | _GEN_952; // @[lut_35.scala 2834:105 lut_35.scala 2872:38]
  wire  _GEN_1064 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_254_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2834:105 lut_35.scala 177:26 lut_35.scala 2874:89]
  wire  _GEN_1072 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_254_data[32] ? 1'h0 : _GEN_956; // @[lut_35.scala 2834:105 lut_35.scala 177:26]
  wire  _GEN_1080 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_254_data[32] ? 1'h0 : _GEN_964; // @[lut_35.scala 2834:105 lut_35.scala 177:26]
  wire  _GEN_1088 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_254_data[32] ? 1'h0 : _GEN_972; // @[lut_35.scala 2834:105 lut_35.scala 177:26]
  wire  _GEN_1096 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_254_data[32] ? 1'h0 : _GEN_980; // @[lut_35.scala 2834:105 lut_35.scala 177:26]
  wire  _GEN_1104 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_254_data[32] ? 1'h0 : _GEN_988; // @[lut_35.scala 2834:105 lut_35.scala 177:26]
  wire  _GEN_1112 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_254_data[32] ? 1'h0 : _GEN_996; // @[lut_35.scala 2834:105 lut_35.scala 177:26]
  wire  _GEN_1120 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_254_data[32] ? 1'h0 : _GEN_1004; // @[lut_35.scala 2834:105 lut_35.scala 177:26]
  wire  _GEN_1128 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_254_data[32] ? 1'h0 : _GEN_1012; // @[lut_35.scala 2834:105 lut_35.scala 177:26]
  wire  _GEN_1136 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_254_data[32] ? 1'h0 : _GEN_1020; // @[lut_35.scala 2834:105 lut_35.scala 177:26]
  wire  _GEN_1144 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_254_data[32] ? 1'h0 : _GEN_1028; // @[lut_35.scala 2834:105 lut_35.scala 177:26]
  wire  _GEN_1152 = io_empty_22 & push_valid & ~push_22_1 & ~LUT_mem_MPORT_254_data[32] ? 1'h0 : _GEN_1036; // @[lut_35.scala 2834:105 lut_35.scala 177:26]
  wire  _GEN_1164 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_252_data[32] ? 1'h0 : _T_526; // @[lut_35.scala 2794:105 lut_35.scala 2819:43]
  wire  _GEN_1165 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_252_data[32] ? 1'h0 : _GEN_1048; // @[lut_35.scala 2794:105 lut_35.scala 2820:43]
  wire  _GEN_1166 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_252_data[32] ? 1'h0 : _GEN_1049; // @[lut_35.scala 2794:105 lut_35.scala 2821:43]
  wire  _GEN_1167 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_252_data[32] ? 1'h0 : _GEN_1050; // @[lut_35.scala 2794:105 lut_35.scala 2822:43]
  wire  _GEN_1168 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_252_data[32] ? 1'h0 : _GEN_1051; // @[lut_35.scala 2794:105 lut_35.scala 2823:43]
  wire  _GEN_1169 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_252_data[32] ? 1'h0 : _GEN_1052; // @[lut_35.scala 2794:105 lut_35.scala 2824:43]
  wire  _GEN_1170 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_252_data[32] ? 1'h0 : _GEN_1053; // @[lut_35.scala 2794:105 lut_35.scala 2825:43]
  wire  _GEN_1171 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_252_data[32] ? 1'h0 : _GEN_1054; // @[lut_35.scala 2794:105 lut_35.scala 2826:43]
  wire  _GEN_1172 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_252_data[32] ? 1'h0 : _GEN_1055; // @[lut_35.scala 2794:105 lut_35.scala 2827:43]
  wire  _GEN_1173 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_252_data[32] ? 1'h0 : _GEN_1056; // @[lut_35.scala 2794:105 lut_35.scala 2828:43]
  wire  _GEN_1174 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_252_data[32] ? 1'h0 : _GEN_1057; // @[lut_35.scala 2794:105 lut_35.scala 2829:43]
  wire  _GEN_1175 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_252_data[32] ? 1'h0 : _GEN_1058; // @[lut_35.scala 2794:105 lut_35.scala 2830:43]
  wire  _GEN_1176 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_252_data[32] ? 1'h0 : _GEN_1059; // @[lut_35.scala 2794:105 lut_35.scala 2831:43]
  wire  _GEN_1177 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_252_data[32] | _GEN_1060; // @[lut_35.scala 2794:105 lut_35.scala 2832:38]
  wire  _GEN_1181 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_252_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2794:105 lut_35.scala 177:26 lut_35.scala 2834:89]
  wire  _GEN_1189 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_252_data[32] ? 1'h0 : _GEN_1064; // @[lut_35.scala 2794:105 lut_35.scala 177:26]
  wire  _GEN_1197 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_252_data[32] ? 1'h0 : _GEN_1072; // @[lut_35.scala 2794:105 lut_35.scala 177:26]
  wire  _GEN_1205 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_252_data[32] ? 1'h0 : _GEN_1080; // @[lut_35.scala 2794:105 lut_35.scala 177:26]
  wire  _GEN_1213 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_252_data[32] ? 1'h0 : _GEN_1088; // @[lut_35.scala 2794:105 lut_35.scala 177:26]
  wire  _GEN_1221 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_252_data[32] ? 1'h0 : _GEN_1096; // @[lut_35.scala 2794:105 lut_35.scala 177:26]
  wire  _GEN_1229 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_252_data[32] ? 1'h0 : _GEN_1104; // @[lut_35.scala 2794:105 lut_35.scala 177:26]
  wire  _GEN_1237 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_252_data[32] ? 1'h0 : _GEN_1112; // @[lut_35.scala 2794:105 lut_35.scala 177:26]
  wire  _GEN_1245 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_252_data[32] ? 1'h0 : _GEN_1120; // @[lut_35.scala 2794:105 lut_35.scala 177:26]
  wire  _GEN_1253 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_252_data[32] ? 1'h0 : _GEN_1128; // @[lut_35.scala 2794:105 lut_35.scala 177:26]
  wire  _GEN_1261 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_252_data[32] ? 1'h0 : _GEN_1136; // @[lut_35.scala 2794:105 lut_35.scala 177:26]
  wire  _GEN_1269 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_252_data[32] ? 1'h0 : _GEN_1144; // @[lut_35.scala 2794:105 lut_35.scala 177:26]
  wire  _GEN_1277 = io_empty_21 & push_valid & ~push_21_1 & ~LUT_mem_MPORT_252_data[32] ? 1'h0 : _GEN_1152; // @[lut_35.scala 2794:105 lut_35.scala 177:26]
  wire  _GEN_1289 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_250_data[32] ? 1'h0 : _T_517; // @[lut_35.scala 2754:105 lut_35.scala 2778:43]
  wire  _GEN_1290 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_250_data[32] ? 1'h0 : _GEN_1164; // @[lut_35.scala 2754:105 lut_35.scala 2779:43]
  wire  _GEN_1291 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_250_data[32] ? 1'h0 : _GEN_1165; // @[lut_35.scala 2754:105 lut_35.scala 2780:43]
  wire  _GEN_1292 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_250_data[32] ? 1'h0 : _GEN_1166; // @[lut_35.scala 2754:105 lut_35.scala 2781:43]
  wire  _GEN_1293 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_250_data[32] ? 1'h0 : _GEN_1167; // @[lut_35.scala 2754:105 lut_35.scala 2782:43]
  wire  _GEN_1294 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_250_data[32] ? 1'h0 : _GEN_1168; // @[lut_35.scala 2754:105 lut_35.scala 2783:43]
  wire  _GEN_1295 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_250_data[32] ? 1'h0 : _GEN_1169; // @[lut_35.scala 2754:105 lut_35.scala 2784:43]
  wire  _GEN_1296 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_250_data[32] ? 1'h0 : _GEN_1170; // @[lut_35.scala 2754:105 lut_35.scala 2785:43]
  wire  _GEN_1297 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_250_data[32] ? 1'h0 : _GEN_1171; // @[lut_35.scala 2754:105 lut_35.scala 2786:43]
  wire  _GEN_1298 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_250_data[32] ? 1'h0 : _GEN_1172; // @[lut_35.scala 2754:105 lut_35.scala 2787:43]
  wire  _GEN_1299 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_250_data[32] ? 1'h0 : _GEN_1173; // @[lut_35.scala 2754:105 lut_35.scala 2788:43]
  wire  _GEN_1300 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_250_data[32] ? 1'h0 : _GEN_1174; // @[lut_35.scala 2754:105 lut_35.scala 2789:43]
  wire  _GEN_1301 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_250_data[32] ? 1'h0 : _GEN_1175; // @[lut_35.scala 2754:105 lut_35.scala 2790:43]
  wire  _GEN_1302 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_250_data[32] ? 1'h0 : _GEN_1176; // @[lut_35.scala 2754:105 lut_35.scala 2791:43]
  wire  _GEN_1303 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_250_data[32] | _GEN_1177; // @[lut_35.scala 2754:105 lut_35.scala 2792:38]
  wire  _GEN_1307 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_250_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2754:105 lut_35.scala 177:26 lut_35.scala 2794:89]
  wire  _GEN_1315 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_250_data[32] ? 1'h0 : _GEN_1181; // @[lut_35.scala 2754:105 lut_35.scala 177:26]
  wire  _GEN_1323 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_250_data[32] ? 1'h0 : _GEN_1189; // @[lut_35.scala 2754:105 lut_35.scala 177:26]
  wire  _GEN_1331 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_250_data[32] ? 1'h0 : _GEN_1197; // @[lut_35.scala 2754:105 lut_35.scala 177:26]
  wire  _GEN_1339 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_250_data[32] ? 1'h0 : _GEN_1205; // @[lut_35.scala 2754:105 lut_35.scala 177:26]
  wire  _GEN_1347 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_250_data[32] ? 1'h0 : _GEN_1213; // @[lut_35.scala 2754:105 lut_35.scala 177:26]
  wire  _GEN_1355 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_250_data[32] ? 1'h0 : _GEN_1221; // @[lut_35.scala 2754:105 lut_35.scala 177:26]
  wire  _GEN_1363 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_250_data[32] ? 1'h0 : _GEN_1229; // @[lut_35.scala 2754:105 lut_35.scala 177:26]
  wire  _GEN_1371 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_250_data[32] ? 1'h0 : _GEN_1237; // @[lut_35.scala 2754:105 lut_35.scala 177:26]
  wire  _GEN_1379 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_250_data[32] ? 1'h0 : _GEN_1245; // @[lut_35.scala 2754:105 lut_35.scala 177:26]
  wire  _GEN_1387 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_250_data[32] ? 1'h0 : _GEN_1253; // @[lut_35.scala 2754:105 lut_35.scala 177:26]
  wire  _GEN_1395 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_250_data[32] ? 1'h0 : _GEN_1261; // @[lut_35.scala 2754:105 lut_35.scala 177:26]
  wire  _GEN_1403 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_250_data[32] ? 1'h0 : _GEN_1269; // @[lut_35.scala 2754:105 lut_35.scala 177:26]
  wire  _GEN_1411 = io_empty_20 & push_valid & ~push_20_1 & ~LUT_mem_MPORT_250_data[32] ? 1'h0 : _GEN_1277; // @[lut_35.scala 2754:105 lut_35.scala 177:26]
  wire  _GEN_1423 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_248_data[32] ? 1'h0 : _T_508; // @[lut_35.scala 2714:105 lut_35.scala 2737:43]
  wire  _GEN_1424 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_248_data[32] ? 1'h0 : _GEN_1289; // @[lut_35.scala 2714:105 lut_35.scala 2738:43]
  wire  _GEN_1425 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_248_data[32] ? 1'h0 : _GEN_1290; // @[lut_35.scala 2714:105 lut_35.scala 2739:43]
  wire  _GEN_1426 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_248_data[32] ? 1'h0 : _GEN_1291; // @[lut_35.scala 2714:105 lut_35.scala 2740:43]
  wire  _GEN_1427 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_248_data[32] ? 1'h0 : _GEN_1292; // @[lut_35.scala 2714:105 lut_35.scala 2741:43]
  wire  _GEN_1428 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_248_data[32] ? 1'h0 : _GEN_1293; // @[lut_35.scala 2714:105 lut_35.scala 2742:43]
  wire  _GEN_1429 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_248_data[32] ? 1'h0 : _GEN_1294; // @[lut_35.scala 2714:105 lut_35.scala 2743:43]
  wire  _GEN_1430 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_248_data[32] ? 1'h0 : _GEN_1295; // @[lut_35.scala 2714:105 lut_35.scala 2744:43]
  wire  _GEN_1431 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_248_data[32] ? 1'h0 : _GEN_1296; // @[lut_35.scala 2714:105 lut_35.scala 2745:43]
  wire  _GEN_1432 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_248_data[32] ? 1'h0 : _GEN_1297; // @[lut_35.scala 2714:105 lut_35.scala 2746:43]
  wire  _GEN_1433 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_248_data[32] ? 1'h0 : _GEN_1298; // @[lut_35.scala 2714:105 lut_35.scala 2747:43]
  wire  _GEN_1434 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_248_data[32] ? 1'h0 : _GEN_1299; // @[lut_35.scala 2714:105 lut_35.scala 2748:43]
  wire  _GEN_1435 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_248_data[32] ? 1'h0 : _GEN_1300; // @[lut_35.scala 2714:105 lut_35.scala 2749:43]
  wire  _GEN_1436 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_248_data[32] ? 1'h0 : _GEN_1301; // @[lut_35.scala 2714:105 lut_35.scala 2750:43]
  wire  _GEN_1437 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_248_data[32] ? 1'h0 : _GEN_1302; // @[lut_35.scala 2714:105 lut_35.scala 2751:43]
  wire  _GEN_1438 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_248_data[32] | _GEN_1303; // @[lut_35.scala 2714:105 lut_35.scala 2752:38]
  wire  _GEN_1442 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_248_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2714:105 lut_35.scala 177:26 lut_35.scala 2754:89]
  wire  _GEN_1450 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_248_data[32] ? 1'h0 : _GEN_1307; // @[lut_35.scala 2714:105 lut_35.scala 177:26]
  wire  _GEN_1458 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_248_data[32] ? 1'h0 : _GEN_1315; // @[lut_35.scala 2714:105 lut_35.scala 177:26]
  wire  _GEN_1466 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_248_data[32] ? 1'h0 : _GEN_1323; // @[lut_35.scala 2714:105 lut_35.scala 177:26]
  wire  _GEN_1474 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_248_data[32] ? 1'h0 : _GEN_1331; // @[lut_35.scala 2714:105 lut_35.scala 177:26]
  wire  _GEN_1482 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_248_data[32] ? 1'h0 : _GEN_1339; // @[lut_35.scala 2714:105 lut_35.scala 177:26]
  wire  _GEN_1490 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_248_data[32] ? 1'h0 : _GEN_1347; // @[lut_35.scala 2714:105 lut_35.scala 177:26]
  wire  _GEN_1498 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_248_data[32] ? 1'h0 : _GEN_1355; // @[lut_35.scala 2714:105 lut_35.scala 177:26]
  wire  _GEN_1506 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_248_data[32] ? 1'h0 : _GEN_1363; // @[lut_35.scala 2714:105 lut_35.scala 177:26]
  wire  _GEN_1514 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_248_data[32] ? 1'h0 : _GEN_1371; // @[lut_35.scala 2714:105 lut_35.scala 177:26]
  wire  _GEN_1522 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_248_data[32] ? 1'h0 : _GEN_1379; // @[lut_35.scala 2714:105 lut_35.scala 177:26]
  wire  _GEN_1530 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_248_data[32] ? 1'h0 : _GEN_1387; // @[lut_35.scala 2714:105 lut_35.scala 177:26]
  wire  _GEN_1538 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_248_data[32] ? 1'h0 : _GEN_1395; // @[lut_35.scala 2714:105 lut_35.scala 177:26]
  wire  _GEN_1546 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_248_data[32] ? 1'h0 : _GEN_1403; // @[lut_35.scala 2714:105 lut_35.scala 177:26]
  wire  _GEN_1554 = io_empty_19 & push_valid & ~push_19_1 & ~LUT_mem_MPORT_248_data[32] ? 1'h0 : _GEN_1411; // @[lut_35.scala 2714:105 lut_35.scala 177:26]
  wire  _GEN_1566 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_246_data[32] ? 1'h0 : _T_499; // @[lut_35.scala 2674:105 lut_35.scala 2696:43]
  wire  _GEN_1567 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_246_data[32] ? 1'h0 : _GEN_1423; // @[lut_35.scala 2674:105 lut_35.scala 2697:43]
  wire  _GEN_1568 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_246_data[32] ? 1'h0 : _GEN_1424; // @[lut_35.scala 2674:105 lut_35.scala 2698:43]
  wire  _GEN_1569 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_246_data[32] ? 1'h0 : _GEN_1425; // @[lut_35.scala 2674:105 lut_35.scala 2699:43]
  wire  _GEN_1570 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_246_data[32] ? 1'h0 : _GEN_1426; // @[lut_35.scala 2674:105 lut_35.scala 2700:43]
  wire  _GEN_1571 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_246_data[32] ? 1'h0 : _GEN_1427; // @[lut_35.scala 2674:105 lut_35.scala 2701:43]
  wire  _GEN_1572 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_246_data[32] ? 1'h0 : _GEN_1428; // @[lut_35.scala 2674:105 lut_35.scala 2702:43]
  wire  _GEN_1573 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_246_data[32] ? 1'h0 : _GEN_1429; // @[lut_35.scala 2674:105 lut_35.scala 2703:43]
  wire  _GEN_1574 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_246_data[32] ? 1'h0 : _GEN_1430; // @[lut_35.scala 2674:105 lut_35.scala 2704:43]
  wire  _GEN_1575 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_246_data[32] ? 1'h0 : _GEN_1431; // @[lut_35.scala 2674:105 lut_35.scala 2705:43]
  wire  _GEN_1576 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_246_data[32] ? 1'h0 : _GEN_1432; // @[lut_35.scala 2674:105 lut_35.scala 2706:43]
  wire  _GEN_1577 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_246_data[32] ? 1'h0 : _GEN_1433; // @[lut_35.scala 2674:105 lut_35.scala 2707:43]
  wire  _GEN_1578 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_246_data[32] ? 1'h0 : _GEN_1434; // @[lut_35.scala 2674:105 lut_35.scala 2708:43]
  wire  _GEN_1579 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_246_data[32] ? 1'h0 : _GEN_1435; // @[lut_35.scala 2674:105 lut_35.scala 2709:43]
  wire  _GEN_1580 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_246_data[32] ? 1'h0 : _GEN_1436; // @[lut_35.scala 2674:105 lut_35.scala 2710:43]
  wire  _GEN_1581 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_246_data[32] ? 1'h0 : _GEN_1437; // @[lut_35.scala 2674:105 lut_35.scala 2711:43]
  wire  _GEN_1582 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_246_data[32] | _GEN_1438; // @[lut_35.scala 2674:105 lut_35.scala 2712:38]
  wire  _GEN_1586 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_246_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2674:105 lut_35.scala 177:26 lut_35.scala 2714:89]
  wire  _GEN_1594 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_246_data[32] ? 1'h0 : _GEN_1442; // @[lut_35.scala 2674:105 lut_35.scala 177:26]
  wire  _GEN_1602 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_246_data[32] ? 1'h0 : _GEN_1450; // @[lut_35.scala 2674:105 lut_35.scala 177:26]
  wire  _GEN_1610 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_246_data[32] ? 1'h0 : _GEN_1458; // @[lut_35.scala 2674:105 lut_35.scala 177:26]
  wire  _GEN_1618 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_246_data[32] ? 1'h0 : _GEN_1466; // @[lut_35.scala 2674:105 lut_35.scala 177:26]
  wire  _GEN_1626 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_246_data[32] ? 1'h0 : _GEN_1474; // @[lut_35.scala 2674:105 lut_35.scala 177:26]
  wire  _GEN_1634 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_246_data[32] ? 1'h0 : _GEN_1482; // @[lut_35.scala 2674:105 lut_35.scala 177:26]
  wire  _GEN_1642 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_246_data[32] ? 1'h0 : _GEN_1490; // @[lut_35.scala 2674:105 lut_35.scala 177:26]
  wire  _GEN_1650 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_246_data[32] ? 1'h0 : _GEN_1498; // @[lut_35.scala 2674:105 lut_35.scala 177:26]
  wire  _GEN_1658 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_246_data[32] ? 1'h0 : _GEN_1506; // @[lut_35.scala 2674:105 lut_35.scala 177:26]
  wire  _GEN_1666 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_246_data[32] ? 1'h0 : _GEN_1514; // @[lut_35.scala 2674:105 lut_35.scala 177:26]
  wire  _GEN_1674 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_246_data[32] ? 1'h0 : _GEN_1522; // @[lut_35.scala 2674:105 lut_35.scala 177:26]
  wire  _GEN_1682 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_246_data[32] ? 1'h0 : _GEN_1530; // @[lut_35.scala 2674:105 lut_35.scala 177:26]
  wire  _GEN_1690 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_246_data[32] ? 1'h0 : _GEN_1538; // @[lut_35.scala 2674:105 lut_35.scala 177:26]
  wire  _GEN_1698 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_246_data[32] ? 1'h0 : _GEN_1546; // @[lut_35.scala 2674:105 lut_35.scala 177:26]
  wire  _GEN_1706 = io_empty_18 & push_valid & ~push_18_1 & ~LUT_mem_MPORT_246_data[32] ? 1'h0 : _GEN_1554; // @[lut_35.scala 2674:105 lut_35.scala 177:26]
  wire  _GEN_1718 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_244_data[32] ? 1'h0 : _T_490; // @[lut_35.scala 2634:105 lut_35.scala 2655:43]
  wire  _GEN_1719 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_244_data[32] ? 1'h0 : _GEN_1566; // @[lut_35.scala 2634:105 lut_35.scala 2656:43]
  wire  _GEN_1720 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_244_data[32] ? 1'h0 : _GEN_1567; // @[lut_35.scala 2634:105 lut_35.scala 2657:43]
  wire  _GEN_1721 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_244_data[32] ? 1'h0 : _GEN_1568; // @[lut_35.scala 2634:105 lut_35.scala 2658:43]
  wire  _GEN_1722 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_244_data[32] ? 1'h0 : _GEN_1569; // @[lut_35.scala 2634:105 lut_35.scala 2659:43]
  wire  _GEN_1723 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_244_data[32] ? 1'h0 : _GEN_1570; // @[lut_35.scala 2634:105 lut_35.scala 2660:43]
  wire  _GEN_1724 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_244_data[32] ? 1'h0 : _GEN_1571; // @[lut_35.scala 2634:105 lut_35.scala 2661:43]
  wire  _GEN_1725 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_244_data[32] ? 1'h0 : _GEN_1572; // @[lut_35.scala 2634:105 lut_35.scala 2662:43]
  wire  _GEN_1726 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_244_data[32] ? 1'h0 : _GEN_1573; // @[lut_35.scala 2634:105 lut_35.scala 2663:43]
  wire  _GEN_1727 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_244_data[32] ? 1'h0 : _GEN_1574; // @[lut_35.scala 2634:105 lut_35.scala 2664:43]
  wire  _GEN_1728 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_244_data[32] ? 1'h0 : _GEN_1575; // @[lut_35.scala 2634:105 lut_35.scala 2665:43]
  wire  _GEN_1729 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_244_data[32] ? 1'h0 : _GEN_1576; // @[lut_35.scala 2634:105 lut_35.scala 2666:43]
  wire  _GEN_1730 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_244_data[32] ? 1'h0 : _GEN_1577; // @[lut_35.scala 2634:105 lut_35.scala 2667:43]
  wire  _GEN_1731 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_244_data[32] ? 1'h0 : _GEN_1578; // @[lut_35.scala 2634:105 lut_35.scala 2668:43]
  wire  _GEN_1732 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_244_data[32] ? 1'h0 : _GEN_1579; // @[lut_35.scala 2634:105 lut_35.scala 2669:43]
  wire  _GEN_1733 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_244_data[32] ? 1'h0 : _GEN_1580; // @[lut_35.scala 2634:105 lut_35.scala 2670:43]
  wire  _GEN_1734 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_244_data[32] ? 1'h0 : _GEN_1581; // @[lut_35.scala 2634:105 lut_35.scala 2671:43]
  wire  _GEN_1735 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_244_data[32] | _GEN_1582; // @[lut_35.scala 2634:105 lut_35.scala 2672:38]
  wire  _GEN_1739 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_244_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2634:105 lut_35.scala 177:26 lut_35.scala 2674:89]
  wire  _GEN_1747 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_244_data[32] ? 1'h0 : _GEN_1586; // @[lut_35.scala 2634:105 lut_35.scala 177:26]
  wire  _GEN_1755 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_244_data[32] ? 1'h0 : _GEN_1594; // @[lut_35.scala 2634:105 lut_35.scala 177:26]
  wire  _GEN_1763 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_244_data[32] ? 1'h0 : _GEN_1602; // @[lut_35.scala 2634:105 lut_35.scala 177:26]
  wire  _GEN_1771 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_244_data[32] ? 1'h0 : _GEN_1610; // @[lut_35.scala 2634:105 lut_35.scala 177:26]
  wire  _GEN_1779 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_244_data[32] ? 1'h0 : _GEN_1618; // @[lut_35.scala 2634:105 lut_35.scala 177:26]
  wire  _GEN_1787 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_244_data[32] ? 1'h0 : _GEN_1626; // @[lut_35.scala 2634:105 lut_35.scala 177:26]
  wire  _GEN_1795 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_244_data[32] ? 1'h0 : _GEN_1634; // @[lut_35.scala 2634:105 lut_35.scala 177:26]
  wire  _GEN_1803 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_244_data[32] ? 1'h0 : _GEN_1642; // @[lut_35.scala 2634:105 lut_35.scala 177:26]
  wire  _GEN_1811 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_244_data[32] ? 1'h0 : _GEN_1650; // @[lut_35.scala 2634:105 lut_35.scala 177:26]
  wire  _GEN_1819 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_244_data[32] ? 1'h0 : _GEN_1658; // @[lut_35.scala 2634:105 lut_35.scala 177:26]
  wire  _GEN_1827 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_244_data[32] ? 1'h0 : _GEN_1666; // @[lut_35.scala 2634:105 lut_35.scala 177:26]
  wire  _GEN_1835 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_244_data[32] ? 1'h0 : _GEN_1674; // @[lut_35.scala 2634:105 lut_35.scala 177:26]
  wire  _GEN_1843 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_244_data[32] ? 1'h0 : _GEN_1682; // @[lut_35.scala 2634:105 lut_35.scala 177:26]
  wire  _GEN_1851 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_244_data[32] ? 1'h0 : _GEN_1690; // @[lut_35.scala 2634:105 lut_35.scala 177:26]
  wire  _GEN_1859 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_244_data[32] ? 1'h0 : _GEN_1698; // @[lut_35.scala 2634:105 lut_35.scala 177:26]
  wire  _GEN_1867 = io_empty_17 & push_valid & ~push_17_1 & ~LUT_mem_MPORT_244_data[32] ? 1'h0 : _GEN_1706; // @[lut_35.scala 2634:105 lut_35.scala 177:26]
  wire  _GEN_1879 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_242_data[32] ? 1'h0 : _T_481; // @[lut_35.scala 2594:105 lut_35.scala 2614:43]
  wire  _GEN_1880 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_242_data[32] ? 1'h0 : _GEN_1718; // @[lut_35.scala 2594:105 lut_35.scala 2615:43]
  wire  _GEN_1881 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_242_data[32] ? 1'h0 : _GEN_1719; // @[lut_35.scala 2594:105 lut_35.scala 2616:43]
  wire  _GEN_1882 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_242_data[32] ? 1'h0 : _GEN_1720; // @[lut_35.scala 2594:105 lut_35.scala 2617:43]
  wire  _GEN_1883 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_242_data[32] ? 1'h0 : _GEN_1721; // @[lut_35.scala 2594:105 lut_35.scala 2618:43]
  wire  _GEN_1884 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_242_data[32] ? 1'h0 : _GEN_1722; // @[lut_35.scala 2594:105 lut_35.scala 2619:43]
  wire  _GEN_1885 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_242_data[32] ? 1'h0 : _GEN_1723; // @[lut_35.scala 2594:105 lut_35.scala 2620:43]
  wire  _GEN_1886 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_242_data[32] ? 1'h0 : _GEN_1724; // @[lut_35.scala 2594:105 lut_35.scala 2621:43]
  wire  _GEN_1887 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_242_data[32] ? 1'h0 : _GEN_1725; // @[lut_35.scala 2594:105 lut_35.scala 2622:43]
  wire  _GEN_1888 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_242_data[32] ? 1'h0 : _GEN_1726; // @[lut_35.scala 2594:105 lut_35.scala 2623:43]
  wire  _GEN_1889 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_242_data[32] ? 1'h0 : _GEN_1727; // @[lut_35.scala 2594:105 lut_35.scala 2624:43]
  wire  _GEN_1890 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_242_data[32] ? 1'h0 : _GEN_1728; // @[lut_35.scala 2594:105 lut_35.scala 2625:43]
  wire  _GEN_1891 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_242_data[32] ? 1'h0 : _GEN_1729; // @[lut_35.scala 2594:105 lut_35.scala 2626:43]
  wire  _GEN_1892 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_242_data[32] ? 1'h0 : _GEN_1730; // @[lut_35.scala 2594:105 lut_35.scala 2627:43]
  wire  _GEN_1893 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_242_data[32] ? 1'h0 : _GEN_1731; // @[lut_35.scala 2594:105 lut_35.scala 2628:43]
  wire  _GEN_1894 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_242_data[32] ? 1'h0 : _GEN_1732; // @[lut_35.scala 2594:105 lut_35.scala 2629:43]
  wire  _GEN_1895 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_242_data[32] ? 1'h0 : _GEN_1733; // @[lut_35.scala 2594:105 lut_35.scala 2630:43]
  wire  _GEN_1896 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_242_data[32] ? 1'h0 : _GEN_1734; // @[lut_35.scala 2594:105 lut_35.scala 2631:43]
  wire  _GEN_1897 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_242_data[32] | _GEN_1735; // @[lut_35.scala 2594:105 lut_35.scala 2632:38]
  wire  _GEN_1901 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_242_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2594:105 lut_35.scala 177:26 lut_35.scala 2634:89]
  wire  _GEN_1909 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_242_data[32] ? 1'h0 : _GEN_1739; // @[lut_35.scala 2594:105 lut_35.scala 177:26]
  wire  _GEN_1917 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_242_data[32] ? 1'h0 : _GEN_1747; // @[lut_35.scala 2594:105 lut_35.scala 177:26]
  wire  _GEN_1925 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_242_data[32] ? 1'h0 : _GEN_1755; // @[lut_35.scala 2594:105 lut_35.scala 177:26]
  wire  _GEN_1933 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_242_data[32] ? 1'h0 : _GEN_1763; // @[lut_35.scala 2594:105 lut_35.scala 177:26]
  wire  _GEN_1941 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_242_data[32] ? 1'h0 : _GEN_1771; // @[lut_35.scala 2594:105 lut_35.scala 177:26]
  wire  _GEN_1949 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_242_data[32] ? 1'h0 : _GEN_1779; // @[lut_35.scala 2594:105 lut_35.scala 177:26]
  wire  _GEN_1957 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_242_data[32] ? 1'h0 : _GEN_1787; // @[lut_35.scala 2594:105 lut_35.scala 177:26]
  wire  _GEN_1965 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_242_data[32] ? 1'h0 : _GEN_1795; // @[lut_35.scala 2594:105 lut_35.scala 177:26]
  wire  _GEN_1973 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_242_data[32] ? 1'h0 : _GEN_1803; // @[lut_35.scala 2594:105 lut_35.scala 177:26]
  wire  _GEN_1981 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_242_data[32] ? 1'h0 : _GEN_1811; // @[lut_35.scala 2594:105 lut_35.scala 177:26]
  wire  _GEN_1989 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_242_data[32] ? 1'h0 : _GEN_1819; // @[lut_35.scala 2594:105 lut_35.scala 177:26]
  wire  _GEN_1997 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_242_data[32] ? 1'h0 : _GEN_1827; // @[lut_35.scala 2594:105 lut_35.scala 177:26]
  wire  _GEN_2005 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_242_data[32] ? 1'h0 : _GEN_1835; // @[lut_35.scala 2594:105 lut_35.scala 177:26]
  wire  _GEN_2013 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_242_data[32] ? 1'h0 : _GEN_1843; // @[lut_35.scala 2594:105 lut_35.scala 177:26]
  wire  _GEN_2021 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_242_data[32] ? 1'h0 : _GEN_1851; // @[lut_35.scala 2594:105 lut_35.scala 177:26]
  wire  _GEN_2029 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_242_data[32] ? 1'h0 : _GEN_1859; // @[lut_35.scala 2594:105 lut_35.scala 177:26]
  wire  _GEN_2037 = io_empty_16 & push_valid & ~push_16_1 & ~LUT_mem_MPORT_242_data[32] ? 1'h0 : _GEN_1867; // @[lut_35.scala 2594:105 lut_35.scala 177:26]
  wire  _GEN_2049 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_240_data[32] ? 1'h0 : _T_472; // @[lut_35.scala 2554:105 lut_35.scala 2573:43]
  wire  _GEN_2050 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_240_data[32] ? 1'h0 : _GEN_1879; // @[lut_35.scala 2554:105 lut_35.scala 2574:43]
  wire  _GEN_2051 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_240_data[32] ? 1'h0 : _GEN_1880; // @[lut_35.scala 2554:105 lut_35.scala 2575:43]
  wire  _GEN_2052 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_240_data[32] ? 1'h0 : _GEN_1881; // @[lut_35.scala 2554:105 lut_35.scala 2576:43]
  wire  _GEN_2053 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_240_data[32] ? 1'h0 : _GEN_1882; // @[lut_35.scala 2554:105 lut_35.scala 2577:43]
  wire  _GEN_2054 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_240_data[32] ? 1'h0 : _GEN_1883; // @[lut_35.scala 2554:105 lut_35.scala 2578:43]
  wire  _GEN_2055 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_240_data[32] ? 1'h0 : _GEN_1884; // @[lut_35.scala 2554:105 lut_35.scala 2579:43]
  wire  _GEN_2056 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_240_data[32] ? 1'h0 : _GEN_1885; // @[lut_35.scala 2554:105 lut_35.scala 2580:43]
  wire  _GEN_2057 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_240_data[32] ? 1'h0 : _GEN_1886; // @[lut_35.scala 2554:105 lut_35.scala 2581:43]
  wire  _GEN_2058 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_240_data[32] ? 1'h0 : _GEN_1887; // @[lut_35.scala 2554:105 lut_35.scala 2582:43]
  wire  _GEN_2059 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_240_data[32] ? 1'h0 : _GEN_1888; // @[lut_35.scala 2554:105 lut_35.scala 2583:43]
  wire  _GEN_2060 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_240_data[32] ? 1'h0 : _GEN_1889; // @[lut_35.scala 2554:105 lut_35.scala 2584:43]
  wire  _GEN_2061 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_240_data[32] ? 1'h0 : _GEN_1890; // @[lut_35.scala 2554:105 lut_35.scala 2585:43]
  wire  _GEN_2062 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_240_data[32] ? 1'h0 : _GEN_1891; // @[lut_35.scala 2554:105 lut_35.scala 2586:43]
  wire  _GEN_2063 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_240_data[32] ? 1'h0 : _GEN_1892; // @[lut_35.scala 2554:105 lut_35.scala 2587:43]
  wire  _GEN_2064 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_240_data[32] ? 1'h0 : _GEN_1893; // @[lut_35.scala 2554:105 lut_35.scala 2588:43]
  wire  _GEN_2065 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_240_data[32] ? 1'h0 : _GEN_1894; // @[lut_35.scala 2554:105 lut_35.scala 2589:43]
  wire  _GEN_2066 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_240_data[32] ? 1'h0 : _GEN_1895; // @[lut_35.scala 2554:105 lut_35.scala 2590:43]
  wire  _GEN_2067 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_240_data[32] ? 1'h0 : _GEN_1896; // @[lut_35.scala 2554:105 lut_35.scala 2591:43]
  wire  _GEN_2068 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_240_data[32] | _GEN_1897; // @[lut_35.scala 2554:105 lut_35.scala 2592:38]
  wire  _GEN_2072 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_240_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2554:105 lut_35.scala 177:26 lut_35.scala 2594:89]
  wire  _GEN_2080 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_240_data[32] ? 1'h0 : _GEN_1901; // @[lut_35.scala 2554:105 lut_35.scala 177:26]
  wire  _GEN_2088 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_240_data[32] ? 1'h0 : _GEN_1909; // @[lut_35.scala 2554:105 lut_35.scala 177:26]
  wire  _GEN_2096 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_240_data[32] ? 1'h0 : _GEN_1917; // @[lut_35.scala 2554:105 lut_35.scala 177:26]
  wire  _GEN_2104 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_240_data[32] ? 1'h0 : _GEN_1925; // @[lut_35.scala 2554:105 lut_35.scala 177:26]
  wire  _GEN_2112 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_240_data[32] ? 1'h0 : _GEN_1933; // @[lut_35.scala 2554:105 lut_35.scala 177:26]
  wire  _GEN_2120 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_240_data[32] ? 1'h0 : _GEN_1941; // @[lut_35.scala 2554:105 lut_35.scala 177:26]
  wire  _GEN_2128 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_240_data[32] ? 1'h0 : _GEN_1949; // @[lut_35.scala 2554:105 lut_35.scala 177:26]
  wire  _GEN_2136 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_240_data[32] ? 1'h0 : _GEN_1957; // @[lut_35.scala 2554:105 lut_35.scala 177:26]
  wire  _GEN_2144 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_240_data[32] ? 1'h0 : _GEN_1965; // @[lut_35.scala 2554:105 lut_35.scala 177:26]
  wire  _GEN_2152 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_240_data[32] ? 1'h0 : _GEN_1973; // @[lut_35.scala 2554:105 lut_35.scala 177:26]
  wire  _GEN_2160 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_240_data[32] ? 1'h0 : _GEN_1981; // @[lut_35.scala 2554:105 lut_35.scala 177:26]
  wire  _GEN_2168 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_240_data[32] ? 1'h0 : _GEN_1989; // @[lut_35.scala 2554:105 lut_35.scala 177:26]
  wire  _GEN_2176 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_240_data[32] ? 1'h0 : _GEN_1997; // @[lut_35.scala 2554:105 lut_35.scala 177:26]
  wire  _GEN_2184 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_240_data[32] ? 1'h0 : _GEN_2005; // @[lut_35.scala 2554:105 lut_35.scala 177:26]
  wire  _GEN_2192 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_240_data[32] ? 1'h0 : _GEN_2013; // @[lut_35.scala 2554:105 lut_35.scala 177:26]
  wire  _GEN_2200 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_240_data[32] ? 1'h0 : _GEN_2021; // @[lut_35.scala 2554:105 lut_35.scala 177:26]
  wire  _GEN_2208 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_240_data[32] ? 1'h0 : _GEN_2029; // @[lut_35.scala 2554:105 lut_35.scala 177:26]
  wire  _GEN_2216 = io_empty_15 & push_valid & ~push_15_1 & ~LUT_mem_MPORT_240_data[32] ? 1'h0 : _GEN_2037; // @[lut_35.scala 2554:105 lut_35.scala 177:26]
  wire  _GEN_2228 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_238_data[32] ? 1'h0 : _T_463; // @[lut_35.scala 2514:105 lut_35.scala 2532:43]
  wire  _GEN_2229 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_238_data[32] ? 1'h0 : _GEN_2049; // @[lut_35.scala 2514:105 lut_35.scala 2533:43]
  wire  _GEN_2230 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_238_data[32] ? 1'h0 : _GEN_2050; // @[lut_35.scala 2514:105 lut_35.scala 2534:43]
  wire  _GEN_2231 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_238_data[32] ? 1'h0 : _GEN_2051; // @[lut_35.scala 2514:105 lut_35.scala 2535:43]
  wire  _GEN_2232 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_238_data[32] ? 1'h0 : _GEN_2052; // @[lut_35.scala 2514:105 lut_35.scala 2536:43]
  wire  _GEN_2233 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_238_data[32] ? 1'h0 : _GEN_2053; // @[lut_35.scala 2514:105 lut_35.scala 2537:43]
  wire  _GEN_2234 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_238_data[32] ? 1'h0 : _GEN_2054; // @[lut_35.scala 2514:105 lut_35.scala 2538:43]
  wire  _GEN_2235 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_238_data[32] ? 1'h0 : _GEN_2055; // @[lut_35.scala 2514:105 lut_35.scala 2539:43]
  wire  _GEN_2236 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_238_data[32] ? 1'h0 : _GEN_2056; // @[lut_35.scala 2514:105 lut_35.scala 2540:43]
  wire  _GEN_2237 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_238_data[32] ? 1'h0 : _GEN_2057; // @[lut_35.scala 2514:105 lut_35.scala 2541:43]
  wire  _GEN_2238 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_238_data[32] ? 1'h0 : _GEN_2058; // @[lut_35.scala 2514:105 lut_35.scala 2542:43]
  wire  _GEN_2239 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_238_data[32] ? 1'h0 : _GEN_2059; // @[lut_35.scala 2514:105 lut_35.scala 2543:43]
  wire  _GEN_2240 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_238_data[32] ? 1'h0 : _GEN_2060; // @[lut_35.scala 2514:105 lut_35.scala 2544:43]
  wire  _GEN_2241 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_238_data[32] ? 1'h0 : _GEN_2061; // @[lut_35.scala 2514:105 lut_35.scala 2545:43]
  wire  _GEN_2242 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_238_data[32] ? 1'h0 : _GEN_2062; // @[lut_35.scala 2514:105 lut_35.scala 2546:43]
  wire  _GEN_2243 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_238_data[32] ? 1'h0 : _GEN_2063; // @[lut_35.scala 2514:105 lut_35.scala 2547:43]
  wire  _GEN_2244 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_238_data[32] ? 1'h0 : _GEN_2064; // @[lut_35.scala 2514:105 lut_35.scala 2548:43]
  wire  _GEN_2245 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_238_data[32] ? 1'h0 : _GEN_2065; // @[lut_35.scala 2514:105 lut_35.scala 2549:43]
  wire  _GEN_2246 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_238_data[32] ? 1'h0 : _GEN_2066; // @[lut_35.scala 2514:105 lut_35.scala 2550:43]
  wire  _GEN_2247 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_238_data[32] ? 1'h0 : _GEN_2067; // @[lut_35.scala 2514:105 lut_35.scala 2551:43]
  wire  _GEN_2248 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_238_data[32] | _GEN_2068; // @[lut_35.scala 2514:105 lut_35.scala 2552:38]
  wire  _GEN_2252 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_238_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2514:105 lut_35.scala 177:26 lut_35.scala 2554:89]
  wire  _GEN_2260 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_238_data[32] ? 1'h0 : _GEN_2072; // @[lut_35.scala 2514:105 lut_35.scala 177:26]
  wire  _GEN_2268 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_238_data[32] ? 1'h0 : _GEN_2080; // @[lut_35.scala 2514:105 lut_35.scala 177:26]
  wire  _GEN_2276 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_238_data[32] ? 1'h0 : _GEN_2088; // @[lut_35.scala 2514:105 lut_35.scala 177:26]
  wire  _GEN_2284 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_238_data[32] ? 1'h0 : _GEN_2096; // @[lut_35.scala 2514:105 lut_35.scala 177:26]
  wire  _GEN_2292 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_238_data[32] ? 1'h0 : _GEN_2104; // @[lut_35.scala 2514:105 lut_35.scala 177:26]
  wire  _GEN_2300 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_238_data[32] ? 1'h0 : _GEN_2112; // @[lut_35.scala 2514:105 lut_35.scala 177:26]
  wire  _GEN_2308 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_238_data[32] ? 1'h0 : _GEN_2120; // @[lut_35.scala 2514:105 lut_35.scala 177:26]
  wire  _GEN_2316 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_238_data[32] ? 1'h0 : _GEN_2128; // @[lut_35.scala 2514:105 lut_35.scala 177:26]
  wire  _GEN_2324 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_238_data[32] ? 1'h0 : _GEN_2136; // @[lut_35.scala 2514:105 lut_35.scala 177:26]
  wire  _GEN_2332 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_238_data[32] ? 1'h0 : _GEN_2144; // @[lut_35.scala 2514:105 lut_35.scala 177:26]
  wire  _GEN_2340 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_238_data[32] ? 1'h0 : _GEN_2152; // @[lut_35.scala 2514:105 lut_35.scala 177:26]
  wire  _GEN_2348 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_238_data[32] ? 1'h0 : _GEN_2160; // @[lut_35.scala 2514:105 lut_35.scala 177:26]
  wire  _GEN_2356 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_238_data[32] ? 1'h0 : _GEN_2168; // @[lut_35.scala 2514:105 lut_35.scala 177:26]
  wire  _GEN_2364 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_238_data[32] ? 1'h0 : _GEN_2176; // @[lut_35.scala 2514:105 lut_35.scala 177:26]
  wire  _GEN_2372 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_238_data[32] ? 1'h0 : _GEN_2184; // @[lut_35.scala 2514:105 lut_35.scala 177:26]
  wire  _GEN_2380 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_238_data[32] ? 1'h0 : _GEN_2192; // @[lut_35.scala 2514:105 lut_35.scala 177:26]
  wire  _GEN_2388 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_238_data[32] ? 1'h0 : _GEN_2200; // @[lut_35.scala 2514:105 lut_35.scala 177:26]
  wire  _GEN_2396 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_238_data[32] ? 1'h0 : _GEN_2208; // @[lut_35.scala 2514:105 lut_35.scala 177:26]
  wire  _GEN_2404 = io_empty_14 & push_valid & ~push_14_1 & ~LUT_mem_MPORT_238_data[32] ? 1'h0 : _GEN_2216; // @[lut_35.scala 2514:105 lut_35.scala 177:26]
  wire  _GEN_2416 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] ? 1'h0 : _T_454; // @[lut_35.scala 2474:105 lut_35.scala 2491:43]
  wire  _GEN_2417 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] ? 1'h0 : _GEN_2228; // @[lut_35.scala 2474:105 lut_35.scala 2492:43]
  wire  _GEN_2418 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] ? 1'h0 : _GEN_2229; // @[lut_35.scala 2474:105 lut_35.scala 2493:43]
  wire  _GEN_2419 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] ? 1'h0 : _GEN_2230; // @[lut_35.scala 2474:105 lut_35.scala 2494:43]
  wire  _GEN_2420 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] ? 1'h0 : _GEN_2231; // @[lut_35.scala 2474:105 lut_35.scala 2495:43]
  wire  _GEN_2421 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] ? 1'h0 : _GEN_2232; // @[lut_35.scala 2474:105 lut_35.scala 2496:43]
  wire  _GEN_2422 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] ? 1'h0 : _GEN_2233; // @[lut_35.scala 2474:105 lut_35.scala 2497:43]
  wire  _GEN_2423 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] ? 1'h0 : _GEN_2234; // @[lut_35.scala 2474:105 lut_35.scala 2498:43]
  wire  _GEN_2424 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] ? 1'h0 : _GEN_2235; // @[lut_35.scala 2474:105 lut_35.scala 2499:43]
  wire  _GEN_2425 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] ? 1'h0 : _GEN_2236; // @[lut_35.scala 2474:105 lut_35.scala 2500:43]
  wire  _GEN_2426 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] ? 1'h0 : _GEN_2237; // @[lut_35.scala 2474:105 lut_35.scala 2501:43]
  wire  _GEN_2427 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] ? 1'h0 : _GEN_2238; // @[lut_35.scala 2474:105 lut_35.scala 2502:43]
  wire  _GEN_2428 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] ? 1'h0 : _GEN_2239; // @[lut_35.scala 2474:105 lut_35.scala 2503:43]
  wire  _GEN_2429 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] ? 1'h0 : _GEN_2240; // @[lut_35.scala 2474:105 lut_35.scala 2504:43]
  wire  _GEN_2430 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] ? 1'h0 : _GEN_2241; // @[lut_35.scala 2474:105 lut_35.scala 2505:43]
  wire  _GEN_2431 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] ? 1'h0 : _GEN_2242; // @[lut_35.scala 2474:105 lut_35.scala 2506:43]
  wire  _GEN_2432 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] ? 1'h0 : _GEN_2243; // @[lut_35.scala 2474:105 lut_35.scala 2507:43]
  wire  _GEN_2433 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] ? 1'h0 : _GEN_2244; // @[lut_35.scala 2474:105 lut_35.scala 2508:43]
  wire  _GEN_2434 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] ? 1'h0 : _GEN_2245; // @[lut_35.scala 2474:105 lut_35.scala 2509:43]
  wire  _GEN_2435 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] ? 1'h0 : _GEN_2246; // @[lut_35.scala 2474:105 lut_35.scala 2510:43]
  wire  _GEN_2436 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] ? 1'h0 : _GEN_2247; // @[lut_35.scala 2474:105 lut_35.scala 2511:43]
  wire  _GEN_2437 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] | _GEN_2248; // @[lut_35.scala 2474:105 lut_35.scala 2512:38]
  wire  _GEN_2441 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2474:105 lut_35.scala 177:26 lut_35.scala 2514:89]
  wire  _GEN_2449 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] ? 1'h0 : _GEN_2252; // @[lut_35.scala 2474:105 lut_35.scala 177:26]
  wire  _GEN_2457 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] ? 1'h0 : _GEN_2260; // @[lut_35.scala 2474:105 lut_35.scala 177:26]
  wire  _GEN_2465 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] ? 1'h0 : _GEN_2268; // @[lut_35.scala 2474:105 lut_35.scala 177:26]
  wire  _GEN_2473 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] ? 1'h0 : _GEN_2276; // @[lut_35.scala 2474:105 lut_35.scala 177:26]
  wire  _GEN_2481 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] ? 1'h0 : _GEN_2284; // @[lut_35.scala 2474:105 lut_35.scala 177:26]
  wire  _GEN_2489 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] ? 1'h0 : _GEN_2292; // @[lut_35.scala 2474:105 lut_35.scala 177:26]
  wire  _GEN_2497 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] ? 1'h0 : _GEN_2300; // @[lut_35.scala 2474:105 lut_35.scala 177:26]
  wire  _GEN_2505 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] ? 1'h0 : _GEN_2308; // @[lut_35.scala 2474:105 lut_35.scala 177:26]
  wire  _GEN_2513 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] ? 1'h0 : _GEN_2316; // @[lut_35.scala 2474:105 lut_35.scala 177:26]
  wire  _GEN_2521 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] ? 1'h0 : _GEN_2324; // @[lut_35.scala 2474:105 lut_35.scala 177:26]
  wire  _GEN_2529 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] ? 1'h0 : _GEN_2332; // @[lut_35.scala 2474:105 lut_35.scala 177:26]
  wire  _GEN_2537 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] ? 1'h0 : _GEN_2340; // @[lut_35.scala 2474:105 lut_35.scala 177:26]
  wire  _GEN_2545 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] ? 1'h0 : _GEN_2348; // @[lut_35.scala 2474:105 lut_35.scala 177:26]
  wire  _GEN_2553 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] ? 1'h0 : _GEN_2356; // @[lut_35.scala 2474:105 lut_35.scala 177:26]
  wire  _GEN_2561 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] ? 1'h0 : _GEN_2364; // @[lut_35.scala 2474:105 lut_35.scala 177:26]
  wire  _GEN_2569 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] ? 1'h0 : _GEN_2372; // @[lut_35.scala 2474:105 lut_35.scala 177:26]
  wire  _GEN_2577 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] ? 1'h0 : _GEN_2380; // @[lut_35.scala 2474:105 lut_35.scala 177:26]
  wire  _GEN_2585 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] ? 1'h0 : _GEN_2388; // @[lut_35.scala 2474:105 lut_35.scala 177:26]
  wire  _GEN_2593 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] ? 1'h0 : _GEN_2396; // @[lut_35.scala 2474:105 lut_35.scala 177:26]
  wire  _GEN_2601 = io_empty_13 & push_valid & ~push_13_1 & ~LUT_mem_MPORT_236_data[32] ? 1'h0 : _GEN_2404; // @[lut_35.scala 2474:105 lut_35.scala 177:26]
  wire  _GEN_2613 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _T_445; // @[lut_35.scala 2434:105 lut_35.scala 2450:43]
  wire  _GEN_2614 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _GEN_2416; // @[lut_35.scala 2434:105 lut_35.scala 2451:43]
  wire  _GEN_2615 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _GEN_2417; // @[lut_35.scala 2434:105 lut_35.scala 2452:43]
  wire  _GEN_2616 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _GEN_2418; // @[lut_35.scala 2434:105 lut_35.scala 2453:43]
  wire  _GEN_2617 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _GEN_2419; // @[lut_35.scala 2434:105 lut_35.scala 2454:43]
  wire  _GEN_2618 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _GEN_2420; // @[lut_35.scala 2434:105 lut_35.scala 2455:43]
  wire  _GEN_2619 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _GEN_2421; // @[lut_35.scala 2434:105 lut_35.scala 2456:43]
  wire  _GEN_2620 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _GEN_2422; // @[lut_35.scala 2434:105 lut_35.scala 2457:43]
  wire  _GEN_2621 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _GEN_2423; // @[lut_35.scala 2434:105 lut_35.scala 2458:43]
  wire  _GEN_2622 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _GEN_2424; // @[lut_35.scala 2434:105 lut_35.scala 2459:43]
  wire  _GEN_2623 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _GEN_2425; // @[lut_35.scala 2434:105 lut_35.scala 2460:43]
  wire  _GEN_2624 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _GEN_2426; // @[lut_35.scala 2434:105 lut_35.scala 2461:43]
  wire  _GEN_2625 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _GEN_2427; // @[lut_35.scala 2434:105 lut_35.scala 2462:43]
  wire  _GEN_2626 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _GEN_2428; // @[lut_35.scala 2434:105 lut_35.scala 2463:43]
  wire  _GEN_2627 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _GEN_2429; // @[lut_35.scala 2434:105 lut_35.scala 2464:43]
  wire  _GEN_2628 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _GEN_2430; // @[lut_35.scala 2434:105 lut_35.scala 2465:43]
  wire  _GEN_2629 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _GEN_2431; // @[lut_35.scala 2434:105 lut_35.scala 2466:43]
  wire  _GEN_2630 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _GEN_2432; // @[lut_35.scala 2434:105 lut_35.scala 2467:43]
  wire  _GEN_2631 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _GEN_2433; // @[lut_35.scala 2434:105 lut_35.scala 2468:43]
  wire  _GEN_2632 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _GEN_2434; // @[lut_35.scala 2434:105 lut_35.scala 2469:43]
  wire  _GEN_2633 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _GEN_2435; // @[lut_35.scala 2434:105 lut_35.scala 2470:43]
  wire  _GEN_2634 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _GEN_2436; // @[lut_35.scala 2434:105 lut_35.scala 2471:43]
  wire  _GEN_2635 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] | _GEN_2437; // @[lut_35.scala 2434:105 lut_35.scala 2472:38]
  wire  _GEN_2639 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2434:105 lut_35.scala 177:26 lut_35.scala 2474:89]
  wire  _GEN_2647 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _GEN_2441; // @[lut_35.scala 2434:105 lut_35.scala 177:26]
  wire  _GEN_2655 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _GEN_2449; // @[lut_35.scala 2434:105 lut_35.scala 177:26]
  wire  _GEN_2663 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _GEN_2457; // @[lut_35.scala 2434:105 lut_35.scala 177:26]
  wire  _GEN_2671 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _GEN_2465; // @[lut_35.scala 2434:105 lut_35.scala 177:26]
  wire  _GEN_2679 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _GEN_2473; // @[lut_35.scala 2434:105 lut_35.scala 177:26]
  wire  _GEN_2687 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _GEN_2481; // @[lut_35.scala 2434:105 lut_35.scala 177:26]
  wire  _GEN_2695 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _GEN_2489; // @[lut_35.scala 2434:105 lut_35.scala 177:26]
  wire  _GEN_2703 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _GEN_2497; // @[lut_35.scala 2434:105 lut_35.scala 177:26]
  wire  _GEN_2711 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _GEN_2505; // @[lut_35.scala 2434:105 lut_35.scala 177:26]
  wire  _GEN_2719 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _GEN_2513; // @[lut_35.scala 2434:105 lut_35.scala 177:26]
  wire  _GEN_2727 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _GEN_2521; // @[lut_35.scala 2434:105 lut_35.scala 177:26]
  wire  _GEN_2735 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _GEN_2529; // @[lut_35.scala 2434:105 lut_35.scala 177:26]
  wire  _GEN_2743 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _GEN_2537; // @[lut_35.scala 2434:105 lut_35.scala 177:26]
  wire  _GEN_2751 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _GEN_2545; // @[lut_35.scala 2434:105 lut_35.scala 177:26]
  wire  _GEN_2759 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _GEN_2553; // @[lut_35.scala 2434:105 lut_35.scala 177:26]
  wire  _GEN_2767 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _GEN_2561; // @[lut_35.scala 2434:105 lut_35.scala 177:26]
  wire  _GEN_2775 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _GEN_2569; // @[lut_35.scala 2434:105 lut_35.scala 177:26]
  wire  _GEN_2783 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _GEN_2577; // @[lut_35.scala 2434:105 lut_35.scala 177:26]
  wire  _GEN_2791 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _GEN_2585; // @[lut_35.scala 2434:105 lut_35.scala 177:26]
  wire  _GEN_2799 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _GEN_2593; // @[lut_35.scala 2434:105 lut_35.scala 177:26]
  wire  _GEN_2807 = io_empty_12 & push_valid & ~push_12_1 & ~LUT_mem_MPORT_234_data[32] ? 1'h0 : _GEN_2601; // @[lut_35.scala 2434:105 lut_35.scala 177:26]
  wire  _GEN_2819 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _T_436; // @[lut_35.scala 2394:105 lut_35.scala 2409:43]
  wire  _GEN_2820 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2613; // @[lut_35.scala 2394:105 lut_35.scala 2410:43]
  wire  _GEN_2821 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2614; // @[lut_35.scala 2394:105 lut_35.scala 2411:43]
  wire  _GEN_2822 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2615; // @[lut_35.scala 2394:105 lut_35.scala 2412:43]
  wire  _GEN_2823 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2616; // @[lut_35.scala 2394:105 lut_35.scala 2413:43]
  wire  _GEN_2824 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2617; // @[lut_35.scala 2394:105 lut_35.scala 2414:43]
  wire  _GEN_2825 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2618; // @[lut_35.scala 2394:105 lut_35.scala 2415:43]
  wire  _GEN_2826 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2619; // @[lut_35.scala 2394:105 lut_35.scala 2416:43]
  wire  _GEN_2827 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2620; // @[lut_35.scala 2394:105 lut_35.scala 2417:43]
  wire  _GEN_2828 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2621; // @[lut_35.scala 2394:105 lut_35.scala 2418:43]
  wire  _GEN_2829 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2622; // @[lut_35.scala 2394:105 lut_35.scala 2419:43]
  wire  _GEN_2830 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2623; // @[lut_35.scala 2394:105 lut_35.scala 2420:43]
  wire  _GEN_2831 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2624; // @[lut_35.scala 2394:105 lut_35.scala 2421:43]
  wire  _GEN_2832 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2625; // @[lut_35.scala 2394:105 lut_35.scala 2422:43]
  wire  _GEN_2833 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2626; // @[lut_35.scala 2394:105 lut_35.scala 2423:43]
  wire  _GEN_2834 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2627; // @[lut_35.scala 2394:105 lut_35.scala 2424:43]
  wire  _GEN_2835 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2628; // @[lut_35.scala 2394:105 lut_35.scala 2425:43]
  wire  _GEN_2836 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2629; // @[lut_35.scala 2394:105 lut_35.scala 2426:43]
  wire  _GEN_2837 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2630; // @[lut_35.scala 2394:105 lut_35.scala 2427:43]
  wire  _GEN_2838 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2631; // @[lut_35.scala 2394:105 lut_35.scala 2428:43]
  wire  _GEN_2839 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2632; // @[lut_35.scala 2394:105 lut_35.scala 2429:43]
  wire  _GEN_2840 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2633; // @[lut_35.scala 2394:105 lut_35.scala 2430:43]
  wire  _GEN_2841 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2634; // @[lut_35.scala 2394:105 lut_35.scala 2431:43]
  wire  _GEN_2842 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] | _GEN_2635; // @[lut_35.scala 2394:105 lut_35.scala 2432:38]
  wire  _GEN_2846 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2394:105 lut_35.scala 177:26 lut_35.scala 2434:89]
  wire  _GEN_2854 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2639; // @[lut_35.scala 2394:105 lut_35.scala 177:26]
  wire  _GEN_2862 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2647; // @[lut_35.scala 2394:105 lut_35.scala 177:26]
  wire  _GEN_2870 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2655; // @[lut_35.scala 2394:105 lut_35.scala 177:26]
  wire  _GEN_2878 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2663; // @[lut_35.scala 2394:105 lut_35.scala 177:26]
  wire  _GEN_2886 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2671; // @[lut_35.scala 2394:105 lut_35.scala 177:26]
  wire  _GEN_2894 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2679; // @[lut_35.scala 2394:105 lut_35.scala 177:26]
  wire  _GEN_2902 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2687; // @[lut_35.scala 2394:105 lut_35.scala 177:26]
  wire  _GEN_2910 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2695; // @[lut_35.scala 2394:105 lut_35.scala 177:26]
  wire  _GEN_2918 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2703; // @[lut_35.scala 2394:105 lut_35.scala 177:26]
  wire  _GEN_2926 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2711; // @[lut_35.scala 2394:105 lut_35.scala 177:26]
  wire  _GEN_2934 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2719; // @[lut_35.scala 2394:105 lut_35.scala 177:26]
  wire  _GEN_2942 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2727; // @[lut_35.scala 2394:105 lut_35.scala 177:26]
  wire  _GEN_2950 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2735; // @[lut_35.scala 2394:105 lut_35.scala 177:26]
  wire  _GEN_2958 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2743; // @[lut_35.scala 2394:105 lut_35.scala 177:26]
  wire  _GEN_2966 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2751; // @[lut_35.scala 2394:105 lut_35.scala 177:26]
  wire  _GEN_2974 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2759; // @[lut_35.scala 2394:105 lut_35.scala 177:26]
  wire  _GEN_2982 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2767; // @[lut_35.scala 2394:105 lut_35.scala 177:26]
  wire  _GEN_2990 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2775; // @[lut_35.scala 2394:105 lut_35.scala 177:26]
  wire  _GEN_2998 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2783; // @[lut_35.scala 2394:105 lut_35.scala 177:26]
  wire  _GEN_3006 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2791; // @[lut_35.scala 2394:105 lut_35.scala 177:26]
  wire  _GEN_3014 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2799; // @[lut_35.scala 2394:105 lut_35.scala 177:26]
  wire  _GEN_3022 = io_empty_11 & push_valid & ~push_11_1 & ~LUT_mem_MPORT_232_data[32] ? 1'h0 : _GEN_2807; // @[lut_35.scala 2394:105 lut_35.scala 177:26]
  wire  _GEN_3034 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _T_427; // @[lut_35.scala 2354:105 lut_35.scala 2368:43]
  wire  _GEN_3035 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2819; // @[lut_35.scala 2354:105 lut_35.scala 2369:43]
  wire  _GEN_3036 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2820; // @[lut_35.scala 2354:105 lut_35.scala 2370:43]
  wire  _GEN_3037 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2821; // @[lut_35.scala 2354:105 lut_35.scala 2371:43]
  wire  _GEN_3038 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2822; // @[lut_35.scala 2354:105 lut_35.scala 2372:43]
  wire  _GEN_3039 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2823; // @[lut_35.scala 2354:105 lut_35.scala 2373:43]
  wire  _GEN_3040 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2824; // @[lut_35.scala 2354:105 lut_35.scala 2374:43]
  wire  _GEN_3041 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2825; // @[lut_35.scala 2354:105 lut_35.scala 2375:43]
  wire  _GEN_3042 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2826; // @[lut_35.scala 2354:105 lut_35.scala 2376:43]
  wire  _GEN_3043 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2827; // @[lut_35.scala 2354:105 lut_35.scala 2377:43]
  wire  _GEN_3044 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2828; // @[lut_35.scala 2354:105 lut_35.scala 2378:43]
  wire  _GEN_3045 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2829; // @[lut_35.scala 2354:105 lut_35.scala 2379:43]
  wire  _GEN_3046 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2830; // @[lut_35.scala 2354:105 lut_35.scala 2380:43]
  wire  _GEN_3047 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2831; // @[lut_35.scala 2354:105 lut_35.scala 2381:43]
  wire  _GEN_3048 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2832; // @[lut_35.scala 2354:105 lut_35.scala 2382:43]
  wire  _GEN_3049 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2833; // @[lut_35.scala 2354:105 lut_35.scala 2383:43]
  wire  _GEN_3050 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2834; // @[lut_35.scala 2354:105 lut_35.scala 2384:43]
  wire  _GEN_3051 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2835; // @[lut_35.scala 2354:105 lut_35.scala 2385:43]
  wire  _GEN_3052 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2836; // @[lut_35.scala 2354:105 lut_35.scala 2386:43]
  wire  _GEN_3053 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2837; // @[lut_35.scala 2354:105 lut_35.scala 2387:43]
  wire  _GEN_3054 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2838; // @[lut_35.scala 2354:105 lut_35.scala 2388:43]
  wire  _GEN_3055 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2839; // @[lut_35.scala 2354:105 lut_35.scala 2389:43]
  wire  _GEN_3056 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2840; // @[lut_35.scala 2354:105 lut_35.scala 2390:43]
  wire  _GEN_3057 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2841; // @[lut_35.scala 2354:105 lut_35.scala 2391:43]
  wire  _GEN_3058 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] | _GEN_2842; // @[lut_35.scala 2354:105 lut_35.scala 2392:38]
  wire  _GEN_3062 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2354:105 lut_35.scala 177:26 lut_35.scala 2394:89]
  wire  _GEN_3070 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2846; // @[lut_35.scala 2354:105 lut_35.scala 177:26]
  wire  _GEN_3078 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2854; // @[lut_35.scala 2354:105 lut_35.scala 177:26]
  wire  _GEN_3086 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2862; // @[lut_35.scala 2354:105 lut_35.scala 177:26]
  wire  _GEN_3094 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2870; // @[lut_35.scala 2354:105 lut_35.scala 177:26]
  wire  _GEN_3102 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2878; // @[lut_35.scala 2354:105 lut_35.scala 177:26]
  wire  _GEN_3110 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2886; // @[lut_35.scala 2354:105 lut_35.scala 177:26]
  wire  _GEN_3118 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2894; // @[lut_35.scala 2354:105 lut_35.scala 177:26]
  wire  _GEN_3126 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2902; // @[lut_35.scala 2354:105 lut_35.scala 177:26]
  wire  _GEN_3134 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2910; // @[lut_35.scala 2354:105 lut_35.scala 177:26]
  wire  _GEN_3142 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2918; // @[lut_35.scala 2354:105 lut_35.scala 177:26]
  wire  _GEN_3150 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2926; // @[lut_35.scala 2354:105 lut_35.scala 177:26]
  wire  _GEN_3158 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2934; // @[lut_35.scala 2354:105 lut_35.scala 177:26]
  wire  _GEN_3166 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2942; // @[lut_35.scala 2354:105 lut_35.scala 177:26]
  wire  _GEN_3174 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2950; // @[lut_35.scala 2354:105 lut_35.scala 177:26]
  wire  _GEN_3182 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2958; // @[lut_35.scala 2354:105 lut_35.scala 177:26]
  wire  _GEN_3190 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2966; // @[lut_35.scala 2354:105 lut_35.scala 177:26]
  wire  _GEN_3198 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2974; // @[lut_35.scala 2354:105 lut_35.scala 177:26]
  wire  _GEN_3206 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2982; // @[lut_35.scala 2354:105 lut_35.scala 177:26]
  wire  _GEN_3214 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2990; // @[lut_35.scala 2354:105 lut_35.scala 177:26]
  wire  _GEN_3222 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_2998; // @[lut_35.scala 2354:105 lut_35.scala 177:26]
  wire  _GEN_3230 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_3006; // @[lut_35.scala 2354:105 lut_35.scala 177:26]
  wire  _GEN_3238 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_3014; // @[lut_35.scala 2354:105 lut_35.scala 177:26]
  wire  _GEN_3246 = io_empty_10 & push_valid & ~push_10_1 & ~LUT_mem_MPORT_230_data[32] ? 1'h0 : _GEN_3022; // @[lut_35.scala 2354:105 lut_35.scala 177:26]
  wire  _GEN_3258 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _T_418; // @[lut_35.scala 2314:102 lut_35.scala 2327:43]
  wire  _GEN_3259 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3034; // @[lut_35.scala 2314:102 lut_35.scala 2328:43]
  wire  _GEN_3260 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3035; // @[lut_35.scala 2314:102 lut_35.scala 2329:43]
  wire  _GEN_3261 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3036; // @[lut_35.scala 2314:102 lut_35.scala 2330:43]
  wire  _GEN_3262 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3037; // @[lut_35.scala 2314:102 lut_35.scala 2331:43]
  wire  _GEN_3263 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3038; // @[lut_35.scala 2314:102 lut_35.scala 2332:43]
  wire  _GEN_3264 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3039; // @[lut_35.scala 2314:102 lut_35.scala 2333:43]
  wire  _GEN_3265 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3040; // @[lut_35.scala 2314:102 lut_35.scala 2334:43]
  wire  _GEN_3266 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3041; // @[lut_35.scala 2314:102 lut_35.scala 2335:43]
  wire  _GEN_3267 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3042; // @[lut_35.scala 2314:102 lut_35.scala 2336:43]
  wire  _GEN_3268 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3043; // @[lut_35.scala 2314:102 lut_35.scala 2337:43]
  wire  _GEN_3269 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3044; // @[lut_35.scala 2314:102 lut_35.scala 2338:43]
  wire  _GEN_3270 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3045; // @[lut_35.scala 2314:102 lut_35.scala 2339:43]
  wire  _GEN_3271 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3046; // @[lut_35.scala 2314:102 lut_35.scala 2340:43]
  wire  _GEN_3272 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3047; // @[lut_35.scala 2314:102 lut_35.scala 2341:43]
  wire  _GEN_3273 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3048; // @[lut_35.scala 2314:102 lut_35.scala 2342:43]
  wire  _GEN_3274 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3049; // @[lut_35.scala 2314:102 lut_35.scala 2343:43]
  wire  _GEN_3275 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3050; // @[lut_35.scala 2314:102 lut_35.scala 2344:43]
  wire  _GEN_3276 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3051; // @[lut_35.scala 2314:102 lut_35.scala 2345:43]
  wire  _GEN_3277 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3052; // @[lut_35.scala 2314:102 lut_35.scala 2346:43]
  wire  _GEN_3278 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3053; // @[lut_35.scala 2314:102 lut_35.scala 2347:43]
  wire  _GEN_3279 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3054; // @[lut_35.scala 2314:102 lut_35.scala 2348:43]
  wire  _GEN_3280 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3055; // @[lut_35.scala 2314:102 lut_35.scala 2349:43]
  wire  _GEN_3281 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3056; // @[lut_35.scala 2314:102 lut_35.scala 2350:43]
  wire  _GEN_3282 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3057; // @[lut_35.scala 2314:102 lut_35.scala 2351:43]
  wire  _GEN_3283 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] | _GEN_3058; // @[lut_35.scala 2314:102 lut_35.scala 2352:38]
  wire  _GEN_3287 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2314:102 lut_35.scala 177:26 lut_35.scala 2354:89]
  wire  _GEN_3295 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3062; // @[lut_35.scala 2314:102 lut_35.scala 177:26]
  wire  _GEN_3303 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3070; // @[lut_35.scala 2314:102 lut_35.scala 177:26]
  wire  _GEN_3311 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3078; // @[lut_35.scala 2314:102 lut_35.scala 177:26]
  wire  _GEN_3319 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3086; // @[lut_35.scala 2314:102 lut_35.scala 177:26]
  wire  _GEN_3327 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3094; // @[lut_35.scala 2314:102 lut_35.scala 177:26]
  wire  _GEN_3335 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3102; // @[lut_35.scala 2314:102 lut_35.scala 177:26]
  wire  _GEN_3343 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3110; // @[lut_35.scala 2314:102 lut_35.scala 177:26]
  wire  _GEN_3351 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3118; // @[lut_35.scala 2314:102 lut_35.scala 177:26]
  wire  _GEN_3359 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3126; // @[lut_35.scala 2314:102 lut_35.scala 177:26]
  wire  _GEN_3367 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3134; // @[lut_35.scala 2314:102 lut_35.scala 177:26]
  wire  _GEN_3375 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3142; // @[lut_35.scala 2314:102 lut_35.scala 177:26]
  wire  _GEN_3383 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3150; // @[lut_35.scala 2314:102 lut_35.scala 177:26]
  wire  _GEN_3391 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3158; // @[lut_35.scala 2314:102 lut_35.scala 177:26]
  wire  _GEN_3399 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3166; // @[lut_35.scala 2314:102 lut_35.scala 177:26]
  wire  _GEN_3407 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3174; // @[lut_35.scala 2314:102 lut_35.scala 177:26]
  wire  _GEN_3415 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3182; // @[lut_35.scala 2314:102 lut_35.scala 177:26]
  wire  _GEN_3423 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3190; // @[lut_35.scala 2314:102 lut_35.scala 177:26]
  wire  _GEN_3431 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3198; // @[lut_35.scala 2314:102 lut_35.scala 177:26]
  wire  _GEN_3439 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3206; // @[lut_35.scala 2314:102 lut_35.scala 177:26]
  wire  _GEN_3447 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3214; // @[lut_35.scala 2314:102 lut_35.scala 177:26]
  wire  _GEN_3455 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3222; // @[lut_35.scala 2314:102 lut_35.scala 177:26]
  wire  _GEN_3463 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3230; // @[lut_35.scala 2314:102 lut_35.scala 177:26]
  wire  _GEN_3471 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3238; // @[lut_35.scala 2314:102 lut_35.scala 177:26]
  wire  _GEN_3479 = io_empty_9 & push_valid & ~push_9_1 & ~LUT_mem_MPORT_228_data[32] ? 1'h0 : _GEN_3246; // @[lut_35.scala 2314:102 lut_35.scala 177:26]
  wire  _GEN_3491 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _T_409; // @[lut_35.scala 2274:102 lut_35.scala 2286:42]
  wire  _GEN_3492 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3258; // @[lut_35.scala 2274:102 lut_35.scala 2287:43]
  wire  _GEN_3493 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3259; // @[lut_35.scala 2274:102 lut_35.scala 2288:43]
  wire  _GEN_3494 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3260; // @[lut_35.scala 2274:102 lut_35.scala 2289:43]
  wire  _GEN_3495 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3261; // @[lut_35.scala 2274:102 lut_35.scala 2290:43]
  wire  _GEN_3496 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3262; // @[lut_35.scala 2274:102 lut_35.scala 2291:43]
  wire  _GEN_3497 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3263; // @[lut_35.scala 2274:102 lut_35.scala 2292:43]
  wire  _GEN_3498 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3264; // @[lut_35.scala 2274:102 lut_35.scala 2293:43]
  wire  _GEN_3499 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3265; // @[lut_35.scala 2274:102 lut_35.scala 2294:43]
  wire  _GEN_3500 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3266; // @[lut_35.scala 2274:102 lut_35.scala 2295:43]
  wire  _GEN_3501 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3267; // @[lut_35.scala 2274:102 lut_35.scala 2296:43]
  wire  _GEN_3502 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3268; // @[lut_35.scala 2274:102 lut_35.scala 2297:43]
  wire  _GEN_3503 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3269; // @[lut_35.scala 2274:102 lut_35.scala 2298:43]
  wire  _GEN_3504 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3270; // @[lut_35.scala 2274:102 lut_35.scala 2299:43]
  wire  _GEN_3505 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3271; // @[lut_35.scala 2274:102 lut_35.scala 2300:43]
  wire  _GEN_3506 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3272; // @[lut_35.scala 2274:102 lut_35.scala 2301:43]
  wire  _GEN_3507 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3273; // @[lut_35.scala 2274:102 lut_35.scala 2302:43]
  wire  _GEN_3508 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3274; // @[lut_35.scala 2274:102 lut_35.scala 2303:43]
  wire  _GEN_3509 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3275; // @[lut_35.scala 2274:102 lut_35.scala 2304:43]
  wire  _GEN_3510 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3276; // @[lut_35.scala 2274:102 lut_35.scala 2305:43]
  wire  _GEN_3511 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3277; // @[lut_35.scala 2274:102 lut_35.scala 2306:43]
  wire  _GEN_3512 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3278; // @[lut_35.scala 2274:102 lut_35.scala 2307:43]
  wire  _GEN_3513 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3279; // @[lut_35.scala 2274:102 lut_35.scala 2308:43]
  wire  _GEN_3514 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3280; // @[lut_35.scala 2274:102 lut_35.scala 2309:43]
  wire  _GEN_3515 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3281; // @[lut_35.scala 2274:102 lut_35.scala 2310:43]
  wire  _GEN_3516 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3282; // @[lut_35.scala 2274:102 lut_35.scala 2311:43]
  wire  _GEN_3517 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] | _GEN_3283; // @[lut_35.scala 2274:102 lut_35.scala 2312:38]
  wire  _GEN_3521 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2274:102 lut_35.scala 177:26 lut_35.scala 2314:87]
  wire  _GEN_3529 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3287; // @[lut_35.scala 2274:102 lut_35.scala 177:26]
  wire  _GEN_3537 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3295; // @[lut_35.scala 2274:102 lut_35.scala 177:26]
  wire  _GEN_3545 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3303; // @[lut_35.scala 2274:102 lut_35.scala 177:26]
  wire  _GEN_3553 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3311; // @[lut_35.scala 2274:102 lut_35.scala 177:26]
  wire  _GEN_3561 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3319; // @[lut_35.scala 2274:102 lut_35.scala 177:26]
  wire  _GEN_3569 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3327; // @[lut_35.scala 2274:102 lut_35.scala 177:26]
  wire  _GEN_3577 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3335; // @[lut_35.scala 2274:102 lut_35.scala 177:26]
  wire  _GEN_3585 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3343; // @[lut_35.scala 2274:102 lut_35.scala 177:26]
  wire  _GEN_3593 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3351; // @[lut_35.scala 2274:102 lut_35.scala 177:26]
  wire  _GEN_3601 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3359; // @[lut_35.scala 2274:102 lut_35.scala 177:26]
  wire  _GEN_3609 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3367; // @[lut_35.scala 2274:102 lut_35.scala 177:26]
  wire  _GEN_3617 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3375; // @[lut_35.scala 2274:102 lut_35.scala 177:26]
  wire  _GEN_3625 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3383; // @[lut_35.scala 2274:102 lut_35.scala 177:26]
  wire  _GEN_3633 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3391; // @[lut_35.scala 2274:102 lut_35.scala 177:26]
  wire  _GEN_3641 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3399; // @[lut_35.scala 2274:102 lut_35.scala 177:26]
  wire  _GEN_3649 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3407; // @[lut_35.scala 2274:102 lut_35.scala 177:26]
  wire  _GEN_3657 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3415; // @[lut_35.scala 2274:102 lut_35.scala 177:26]
  wire  _GEN_3665 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3423; // @[lut_35.scala 2274:102 lut_35.scala 177:26]
  wire  _GEN_3673 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3431; // @[lut_35.scala 2274:102 lut_35.scala 177:26]
  wire  _GEN_3681 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3439; // @[lut_35.scala 2274:102 lut_35.scala 177:26]
  wire  _GEN_3689 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3447; // @[lut_35.scala 2274:102 lut_35.scala 177:26]
  wire  _GEN_3697 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3455; // @[lut_35.scala 2274:102 lut_35.scala 177:26]
  wire  _GEN_3705 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3463; // @[lut_35.scala 2274:102 lut_35.scala 177:26]
  wire  _GEN_3713 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3471; // @[lut_35.scala 2274:102 lut_35.scala 177:26]
  wire  _GEN_3721 = io_empty_8 & push_valid & ~push_8_1 & ~LUT_mem_MPORT_226_data[32] ? 1'h0 : _GEN_3479; // @[lut_35.scala 2274:102 lut_35.scala 177:26]
  wire  _GEN_3733 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _T_400; // @[lut_35.scala 2234:102 lut_35.scala 2245:42]
  wire  _GEN_3734 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3491; // @[lut_35.scala 2234:102 lut_35.scala 2246:42]
  wire  _GEN_3735 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3492; // @[lut_35.scala 2234:102 lut_35.scala 2247:43]
  wire  _GEN_3736 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3493; // @[lut_35.scala 2234:102 lut_35.scala 2248:43]
  wire  _GEN_3737 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3494; // @[lut_35.scala 2234:102 lut_35.scala 2249:43]
  wire  _GEN_3738 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3495; // @[lut_35.scala 2234:102 lut_35.scala 2250:43]
  wire  _GEN_3739 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3496; // @[lut_35.scala 2234:102 lut_35.scala 2251:43]
  wire  _GEN_3740 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3497; // @[lut_35.scala 2234:102 lut_35.scala 2252:43]
  wire  _GEN_3741 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3498; // @[lut_35.scala 2234:102 lut_35.scala 2253:43]
  wire  _GEN_3742 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3499; // @[lut_35.scala 2234:102 lut_35.scala 2254:43]
  wire  _GEN_3743 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3500; // @[lut_35.scala 2234:102 lut_35.scala 2255:43]
  wire  _GEN_3744 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3501; // @[lut_35.scala 2234:102 lut_35.scala 2256:43]
  wire  _GEN_3745 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3502; // @[lut_35.scala 2234:102 lut_35.scala 2257:43]
  wire  _GEN_3746 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3503; // @[lut_35.scala 2234:102 lut_35.scala 2258:43]
  wire  _GEN_3747 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3504; // @[lut_35.scala 2234:102 lut_35.scala 2259:43]
  wire  _GEN_3748 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3505; // @[lut_35.scala 2234:102 lut_35.scala 2260:43]
  wire  _GEN_3749 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3506; // @[lut_35.scala 2234:102 lut_35.scala 2261:43]
  wire  _GEN_3750 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3507; // @[lut_35.scala 2234:102 lut_35.scala 2262:43]
  wire  _GEN_3751 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3508; // @[lut_35.scala 2234:102 lut_35.scala 2263:43]
  wire  _GEN_3752 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3509; // @[lut_35.scala 2234:102 lut_35.scala 2264:43]
  wire  _GEN_3753 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3510; // @[lut_35.scala 2234:102 lut_35.scala 2265:43]
  wire  _GEN_3754 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3511; // @[lut_35.scala 2234:102 lut_35.scala 2266:43]
  wire  _GEN_3755 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3512; // @[lut_35.scala 2234:102 lut_35.scala 2267:43]
  wire  _GEN_3756 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3513; // @[lut_35.scala 2234:102 lut_35.scala 2268:43]
  wire  _GEN_3757 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3514; // @[lut_35.scala 2234:102 lut_35.scala 2269:43]
  wire  _GEN_3758 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3515; // @[lut_35.scala 2234:102 lut_35.scala 2270:43]
  wire  _GEN_3759 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3516; // @[lut_35.scala 2234:102 lut_35.scala 2271:43]
  wire  _GEN_3760 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] | _GEN_3517; // @[lut_35.scala 2234:102 lut_35.scala 2272:38]
  wire  _GEN_3764 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2234:102 lut_35.scala 177:26 lut_35.scala 2274:87]
  wire  _GEN_3772 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3521; // @[lut_35.scala 2234:102 lut_35.scala 177:26]
  wire  _GEN_3780 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3529; // @[lut_35.scala 2234:102 lut_35.scala 177:26]
  wire  _GEN_3788 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3537; // @[lut_35.scala 2234:102 lut_35.scala 177:26]
  wire  _GEN_3796 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3545; // @[lut_35.scala 2234:102 lut_35.scala 177:26]
  wire  _GEN_3804 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3553; // @[lut_35.scala 2234:102 lut_35.scala 177:26]
  wire  _GEN_3812 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3561; // @[lut_35.scala 2234:102 lut_35.scala 177:26]
  wire  _GEN_3820 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3569; // @[lut_35.scala 2234:102 lut_35.scala 177:26]
  wire  _GEN_3828 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3577; // @[lut_35.scala 2234:102 lut_35.scala 177:26]
  wire  _GEN_3836 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3585; // @[lut_35.scala 2234:102 lut_35.scala 177:26]
  wire  _GEN_3844 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3593; // @[lut_35.scala 2234:102 lut_35.scala 177:26]
  wire  _GEN_3852 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3601; // @[lut_35.scala 2234:102 lut_35.scala 177:26]
  wire  _GEN_3860 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3609; // @[lut_35.scala 2234:102 lut_35.scala 177:26]
  wire  _GEN_3868 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3617; // @[lut_35.scala 2234:102 lut_35.scala 177:26]
  wire  _GEN_3876 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3625; // @[lut_35.scala 2234:102 lut_35.scala 177:26]
  wire  _GEN_3884 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3633; // @[lut_35.scala 2234:102 lut_35.scala 177:26]
  wire  _GEN_3892 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3641; // @[lut_35.scala 2234:102 lut_35.scala 177:26]
  wire  _GEN_3900 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3649; // @[lut_35.scala 2234:102 lut_35.scala 177:26]
  wire  _GEN_3908 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3657; // @[lut_35.scala 2234:102 lut_35.scala 177:26]
  wire  _GEN_3916 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3665; // @[lut_35.scala 2234:102 lut_35.scala 177:26]
  wire  _GEN_3924 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3673; // @[lut_35.scala 2234:102 lut_35.scala 177:26]
  wire  _GEN_3932 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3681; // @[lut_35.scala 2234:102 lut_35.scala 177:26]
  wire  _GEN_3940 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3689; // @[lut_35.scala 2234:102 lut_35.scala 177:26]
  wire  _GEN_3948 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3697; // @[lut_35.scala 2234:102 lut_35.scala 177:26]
  wire  _GEN_3956 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3705; // @[lut_35.scala 2234:102 lut_35.scala 177:26]
  wire  _GEN_3964 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3713; // @[lut_35.scala 2234:102 lut_35.scala 177:26]
  wire  _GEN_3972 = io_empty_7 & push_valid & ~push_7_1 & ~LUT_mem_MPORT_224_data[32] ? 1'h0 : _GEN_3721; // @[lut_35.scala 2234:102 lut_35.scala 177:26]
  wire  _GEN_3984 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _T_391; // @[lut_35.scala 2194:102 lut_35.scala 2204:42]
  wire  _GEN_3985 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3733; // @[lut_35.scala 2194:102 lut_35.scala 2205:42]
  wire  _GEN_3986 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3734; // @[lut_35.scala 2194:102 lut_35.scala 2206:42]
  wire  _GEN_3987 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3735; // @[lut_35.scala 2194:102 lut_35.scala 2207:43]
  wire  _GEN_3988 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3736; // @[lut_35.scala 2194:102 lut_35.scala 2208:43]
  wire  _GEN_3989 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3737; // @[lut_35.scala 2194:102 lut_35.scala 2209:43]
  wire  _GEN_3990 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3738; // @[lut_35.scala 2194:102 lut_35.scala 2210:43]
  wire  _GEN_3991 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3739; // @[lut_35.scala 2194:102 lut_35.scala 2211:43]
  wire  _GEN_3992 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3740; // @[lut_35.scala 2194:102 lut_35.scala 2212:43]
  wire  _GEN_3993 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3741; // @[lut_35.scala 2194:102 lut_35.scala 2213:43]
  wire  _GEN_3994 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3742; // @[lut_35.scala 2194:102 lut_35.scala 2214:43]
  wire  _GEN_3995 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3743; // @[lut_35.scala 2194:102 lut_35.scala 2215:43]
  wire  _GEN_3996 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3744; // @[lut_35.scala 2194:102 lut_35.scala 2216:43]
  wire  _GEN_3997 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3745; // @[lut_35.scala 2194:102 lut_35.scala 2217:43]
  wire  _GEN_3998 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3746; // @[lut_35.scala 2194:102 lut_35.scala 2218:43]
  wire  _GEN_3999 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3747; // @[lut_35.scala 2194:102 lut_35.scala 2219:43]
  wire  _GEN_4000 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3748; // @[lut_35.scala 2194:102 lut_35.scala 2220:43]
  wire  _GEN_4001 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3749; // @[lut_35.scala 2194:102 lut_35.scala 2221:43]
  wire  _GEN_4002 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3750; // @[lut_35.scala 2194:102 lut_35.scala 2222:43]
  wire  _GEN_4003 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3751; // @[lut_35.scala 2194:102 lut_35.scala 2223:43]
  wire  _GEN_4004 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3752; // @[lut_35.scala 2194:102 lut_35.scala 2224:43]
  wire  _GEN_4005 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3753; // @[lut_35.scala 2194:102 lut_35.scala 2225:43]
  wire  _GEN_4006 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3754; // @[lut_35.scala 2194:102 lut_35.scala 2226:43]
  wire  _GEN_4007 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3755; // @[lut_35.scala 2194:102 lut_35.scala 2227:43]
  wire  _GEN_4008 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3756; // @[lut_35.scala 2194:102 lut_35.scala 2228:43]
  wire  _GEN_4009 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3757; // @[lut_35.scala 2194:102 lut_35.scala 2229:43]
  wire  _GEN_4010 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3758; // @[lut_35.scala 2194:102 lut_35.scala 2230:43]
  wire  _GEN_4011 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3759; // @[lut_35.scala 2194:102 lut_35.scala 2231:43]
  wire  _GEN_4012 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] | _GEN_3760; // @[lut_35.scala 2194:102 lut_35.scala 2232:38]
  wire  _GEN_4016 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2194:102 lut_35.scala 177:26 lut_35.scala 2234:87]
  wire  _GEN_4024 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3764; // @[lut_35.scala 2194:102 lut_35.scala 177:26]
  wire  _GEN_4032 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3772; // @[lut_35.scala 2194:102 lut_35.scala 177:26]
  wire  _GEN_4040 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3780; // @[lut_35.scala 2194:102 lut_35.scala 177:26]
  wire  _GEN_4048 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3788; // @[lut_35.scala 2194:102 lut_35.scala 177:26]
  wire  _GEN_4056 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3796; // @[lut_35.scala 2194:102 lut_35.scala 177:26]
  wire  _GEN_4064 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3804; // @[lut_35.scala 2194:102 lut_35.scala 177:26]
  wire  _GEN_4072 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3812; // @[lut_35.scala 2194:102 lut_35.scala 177:26]
  wire  _GEN_4080 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3820; // @[lut_35.scala 2194:102 lut_35.scala 177:26]
  wire  _GEN_4088 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3828; // @[lut_35.scala 2194:102 lut_35.scala 177:26]
  wire  _GEN_4096 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3836; // @[lut_35.scala 2194:102 lut_35.scala 177:26]
  wire  _GEN_4104 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3844; // @[lut_35.scala 2194:102 lut_35.scala 177:26]
  wire  _GEN_4112 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3852; // @[lut_35.scala 2194:102 lut_35.scala 177:26]
  wire  _GEN_4120 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3860; // @[lut_35.scala 2194:102 lut_35.scala 177:26]
  wire  _GEN_4128 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3868; // @[lut_35.scala 2194:102 lut_35.scala 177:26]
  wire  _GEN_4136 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3876; // @[lut_35.scala 2194:102 lut_35.scala 177:26]
  wire  _GEN_4144 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3884; // @[lut_35.scala 2194:102 lut_35.scala 177:26]
  wire  _GEN_4152 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3892; // @[lut_35.scala 2194:102 lut_35.scala 177:26]
  wire  _GEN_4160 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3900; // @[lut_35.scala 2194:102 lut_35.scala 177:26]
  wire  _GEN_4168 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3908; // @[lut_35.scala 2194:102 lut_35.scala 177:26]
  wire  _GEN_4176 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3916; // @[lut_35.scala 2194:102 lut_35.scala 177:26]
  wire  _GEN_4184 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3924; // @[lut_35.scala 2194:102 lut_35.scala 177:26]
  wire  _GEN_4192 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3932; // @[lut_35.scala 2194:102 lut_35.scala 177:26]
  wire  _GEN_4200 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3940; // @[lut_35.scala 2194:102 lut_35.scala 177:26]
  wire  _GEN_4208 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3948; // @[lut_35.scala 2194:102 lut_35.scala 177:26]
  wire  _GEN_4216 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3956; // @[lut_35.scala 2194:102 lut_35.scala 177:26]
  wire  _GEN_4224 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3964; // @[lut_35.scala 2194:102 lut_35.scala 177:26]
  wire  _GEN_4232 = io_empty_6 & push_valid & ~push_6_1 & ~LUT_mem_MPORT_222_data[32] ? 1'h0 : _GEN_3972; // @[lut_35.scala 2194:102 lut_35.scala 177:26]
  wire  _GEN_4244 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _T_382; // @[lut_35.scala 2154:102 lut_35.scala 2163:42]
  wire  _GEN_4245 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_3984; // @[lut_35.scala 2154:102 lut_35.scala 2164:42]
  wire  _GEN_4246 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_3985; // @[lut_35.scala 2154:102 lut_35.scala 2165:42]
  wire  _GEN_4247 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_3986; // @[lut_35.scala 2154:102 lut_35.scala 2166:42]
  wire  _GEN_4248 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_3987; // @[lut_35.scala 2154:102 lut_35.scala 2167:43]
  wire  _GEN_4249 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_3988; // @[lut_35.scala 2154:102 lut_35.scala 2168:43]
  wire  _GEN_4250 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_3989; // @[lut_35.scala 2154:102 lut_35.scala 2169:43]
  wire  _GEN_4251 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_3990; // @[lut_35.scala 2154:102 lut_35.scala 2170:43]
  wire  _GEN_4252 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_3991; // @[lut_35.scala 2154:102 lut_35.scala 2171:43]
  wire  _GEN_4253 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_3992; // @[lut_35.scala 2154:102 lut_35.scala 2172:43]
  wire  _GEN_4254 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_3993; // @[lut_35.scala 2154:102 lut_35.scala 2173:43]
  wire  _GEN_4255 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_3994; // @[lut_35.scala 2154:102 lut_35.scala 2174:43]
  wire  _GEN_4256 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_3995; // @[lut_35.scala 2154:102 lut_35.scala 2175:43]
  wire  _GEN_4257 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_3996; // @[lut_35.scala 2154:102 lut_35.scala 2176:43]
  wire  _GEN_4258 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_3997; // @[lut_35.scala 2154:102 lut_35.scala 2177:43]
  wire  _GEN_4259 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_3998; // @[lut_35.scala 2154:102 lut_35.scala 2178:43]
  wire  _GEN_4260 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_3999; // @[lut_35.scala 2154:102 lut_35.scala 2179:43]
  wire  _GEN_4261 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_4000; // @[lut_35.scala 2154:102 lut_35.scala 2180:43]
  wire  _GEN_4262 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_4001; // @[lut_35.scala 2154:102 lut_35.scala 2181:43]
  wire  _GEN_4263 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_4002; // @[lut_35.scala 2154:102 lut_35.scala 2182:43]
  wire  _GEN_4264 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_4003; // @[lut_35.scala 2154:102 lut_35.scala 2183:43]
  wire  _GEN_4265 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_4004; // @[lut_35.scala 2154:102 lut_35.scala 2184:43]
  wire  _GEN_4266 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_4005; // @[lut_35.scala 2154:102 lut_35.scala 2185:43]
  wire  _GEN_4267 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_4006; // @[lut_35.scala 2154:102 lut_35.scala 2186:43]
  wire  _GEN_4268 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_4007; // @[lut_35.scala 2154:102 lut_35.scala 2187:43]
  wire  _GEN_4269 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_4008; // @[lut_35.scala 2154:102 lut_35.scala 2188:43]
  wire  _GEN_4270 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_4009; // @[lut_35.scala 2154:102 lut_35.scala 2189:43]
  wire  _GEN_4271 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_4010; // @[lut_35.scala 2154:102 lut_35.scala 2190:43]
  wire  _GEN_4272 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_4011; // @[lut_35.scala 2154:102 lut_35.scala 2191:43]
  wire  _GEN_4273 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] | _GEN_4012; // @[lut_35.scala 2154:102 lut_35.scala 2192:38]
  wire  _GEN_4277 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2154:102 lut_35.scala 177:26 lut_35.scala 2194:87]
  wire  _GEN_4285 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_4016; // @[lut_35.scala 2154:102 lut_35.scala 177:26]
  wire  _GEN_4293 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_4024; // @[lut_35.scala 2154:102 lut_35.scala 177:26]
  wire  _GEN_4301 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_4032; // @[lut_35.scala 2154:102 lut_35.scala 177:26]
  wire  _GEN_4309 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_4040; // @[lut_35.scala 2154:102 lut_35.scala 177:26]
  wire  _GEN_4317 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_4048; // @[lut_35.scala 2154:102 lut_35.scala 177:26]
  wire  _GEN_4325 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_4056; // @[lut_35.scala 2154:102 lut_35.scala 177:26]
  wire  _GEN_4333 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_4064; // @[lut_35.scala 2154:102 lut_35.scala 177:26]
  wire  _GEN_4341 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_4072; // @[lut_35.scala 2154:102 lut_35.scala 177:26]
  wire  _GEN_4349 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_4080; // @[lut_35.scala 2154:102 lut_35.scala 177:26]
  wire  _GEN_4357 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_4088; // @[lut_35.scala 2154:102 lut_35.scala 177:26]
  wire  _GEN_4365 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_4096; // @[lut_35.scala 2154:102 lut_35.scala 177:26]
  wire  _GEN_4373 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_4104; // @[lut_35.scala 2154:102 lut_35.scala 177:26]
  wire  _GEN_4381 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_4112; // @[lut_35.scala 2154:102 lut_35.scala 177:26]
  wire  _GEN_4389 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_4120; // @[lut_35.scala 2154:102 lut_35.scala 177:26]
  wire  _GEN_4397 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_4128; // @[lut_35.scala 2154:102 lut_35.scala 177:26]
  wire  _GEN_4405 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_4136; // @[lut_35.scala 2154:102 lut_35.scala 177:26]
  wire  _GEN_4413 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_4144; // @[lut_35.scala 2154:102 lut_35.scala 177:26]
  wire  _GEN_4421 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_4152; // @[lut_35.scala 2154:102 lut_35.scala 177:26]
  wire  _GEN_4429 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_4160; // @[lut_35.scala 2154:102 lut_35.scala 177:26]
  wire  _GEN_4437 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_4168; // @[lut_35.scala 2154:102 lut_35.scala 177:26]
  wire  _GEN_4445 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_4176; // @[lut_35.scala 2154:102 lut_35.scala 177:26]
  wire  _GEN_4453 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_4184; // @[lut_35.scala 2154:102 lut_35.scala 177:26]
  wire  _GEN_4461 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_4192; // @[lut_35.scala 2154:102 lut_35.scala 177:26]
  wire  _GEN_4469 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_4200; // @[lut_35.scala 2154:102 lut_35.scala 177:26]
  wire  _GEN_4477 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_4208; // @[lut_35.scala 2154:102 lut_35.scala 177:26]
  wire  _GEN_4485 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_4216; // @[lut_35.scala 2154:102 lut_35.scala 177:26]
  wire  _GEN_4493 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_4224; // @[lut_35.scala 2154:102 lut_35.scala 177:26]
  wire  _GEN_4501 = io_empty_5 & push_valid & ~push_5_1 & ~LUT_mem_MPORT_220_data[32] ? 1'h0 : _GEN_4232; // @[lut_35.scala 2154:102 lut_35.scala 177:26]
  wire  _GEN_4513 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _T_373; // @[lut_35.scala 2114:102 lut_35.scala 2122:42]
  wire  _GEN_4514 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4244; // @[lut_35.scala 2114:102 lut_35.scala 2123:42]
  wire  _GEN_4515 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4245; // @[lut_35.scala 2114:102 lut_35.scala 2124:42]
  wire  _GEN_4516 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4246; // @[lut_35.scala 2114:102 lut_35.scala 2125:42]
  wire  _GEN_4517 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4247; // @[lut_35.scala 2114:102 lut_35.scala 2126:42]
  wire  _GEN_4518 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4248; // @[lut_35.scala 2114:102 lut_35.scala 2127:43]
  wire  _GEN_4519 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4249; // @[lut_35.scala 2114:102 lut_35.scala 2128:43]
  wire  _GEN_4520 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4250; // @[lut_35.scala 2114:102 lut_35.scala 2129:43]
  wire  _GEN_4521 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4251; // @[lut_35.scala 2114:102 lut_35.scala 2130:43]
  wire  _GEN_4522 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4252; // @[lut_35.scala 2114:102 lut_35.scala 2131:43]
  wire  _GEN_4523 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4253; // @[lut_35.scala 2114:102 lut_35.scala 2132:43]
  wire  _GEN_4524 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4254; // @[lut_35.scala 2114:102 lut_35.scala 2133:43]
  wire  _GEN_4525 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4255; // @[lut_35.scala 2114:102 lut_35.scala 2134:43]
  wire  _GEN_4526 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4256; // @[lut_35.scala 2114:102 lut_35.scala 2135:43]
  wire  _GEN_4527 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4257; // @[lut_35.scala 2114:102 lut_35.scala 2136:43]
  wire  _GEN_4528 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4258; // @[lut_35.scala 2114:102 lut_35.scala 2137:43]
  wire  _GEN_4529 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4259; // @[lut_35.scala 2114:102 lut_35.scala 2138:43]
  wire  _GEN_4530 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4260; // @[lut_35.scala 2114:102 lut_35.scala 2139:43]
  wire  _GEN_4531 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4261; // @[lut_35.scala 2114:102 lut_35.scala 2140:43]
  wire  _GEN_4532 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4262; // @[lut_35.scala 2114:102 lut_35.scala 2141:43]
  wire  _GEN_4533 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4263; // @[lut_35.scala 2114:102 lut_35.scala 2142:43]
  wire  _GEN_4534 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4264; // @[lut_35.scala 2114:102 lut_35.scala 2143:43]
  wire  _GEN_4535 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4265; // @[lut_35.scala 2114:102 lut_35.scala 2144:43]
  wire  _GEN_4536 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4266; // @[lut_35.scala 2114:102 lut_35.scala 2145:43]
  wire  _GEN_4537 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4267; // @[lut_35.scala 2114:102 lut_35.scala 2146:43]
  wire  _GEN_4538 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4268; // @[lut_35.scala 2114:102 lut_35.scala 2147:43]
  wire  _GEN_4539 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4269; // @[lut_35.scala 2114:102 lut_35.scala 2148:43]
  wire  _GEN_4540 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4270; // @[lut_35.scala 2114:102 lut_35.scala 2149:43]
  wire  _GEN_4541 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4271; // @[lut_35.scala 2114:102 lut_35.scala 2150:43]
  wire  _GEN_4542 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4272; // @[lut_35.scala 2114:102 lut_35.scala 2151:43]
  wire  _GEN_4543 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] | _GEN_4273; // @[lut_35.scala 2114:102 lut_35.scala 2152:38]
  wire  _GEN_4547 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2114:102 lut_35.scala 177:26 lut_35.scala 2154:87]
  wire  _GEN_4555 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4277; // @[lut_35.scala 2114:102 lut_35.scala 177:26]
  wire  _GEN_4563 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4285; // @[lut_35.scala 2114:102 lut_35.scala 177:26]
  wire  _GEN_4571 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4293; // @[lut_35.scala 2114:102 lut_35.scala 177:26]
  wire  _GEN_4579 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4301; // @[lut_35.scala 2114:102 lut_35.scala 177:26]
  wire  _GEN_4587 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4309; // @[lut_35.scala 2114:102 lut_35.scala 177:26]
  wire  _GEN_4595 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4317; // @[lut_35.scala 2114:102 lut_35.scala 177:26]
  wire  _GEN_4603 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4325; // @[lut_35.scala 2114:102 lut_35.scala 177:26]
  wire  _GEN_4611 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4333; // @[lut_35.scala 2114:102 lut_35.scala 177:26]
  wire  _GEN_4619 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4341; // @[lut_35.scala 2114:102 lut_35.scala 177:26]
  wire  _GEN_4627 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4349; // @[lut_35.scala 2114:102 lut_35.scala 177:26]
  wire  _GEN_4635 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4357; // @[lut_35.scala 2114:102 lut_35.scala 177:26]
  wire  _GEN_4643 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4365; // @[lut_35.scala 2114:102 lut_35.scala 177:26]
  wire  _GEN_4651 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4373; // @[lut_35.scala 2114:102 lut_35.scala 177:26]
  wire  _GEN_4659 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4381; // @[lut_35.scala 2114:102 lut_35.scala 177:26]
  wire  _GEN_4667 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4389; // @[lut_35.scala 2114:102 lut_35.scala 177:26]
  wire  _GEN_4675 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4397; // @[lut_35.scala 2114:102 lut_35.scala 177:26]
  wire  _GEN_4683 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4405; // @[lut_35.scala 2114:102 lut_35.scala 177:26]
  wire  _GEN_4691 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4413; // @[lut_35.scala 2114:102 lut_35.scala 177:26]
  wire  _GEN_4699 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4421; // @[lut_35.scala 2114:102 lut_35.scala 177:26]
  wire  _GEN_4707 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4429; // @[lut_35.scala 2114:102 lut_35.scala 177:26]
  wire  _GEN_4715 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4437; // @[lut_35.scala 2114:102 lut_35.scala 177:26]
  wire  _GEN_4723 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4445; // @[lut_35.scala 2114:102 lut_35.scala 177:26]
  wire  _GEN_4731 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4453; // @[lut_35.scala 2114:102 lut_35.scala 177:26]
  wire  _GEN_4739 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4461; // @[lut_35.scala 2114:102 lut_35.scala 177:26]
  wire  _GEN_4747 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4469; // @[lut_35.scala 2114:102 lut_35.scala 177:26]
  wire  _GEN_4755 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4477; // @[lut_35.scala 2114:102 lut_35.scala 177:26]
  wire  _GEN_4763 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4485; // @[lut_35.scala 2114:102 lut_35.scala 177:26]
  wire  _GEN_4771 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4493; // @[lut_35.scala 2114:102 lut_35.scala 177:26]
  wire  _GEN_4779 = io_empty_4 & push_valid & ~push_4_1 & ~LUT_mem_MPORT_218_data[32] ? 1'h0 : _GEN_4501; // @[lut_35.scala 2114:102 lut_35.scala 177:26]
  wire  _GEN_4791 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _T_364; // @[lut_35.scala 2074:102 lut_35.scala 2081:42]
  wire  _GEN_4792 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4513; // @[lut_35.scala 2074:102 lut_35.scala 2082:42]
  wire  _GEN_4793 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4514; // @[lut_35.scala 2074:102 lut_35.scala 2083:42]
  wire  _GEN_4794 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4515; // @[lut_35.scala 2074:102 lut_35.scala 2084:42]
  wire  _GEN_4795 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4516; // @[lut_35.scala 2074:102 lut_35.scala 2085:42]
  wire  _GEN_4796 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4517; // @[lut_35.scala 2074:102 lut_35.scala 2086:42]
  wire  _GEN_4797 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4518; // @[lut_35.scala 2074:102 lut_35.scala 2087:43]
  wire  _GEN_4798 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4519; // @[lut_35.scala 2074:102 lut_35.scala 2088:43]
  wire  _GEN_4799 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4520; // @[lut_35.scala 2074:102 lut_35.scala 2089:43]
  wire  _GEN_4800 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4521; // @[lut_35.scala 2074:102 lut_35.scala 2090:43]
  wire  _GEN_4801 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4522; // @[lut_35.scala 2074:102 lut_35.scala 2091:43]
  wire  _GEN_4802 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4523; // @[lut_35.scala 2074:102 lut_35.scala 2092:43]
  wire  _GEN_4803 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4524; // @[lut_35.scala 2074:102 lut_35.scala 2093:43]
  wire  _GEN_4804 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4525; // @[lut_35.scala 2074:102 lut_35.scala 2094:43]
  wire  _GEN_4805 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4526; // @[lut_35.scala 2074:102 lut_35.scala 2095:43]
  wire  _GEN_4806 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4527; // @[lut_35.scala 2074:102 lut_35.scala 2096:43]
  wire  _GEN_4807 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4528; // @[lut_35.scala 2074:102 lut_35.scala 2097:43]
  wire  _GEN_4808 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4529; // @[lut_35.scala 2074:102 lut_35.scala 2098:43]
  wire  _GEN_4809 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4530; // @[lut_35.scala 2074:102 lut_35.scala 2099:43]
  wire  _GEN_4810 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4531; // @[lut_35.scala 2074:102 lut_35.scala 2100:43]
  wire  _GEN_4811 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4532; // @[lut_35.scala 2074:102 lut_35.scala 2101:43]
  wire  _GEN_4812 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4533; // @[lut_35.scala 2074:102 lut_35.scala 2102:43]
  wire  _GEN_4813 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4534; // @[lut_35.scala 2074:102 lut_35.scala 2103:43]
  wire  _GEN_4814 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4535; // @[lut_35.scala 2074:102 lut_35.scala 2104:43]
  wire  _GEN_4815 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4536; // @[lut_35.scala 2074:102 lut_35.scala 2105:43]
  wire  _GEN_4816 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4537; // @[lut_35.scala 2074:102 lut_35.scala 2106:43]
  wire  _GEN_4817 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4538; // @[lut_35.scala 2074:102 lut_35.scala 2107:43]
  wire  _GEN_4818 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4539; // @[lut_35.scala 2074:102 lut_35.scala 2108:43]
  wire  _GEN_4819 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4540; // @[lut_35.scala 2074:102 lut_35.scala 2109:43]
  wire  _GEN_4820 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4541; // @[lut_35.scala 2074:102 lut_35.scala 2110:43]
  wire  _GEN_4821 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4542; // @[lut_35.scala 2074:102 lut_35.scala 2111:43]
  wire  _GEN_4822 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] | _GEN_4543; // @[lut_35.scala 2074:102 lut_35.scala 2112:38]
  wire  _GEN_4826 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2074:102 lut_35.scala 177:26 lut_35.scala 2114:87]
  wire  _GEN_4834 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4547; // @[lut_35.scala 2074:102 lut_35.scala 177:26]
  wire  _GEN_4842 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4555; // @[lut_35.scala 2074:102 lut_35.scala 177:26]
  wire  _GEN_4850 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4563; // @[lut_35.scala 2074:102 lut_35.scala 177:26]
  wire  _GEN_4858 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4571; // @[lut_35.scala 2074:102 lut_35.scala 177:26]
  wire  _GEN_4866 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4579; // @[lut_35.scala 2074:102 lut_35.scala 177:26]
  wire  _GEN_4874 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4587; // @[lut_35.scala 2074:102 lut_35.scala 177:26]
  wire  _GEN_4882 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4595; // @[lut_35.scala 2074:102 lut_35.scala 177:26]
  wire  _GEN_4890 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4603; // @[lut_35.scala 2074:102 lut_35.scala 177:26]
  wire  _GEN_4898 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4611; // @[lut_35.scala 2074:102 lut_35.scala 177:26]
  wire  _GEN_4906 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4619; // @[lut_35.scala 2074:102 lut_35.scala 177:26]
  wire  _GEN_4914 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4627; // @[lut_35.scala 2074:102 lut_35.scala 177:26]
  wire  _GEN_4922 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4635; // @[lut_35.scala 2074:102 lut_35.scala 177:26]
  wire  _GEN_4930 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4643; // @[lut_35.scala 2074:102 lut_35.scala 177:26]
  wire  _GEN_4938 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4651; // @[lut_35.scala 2074:102 lut_35.scala 177:26]
  wire  _GEN_4946 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4659; // @[lut_35.scala 2074:102 lut_35.scala 177:26]
  wire  _GEN_4954 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4667; // @[lut_35.scala 2074:102 lut_35.scala 177:26]
  wire  _GEN_4962 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4675; // @[lut_35.scala 2074:102 lut_35.scala 177:26]
  wire  _GEN_4970 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4683; // @[lut_35.scala 2074:102 lut_35.scala 177:26]
  wire  _GEN_4978 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4691; // @[lut_35.scala 2074:102 lut_35.scala 177:26]
  wire  _GEN_4986 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4699; // @[lut_35.scala 2074:102 lut_35.scala 177:26]
  wire  _GEN_4994 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4707; // @[lut_35.scala 2074:102 lut_35.scala 177:26]
  wire  _GEN_5002 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4715; // @[lut_35.scala 2074:102 lut_35.scala 177:26]
  wire  _GEN_5010 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4723; // @[lut_35.scala 2074:102 lut_35.scala 177:26]
  wire  _GEN_5018 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4731; // @[lut_35.scala 2074:102 lut_35.scala 177:26]
  wire  _GEN_5026 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4739; // @[lut_35.scala 2074:102 lut_35.scala 177:26]
  wire  _GEN_5034 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4747; // @[lut_35.scala 2074:102 lut_35.scala 177:26]
  wire  _GEN_5042 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4755; // @[lut_35.scala 2074:102 lut_35.scala 177:26]
  wire  _GEN_5050 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4763; // @[lut_35.scala 2074:102 lut_35.scala 177:26]
  wire  _GEN_5058 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4771; // @[lut_35.scala 2074:102 lut_35.scala 177:26]
  wire  _GEN_5066 = io_empty_3 & push_valid & ~push_3_1 & ~LUT_mem_MPORT_216_data[32] ? 1'h0 : _GEN_4779; // @[lut_35.scala 2074:102 lut_35.scala 177:26]
  wire  _GEN_5078 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _T_355; // @[lut_35.scala 2034:102 lut_35.scala 2040:42]
  wire  _GEN_5079 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4791; // @[lut_35.scala 2034:102 lut_35.scala 2041:42]
  wire  _GEN_5080 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4792; // @[lut_35.scala 2034:102 lut_35.scala 2042:42]
  wire  _GEN_5081 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4793; // @[lut_35.scala 2034:102 lut_35.scala 2043:42]
  wire  _GEN_5082 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4794; // @[lut_35.scala 2034:102 lut_35.scala 2044:42]
  wire  _GEN_5083 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4795; // @[lut_35.scala 2034:102 lut_35.scala 2045:42]
  wire  _GEN_5084 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4796; // @[lut_35.scala 2034:102 lut_35.scala 2046:42]
  wire  _GEN_5085 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4797; // @[lut_35.scala 2034:102 lut_35.scala 2047:43]
  wire  _GEN_5086 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4798; // @[lut_35.scala 2034:102 lut_35.scala 2048:43]
  wire  _GEN_5087 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4799; // @[lut_35.scala 2034:102 lut_35.scala 2049:43]
  wire  _GEN_5088 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4800; // @[lut_35.scala 2034:102 lut_35.scala 2050:43]
  wire  _GEN_5089 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4801; // @[lut_35.scala 2034:102 lut_35.scala 2051:43]
  wire  _GEN_5090 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4802; // @[lut_35.scala 2034:102 lut_35.scala 2052:43]
  wire  _GEN_5091 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4803; // @[lut_35.scala 2034:102 lut_35.scala 2053:43]
  wire  _GEN_5092 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4804; // @[lut_35.scala 2034:102 lut_35.scala 2054:43]
  wire  _GEN_5093 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4805; // @[lut_35.scala 2034:102 lut_35.scala 2055:43]
  wire  _GEN_5094 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4806; // @[lut_35.scala 2034:102 lut_35.scala 2056:43]
  wire  _GEN_5095 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4807; // @[lut_35.scala 2034:102 lut_35.scala 2057:43]
  wire  _GEN_5096 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4808; // @[lut_35.scala 2034:102 lut_35.scala 2058:43]
  wire  _GEN_5097 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4809; // @[lut_35.scala 2034:102 lut_35.scala 2059:43]
  wire  _GEN_5098 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4810; // @[lut_35.scala 2034:102 lut_35.scala 2060:43]
  wire  _GEN_5099 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4811; // @[lut_35.scala 2034:102 lut_35.scala 2061:43]
  wire  _GEN_5100 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4812; // @[lut_35.scala 2034:102 lut_35.scala 2062:43]
  wire  _GEN_5101 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4813; // @[lut_35.scala 2034:102 lut_35.scala 2063:43]
  wire  _GEN_5102 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4814; // @[lut_35.scala 2034:102 lut_35.scala 2064:43]
  wire  _GEN_5103 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4815; // @[lut_35.scala 2034:102 lut_35.scala 2065:43]
  wire  _GEN_5104 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4816; // @[lut_35.scala 2034:102 lut_35.scala 2066:43]
  wire  _GEN_5105 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4817; // @[lut_35.scala 2034:102 lut_35.scala 2067:43]
  wire  _GEN_5106 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4818; // @[lut_35.scala 2034:102 lut_35.scala 2068:43]
  wire  _GEN_5107 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4819; // @[lut_35.scala 2034:102 lut_35.scala 2069:43]
  wire  _GEN_5108 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4820; // @[lut_35.scala 2034:102 lut_35.scala 2070:43]
  wire  _GEN_5109 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4821; // @[lut_35.scala 2034:102 lut_35.scala 2071:43]
  wire  _GEN_5110 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] | _GEN_4822; // @[lut_35.scala 2034:102 lut_35.scala 2072:38]
  wire  _GEN_5114 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 2034:102 lut_35.scala 177:26 lut_35.scala 2074:87]
  wire  _GEN_5122 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4826; // @[lut_35.scala 2034:102 lut_35.scala 177:26]
  wire  _GEN_5130 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4834; // @[lut_35.scala 2034:102 lut_35.scala 177:26]
  wire  _GEN_5138 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4842; // @[lut_35.scala 2034:102 lut_35.scala 177:26]
  wire  _GEN_5146 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4850; // @[lut_35.scala 2034:102 lut_35.scala 177:26]
  wire  _GEN_5154 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4858; // @[lut_35.scala 2034:102 lut_35.scala 177:26]
  wire  _GEN_5162 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4866; // @[lut_35.scala 2034:102 lut_35.scala 177:26]
  wire  _GEN_5170 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4874; // @[lut_35.scala 2034:102 lut_35.scala 177:26]
  wire  _GEN_5178 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4882; // @[lut_35.scala 2034:102 lut_35.scala 177:26]
  wire  _GEN_5186 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4890; // @[lut_35.scala 2034:102 lut_35.scala 177:26]
  wire  _GEN_5194 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4898; // @[lut_35.scala 2034:102 lut_35.scala 177:26]
  wire  _GEN_5202 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4906; // @[lut_35.scala 2034:102 lut_35.scala 177:26]
  wire  _GEN_5210 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4914; // @[lut_35.scala 2034:102 lut_35.scala 177:26]
  wire  _GEN_5218 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4922; // @[lut_35.scala 2034:102 lut_35.scala 177:26]
  wire  _GEN_5226 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4930; // @[lut_35.scala 2034:102 lut_35.scala 177:26]
  wire  _GEN_5234 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4938; // @[lut_35.scala 2034:102 lut_35.scala 177:26]
  wire  _GEN_5242 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4946; // @[lut_35.scala 2034:102 lut_35.scala 177:26]
  wire  _GEN_5250 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4954; // @[lut_35.scala 2034:102 lut_35.scala 177:26]
  wire  _GEN_5258 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4962; // @[lut_35.scala 2034:102 lut_35.scala 177:26]
  wire  _GEN_5266 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4970; // @[lut_35.scala 2034:102 lut_35.scala 177:26]
  wire  _GEN_5274 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4978; // @[lut_35.scala 2034:102 lut_35.scala 177:26]
  wire  _GEN_5282 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4986; // @[lut_35.scala 2034:102 lut_35.scala 177:26]
  wire  _GEN_5290 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_4994; // @[lut_35.scala 2034:102 lut_35.scala 177:26]
  wire  _GEN_5298 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_5002; // @[lut_35.scala 2034:102 lut_35.scala 177:26]
  wire  _GEN_5306 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_5010; // @[lut_35.scala 2034:102 lut_35.scala 177:26]
  wire  _GEN_5314 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_5018; // @[lut_35.scala 2034:102 lut_35.scala 177:26]
  wire  _GEN_5322 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_5026; // @[lut_35.scala 2034:102 lut_35.scala 177:26]
  wire  _GEN_5330 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_5034; // @[lut_35.scala 2034:102 lut_35.scala 177:26]
  wire  _GEN_5338 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_5042; // @[lut_35.scala 2034:102 lut_35.scala 177:26]
  wire  _GEN_5346 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_5050; // @[lut_35.scala 2034:102 lut_35.scala 177:26]
  wire  _GEN_5354 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_5058; // @[lut_35.scala 2034:102 lut_35.scala 177:26]
  wire  _GEN_5362 = io_empty_2 & push_valid & ~push_2_1 & ~LUT_mem_MPORT_214_data[32] ? 1'h0 : _GEN_5066; // @[lut_35.scala 2034:102 lut_35.scala 177:26]
  wire  _GEN_5373 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _T_346; // @[lut_35.scala 1994:102 lut_35.scala 1999:42]
  wire  _GEN_5374 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5078; // @[lut_35.scala 1994:102 lut_35.scala 2000:42]
  wire  _GEN_5375 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5079; // @[lut_35.scala 1994:102 lut_35.scala 2001:42]
  wire  _GEN_5376 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5080; // @[lut_35.scala 1994:102 lut_35.scala 2002:42]
  wire  _GEN_5377 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5081; // @[lut_35.scala 1994:102 lut_35.scala 2003:42]
  wire  _GEN_5378 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5082; // @[lut_35.scala 1994:102 lut_35.scala 2004:42]
  wire  _GEN_5379 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5083; // @[lut_35.scala 1994:102 lut_35.scala 2005:42]
  wire  _GEN_5380 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5084; // @[lut_35.scala 1994:102 lut_35.scala 2006:42]
  wire  _GEN_5381 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5085; // @[lut_35.scala 1994:102 lut_35.scala 2007:43]
  wire  _GEN_5382 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5086; // @[lut_35.scala 1994:102 lut_35.scala 2008:43]
  wire  _GEN_5383 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5087; // @[lut_35.scala 1994:102 lut_35.scala 2009:43]
  wire  _GEN_5384 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5088; // @[lut_35.scala 1994:102 lut_35.scala 2010:43]
  wire  _GEN_5385 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5089; // @[lut_35.scala 1994:102 lut_35.scala 2011:43]
  wire  _GEN_5386 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5090; // @[lut_35.scala 1994:102 lut_35.scala 2012:43]
  wire  _GEN_5387 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5091; // @[lut_35.scala 1994:102 lut_35.scala 2013:43]
  wire  _GEN_5388 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5092; // @[lut_35.scala 1994:102 lut_35.scala 2014:43]
  wire  _GEN_5389 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5093; // @[lut_35.scala 1994:102 lut_35.scala 2015:43]
  wire  _GEN_5390 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5094; // @[lut_35.scala 1994:102 lut_35.scala 2016:43]
  wire  _GEN_5391 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5095; // @[lut_35.scala 1994:102 lut_35.scala 2017:43]
  wire  _GEN_5392 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5096; // @[lut_35.scala 1994:102 lut_35.scala 2018:43]
  wire  _GEN_5393 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5097; // @[lut_35.scala 1994:102 lut_35.scala 2019:43]
  wire  _GEN_5394 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5098; // @[lut_35.scala 1994:102 lut_35.scala 2020:43]
  wire  _GEN_5395 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5099; // @[lut_35.scala 1994:102 lut_35.scala 2021:43]
  wire  _GEN_5396 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5100; // @[lut_35.scala 1994:102 lut_35.scala 2022:43]
  wire  _GEN_5397 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5101; // @[lut_35.scala 1994:102 lut_35.scala 2023:43]
  wire  _GEN_5398 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5102; // @[lut_35.scala 1994:102 lut_35.scala 2024:43]
  wire  _GEN_5399 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5103; // @[lut_35.scala 1994:102 lut_35.scala 2025:43]
  wire  _GEN_5400 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5104; // @[lut_35.scala 1994:102 lut_35.scala 2026:43]
  wire  _GEN_5401 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5105; // @[lut_35.scala 1994:102 lut_35.scala 2027:43]
  wire  _GEN_5402 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5106; // @[lut_35.scala 1994:102 lut_35.scala 2028:43]
  wire  _GEN_5403 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5107; // @[lut_35.scala 1994:102 lut_35.scala 2029:43]
  wire  _GEN_5404 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5108; // @[lut_35.scala 1994:102 lut_35.scala 2030:43]
  wire  _GEN_5405 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5109; // @[lut_35.scala 1994:102 lut_35.scala 2031:43]
  wire  _GEN_5406 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] | _GEN_5110; // @[lut_35.scala 1994:102 lut_35.scala 2032:38]
  wire  _GEN_5410 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 1994:102 lut_35.scala 177:26 lut_35.scala 2034:87]
  wire  _GEN_5418 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5114; // @[lut_35.scala 1994:102 lut_35.scala 177:26]
  wire  _GEN_5426 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5122; // @[lut_35.scala 1994:102 lut_35.scala 177:26]
  wire  _GEN_5434 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5130; // @[lut_35.scala 1994:102 lut_35.scala 177:26]
  wire  _GEN_5442 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5138; // @[lut_35.scala 1994:102 lut_35.scala 177:26]
  wire  _GEN_5450 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5146; // @[lut_35.scala 1994:102 lut_35.scala 177:26]
  wire  _GEN_5458 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5154; // @[lut_35.scala 1994:102 lut_35.scala 177:26]
  wire  _GEN_5466 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5162; // @[lut_35.scala 1994:102 lut_35.scala 177:26]
  wire  _GEN_5474 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5170; // @[lut_35.scala 1994:102 lut_35.scala 177:26]
  wire  _GEN_5482 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5178; // @[lut_35.scala 1994:102 lut_35.scala 177:26]
  wire  _GEN_5490 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5186; // @[lut_35.scala 1994:102 lut_35.scala 177:26]
  wire  _GEN_5498 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5194; // @[lut_35.scala 1994:102 lut_35.scala 177:26]
  wire  _GEN_5506 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5202; // @[lut_35.scala 1994:102 lut_35.scala 177:26]
  wire  _GEN_5514 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5210; // @[lut_35.scala 1994:102 lut_35.scala 177:26]
  wire  _GEN_5522 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5218; // @[lut_35.scala 1994:102 lut_35.scala 177:26]
  wire  _GEN_5530 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5226; // @[lut_35.scala 1994:102 lut_35.scala 177:26]
  wire  _GEN_5538 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5234; // @[lut_35.scala 1994:102 lut_35.scala 177:26]
  wire  _GEN_5546 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5242; // @[lut_35.scala 1994:102 lut_35.scala 177:26]
  wire  _GEN_5554 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5250; // @[lut_35.scala 1994:102 lut_35.scala 177:26]
  wire  _GEN_5562 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5258; // @[lut_35.scala 1994:102 lut_35.scala 177:26]
  wire  _GEN_5570 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5266; // @[lut_35.scala 1994:102 lut_35.scala 177:26]
  wire  _GEN_5578 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5274; // @[lut_35.scala 1994:102 lut_35.scala 177:26]
  wire  _GEN_5586 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5282; // @[lut_35.scala 1994:102 lut_35.scala 177:26]
  wire  _GEN_5594 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5290; // @[lut_35.scala 1994:102 lut_35.scala 177:26]
  wire  _GEN_5602 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5298; // @[lut_35.scala 1994:102 lut_35.scala 177:26]
  wire  _GEN_5610 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5306; // @[lut_35.scala 1994:102 lut_35.scala 177:26]
  wire  _GEN_5618 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5314; // @[lut_35.scala 1994:102 lut_35.scala 177:26]
  wire  _GEN_5626 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5322; // @[lut_35.scala 1994:102 lut_35.scala 177:26]
  wire  _GEN_5634 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5330; // @[lut_35.scala 1994:102 lut_35.scala 177:26]
  wire  _GEN_5642 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5338; // @[lut_35.scala 1994:102 lut_35.scala 177:26]
  wire  _GEN_5650 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5346; // @[lut_35.scala 1994:102 lut_35.scala 177:26]
  wire  _GEN_5658 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5354; // @[lut_35.scala 1994:102 lut_35.scala 177:26]
  wire  _GEN_5666 = io_empty_1 & push_valid & ~push_1_1 & ~LUT_mem_MPORT_212_data[32] ? 1'h0 : _GEN_5362; // @[lut_35.scala 1994:102 lut_35.scala 177:26]
  wire  _GEN_5677 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _T_337; // @[lut_35.scala 1954:103 lut_35.scala 1958:42]
  wire  _GEN_5678 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5373; // @[lut_35.scala 1954:103 lut_35.scala 1959:42]
  wire  _GEN_5679 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5374; // @[lut_35.scala 1954:103 lut_35.scala 1960:42]
  wire  _GEN_5680 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5375; // @[lut_35.scala 1954:103 lut_35.scala 1961:42]
  wire  _GEN_5681 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5376; // @[lut_35.scala 1954:103 lut_35.scala 1962:42]
  wire  _GEN_5682 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5377; // @[lut_35.scala 1954:103 lut_35.scala 1963:42]
  wire  _GEN_5683 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5378; // @[lut_35.scala 1954:103 lut_35.scala 1964:42]
  wire  _GEN_5684 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5379; // @[lut_35.scala 1954:103 lut_35.scala 1965:42]
  wire  _GEN_5685 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5380; // @[lut_35.scala 1954:103 lut_35.scala 1966:42]
  wire  _GEN_5686 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5381; // @[lut_35.scala 1954:103 lut_35.scala 1967:43]
  wire  _GEN_5687 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5382; // @[lut_35.scala 1954:103 lut_35.scala 1968:43]
  wire  _GEN_5688 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5383; // @[lut_35.scala 1954:103 lut_35.scala 1969:43]
  wire  _GEN_5689 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5384; // @[lut_35.scala 1954:103 lut_35.scala 1970:43]
  wire  _GEN_5690 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5385; // @[lut_35.scala 1954:103 lut_35.scala 1971:43]
  wire  _GEN_5691 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5386; // @[lut_35.scala 1954:103 lut_35.scala 1972:43]
  wire  _GEN_5692 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5387; // @[lut_35.scala 1954:103 lut_35.scala 1973:43]
  wire  _GEN_5693 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5388; // @[lut_35.scala 1954:103 lut_35.scala 1974:43]
  wire  _GEN_5694 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5389; // @[lut_35.scala 1954:103 lut_35.scala 1975:43]
  wire  _GEN_5695 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5390; // @[lut_35.scala 1954:103 lut_35.scala 1976:43]
  wire  _GEN_5696 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5391; // @[lut_35.scala 1954:103 lut_35.scala 1977:43]
  wire  _GEN_5697 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5392; // @[lut_35.scala 1954:103 lut_35.scala 1978:43]
  wire  _GEN_5698 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5393; // @[lut_35.scala 1954:103 lut_35.scala 1979:43]
  wire  _GEN_5699 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5394; // @[lut_35.scala 1954:103 lut_35.scala 1980:43]
  wire  _GEN_5700 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5395; // @[lut_35.scala 1954:103 lut_35.scala 1981:43]
  wire  _GEN_5701 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5396; // @[lut_35.scala 1954:103 lut_35.scala 1982:43]
  wire  _GEN_5702 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5397; // @[lut_35.scala 1954:103 lut_35.scala 1983:43]
  wire  _GEN_5703 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5398; // @[lut_35.scala 1954:103 lut_35.scala 1984:43]
  wire  _GEN_5704 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5399; // @[lut_35.scala 1954:103 lut_35.scala 1985:43]
  wire  _GEN_5705 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5400; // @[lut_35.scala 1954:103 lut_35.scala 1986:43]
  wire  _GEN_5706 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5401; // @[lut_35.scala 1954:103 lut_35.scala 1987:43]
  wire  _GEN_5707 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5402; // @[lut_35.scala 1954:103 lut_35.scala 1988:43]
  wire  _GEN_5708 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5403; // @[lut_35.scala 1954:103 lut_35.scala 1989:43]
  wire  _GEN_5709 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5404; // @[lut_35.scala 1954:103 lut_35.scala 1990:43]
  wire  _GEN_5710 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5405; // @[lut_35.scala 1954:103 lut_35.scala 1991:43]
  wire  _GEN_5711 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] | _GEN_5406; // @[lut_35.scala 1954:103 lut_35.scala 1992:38]
  wire  _GEN_5715 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : 1'h1; // @[lut_35.scala 1954:103 lut_35.scala 177:26 lut_35.scala 1994:87]
  wire  _GEN_5722 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5410; // @[lut_35.scala 1954:103 lut_35.scala 177:26]
  wire  _GEN_5730 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5418; // @[lut_35.scala 1954:103 lut_35.scala 177:26]
  wire  _GEN_5738 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5426; // @[lut_35.scala 1954:103 lut_35.scala 177:26]
  wire  _GEN_5746 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5434; // @[lut_35.scala 1954:103 lut_35.scala 177:26]
  wire  _GEN_5754 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5442; // @[lut_35.scala 1954:103 lut_35.scala 177:26]
  wire  _GEN_5762 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5450; // @[lut_35.scala 1954:103 lut_35.scala 177:26]
  wire  _GEN_5770 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5458; // @[lut_35.scala 1954:103 lut_35.scala 177:26]
  wire  _GEN_5778 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5466; // @[lut_35.scala 1954:103 lut_35.scala 177:26]
  wire  _GEN_5786 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5474; // @[lut_35.scala 1954:103 lut_35.scala 177:26]
  wire  _GEN_5794 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5482; // @[lut_35.scala 1954:103 lut_35.scala 177:26]
  wire  _GEN_5802 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5490; // @[lut_35.scala 1954:103 lut_35.scala 177:26]
  wire  _GEN_5810 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5498; // @[lut_35.scala 1954:103 lut_35.scala 177:26]
  wire  _GEN_5818 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5506; // @[lut_35.scala 1954:103 lut_35.scala 177:26]
  wire  _GEN_5826 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5514; // @[lut_35.scala 1954:103 lut_35.scala 177:26]
  wire  _GEN_5834 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5522; // @[lut_35.scala 1954:103 lut_35.scala 177:26]
  wire  _GEN_5842 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5530; // @[lut_35.scala 1954:103 lut_35.scala 177:26]
  wire  _GEN_5850 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5538; // @[lut_35.scala 1954:103 lut_35.scala 177:26]
  wire  _GEN_5858 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5546; // @[lut_35.scala 1954:103 lut_35.scala 177:26]
  wire  _GEN_5866 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5554; // @[lut_35.scala 1954:103 lut_35.scala 177:26]
  wire  _GEN_5874 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5562; // @[lut_35.scala 1954:103 lut_35.scala 177:26]
  wire  _GEN_5882 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5570; // @[lut_35.scala 1954:103 lut_35.scala 177:26]
  wire  _GEN_5890 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5578; // @[lut_35.scala 1954:103 lut_35.scala 177:26]
  wire  _GEN_5898 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5586; // @[lut_35.scala 1954:103 lut_35.scala 177:26]
  wire  _GEN_5906 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5594; // @[lut_35.scala 1954:103 lut_35.scala 177:26]
  wire  _GEN_5914 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5602; // @[lut_35.scala 1954:103 lut_35.scala 177:26]
  wire  _GEN_5922 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5610; // @[lut_35.scala 1954:103 lut_35.scala 177:26]
  wire  _GEN_5930 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5618; // @[lut_35.scala 1954:103 lut_35.scala 177:26]
  wire  _GEN_5938 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5626; // @[lut_35.scala 1954:103 lut_35.scala 177:26]
  wire  _GEN_5946 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5634; // @[lut_35.scala 1954:103 lut_35.scala 177:26]
  wire  _GEN_5954 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5642; // @[lut_35.scala 1954:103 lut_35.scala 177:26]
  wire  _GEN_5962 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5650; // @[lut_35.scala 1954:103 lut_35.scala 177:26]
  wire  _GEN_5970 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5658; // @[lut_35.scala 1954:103 lut_35.scala 177:26]
  wire  _GEN_5978 = io_empty_0 & push_valid & ~push_0_1 & ~LUT_mem_MPORT_210_data[32] ? 1'h0 : _GEN_5666; // @[lut_35.scala 1954:103 lut_35.scala 177:26]
  wire  _GEN_5988 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _T_328; // @[lut_35.scala 1953:125 lut_35.scala 177:26]
  wire  _GEN_5992 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5677; // @[lut_35.scala 1953:125 lut_35.scala 3395:32]
  wire  _GEN_5993 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5678; // @[lut_35.scala 1953:125 lut_35.scala 3396:32]
  wire  _GEN_5994 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5679; // @[lut_35.scala 1953:125 lut_35.scala 3397:32]
  wire  _GEN_5995 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5680; // @[lut_35.scala 1953:125 lut_35.scala 3398:32]
  wire  _GEN_5996 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5681; // @[lut_35.scala 1953:125 lut_35.scala 3399:32]
  wire  _GEN_5997 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5682; // @[lut_35.scala 1953:125 lut_35.scala 3400:32]
  wire  _GEN_5998 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5683; // @[lut_35.scala 1953:125 lut_35.scala 3401:32]
  wire  _GEN_5999 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5684; // @[lut_35.scala 1953:125 lut_35.scala 3402:42]
  wire  _GEN_6000 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5685; // @[lut_35.scala 1953:125 lut_35.scala 3403:42]
  wire  _GEN_6001 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5686; // @[lut_35.scala 1953:125 lut_35.scala 3404:43]
  wire  _GEN_6002 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5687; // @[lut_35.scala 1953:125 lut_35.scala 3405:43]
  wire  _GEN_6003 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5688; // @[lut_35.scala 1953:125 lut_35.scala 3406:43]
  wire  _GEN_6004 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5689; // @[lut_35.scala 1953:125 lut_35.scala 3407:43]
  wire  _GEN_6005 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5690; // @[lut_35.scala 1953:125 lut_35.scala 3408:43]
  wire  _GEN_6006 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5691; // @[lut_35.scala 1953:125 lut_35.scala 3409:43]
  wire  _GEN_6007 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5692; // @[lut_35.scala 1953:125 lut_35.scala 3410:43]
  wire  _GEN_6008 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5693; // @[lut_35.scala 1953:125 lut_35.scala 3411:43]
  wire  _GEN_6009 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5694; // @[lut_35.scala 1953:125 lut_35.scala 3412:43]
  wire  _GEN_6010 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5695; // @[lut_35.scala 1953:125 lut_35.scala 3413:43]
  wire  _GEN_6011 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5696; // @[lut_35.scala 1953:125 lut_35.scala 3414:43]
  wire  _GEN_6012 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5697; // @[lut_35.scala 1953:125 lut_35.scala 3415:43]
  wire  _GEN_6013 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5698; // @[lut_35.scala 1953:125 lut_35.scala 3416:43]
  wire  _GEN_6014 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5699; // @[lut_35.scala 1953:125 lut_35.scala 3417:43]
  wire  _GEN_6015 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5700; // @[lut_35.scala 1953:125 lut_35.scala 3418:43]
  wire  _GEN_6016 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5701; // @[lut_35.scala 1953:125 lut_35.scala 3419:43]
  wire  _GEN_6017 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5702; // @[lut_35.scala 1953:125 lut_35.scala 3420:43]
  wire  _GEN_6018 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5703; // @[lut_35.scala 1953:125 lut_35.scala 3421:43]
  wire  _GEN_6019 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5704; // @[lut_35.scala 1953:125 lut_35.scala 3422:43]
  wire  _GEN_6020 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5705; // @[lut_35.scala 1953:125 lut_35.scala 3423:43]
  wire  _GEN_6021 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5706; // @[lut_35.scala 1953:125 lut_35.scala 3424:43]
  wire  _GEN_6022 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5707; // @[lut_35.scala 1953:125 lut_35.scala 3425:43]
  wire  _GEN_6023 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5708; // @[lut_35.scala 1953:125 lut_35.scala 3426:43]
  wire  _GEN_6024 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5709; // @[lut_35.scala 1953:125 lut_35.scala 3427:43]
  wire  _GEN_6025 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5710; // @[lut_35.scala 1953:125 lut_35.scala 3428:43]
  wire  _GEN_6026 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5711; // @[lut_35.scala 1953:125 lut_35.scala 3429:30]
  wire  _GEN_6030 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5715; // @[lut_35.scala 1953:125 lut_35.scala 177:26]
  wire  _GEN_6037 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5722; // @[lut_35.scala 1953:125 lut_35.scala 177:26]
  wire  _GEN_6045 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5730; // @[lut_35.scala 1953:125 lut_35.scala 177:26]
  wire  _GEN_6053 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5738; // @[lut_35.scala 1953:125 lut_35.scala 177:26]
  wire  _GEN_6061 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5746; // @[lut_35.scala 1953:125 lut_35.scala 177:26]
  wire  _GEN_6069 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5754; // @[lut_35.scala 1953:125 lut_35.scala 177:26]
  wire  _GEN_6077 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5762; // @[lut_35.scala 1953:125 lut_35.scala 177:26]
  wire  _GEN_6085 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5770; // @[lut_35.scala 1953:125 lut_35.scala 177:26]
  wire  _GEN_6093 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5778; // @[lut_35.scala 1953:125 lut_35.scala 177:26]
  wire  _GEN_6101 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5786; // @[lut_35.scala 1953:125 lut_35.scala 177:26]
  wire  _GEN_6109 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5794; // @[lut_35.scala 1953:125 lut_35.scala 177:26]
  wire  _GEN_6117 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5802; // @[lut_35.scala 1953:125 lut_35.scala 177:26]
  wire  _GEN_6125 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5810; // @[lut_35.scala 1953:125 lut_35.scala 177:26]
  wire  _GEN_6133 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5818; // @[lut_35.scala 1953:125 lut_35.scala 177:26]
  wire  _GEN_6141 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5826; // @[lut_35.scala 1953:125 lut_35.scala 177:26]
  wire  _GEN_6149 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5834; // @[lut_35.scala 1953:125 lut_35.scala 177:26]
  wire  _GEN_6157 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5842; // @[lut_35.scala 1953:125 lut_35.scala 177:26]
  wire  _GEN_6165 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5850; // @[lut_35.scala 1953:125 lut_35.scala 177:26]
  wire  _GEN_6173 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5858; // @[lut_35.scala 1953:125 lut_35.scala 177:26]
  wire  _GEN_6181 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5866; // @[lut_35.scala 1953:125 lut_35.scala 177:26]
  wire  _GEN_6189 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5874; // @[lut_35.scala 1953:125 lut_35.scala 177:26]
  wire  _GEN_6197 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5882; // @[lut_35.scala 1953:125 lut_35.scala 177:26]
  wire  _GEN_6205 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5890; // @[lut_35.scala 1953:125 lut_35.scala 177:26]
  wire  _GEN_6213 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5898; // @[lut_35.scala 1953:125 lut_35.scala 177:26]
  wire  _GEN_6221 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5906; // @[lut_35.scala 1953:125 lut_35.scala 177:26]
  wire  _GEN_6229 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5914; // @[lut_35.scala 1953:125 lut_35.scala 177:26]
  wire  _GEN_6237 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5922; // @[lut_35.scala 1953:125 lut_35.scala 177:26]
  wire  _GEN_6245 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5930; // @[lut_35.scala 1953:125 lut_35.scala 177:26]
  wire  _GEN_6253 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5938; // @[lut_35.scala 1953:125 lut_35.scala 177:26]
  wire  _GEN_6261 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5946; // @[lut_35.scala 1953:125 lut_35.scala 177:26]
  wire  _GEN_6269 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5954; // @[lut_35.scala 1953:125 lut_35.scala 177:26]
  wire  _GEN_6277 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5962; // @[lut_35.scala 1953:125 lut_35.scala 177:26]
  wire  _GEN_6285 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5970; // @[lut_35.scala 1953:125 lut_35.scala 177:26]
  wire  _GEN_6293 = _T_312 & read_stack32 != push_ray_id & read_stack33 != push_ray_id & read_stack34 != push_ray_id &
    push_valid & _GEN_5978; // @[lut_35.scala 1953:125 lut_35.scala 177:26]
  wire  _GEN_6298 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5988; // @[lut_35.scala 1910:74 lut_35.scala 1911:38]
  wire  _GEN_6299 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5992; // @[lut_35.scala 1910:74 lut_35.scala 1912:38]
  wire  _GEN_6300 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5993; // @[lut_35.scala 1910:74 lut_35.scala 1913:38]
  wire  _GEN_6301 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5994; // @[lut_35.scala 1910:74 lut_35.scala 1914:38]
  wire  _GEN_6302 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5995; // @[lut_35.scala 1910:74 lut_35.scala 1915:38]
  wire  _GEN_6303 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5996; // @[lut_35.scala 1910:74 lut_35.scala 1916:38]
  wire  _GEN_6304 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5997; // @[lut_35.scala 1910:74 lut_35.scala 1917:38]
  wire  _GEN_6305 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5998; // @[lut_35.scala 1910:74 lut_35.scala 1918:38]
  wire  _GEN_6306 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_5999; // @[lut_35.scala 1910:74 lut_35.scala 1919:38]
  wire  _GEN_6307 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6000; // @[lut_35.scala 1910:74 lut_35.scala 1920:38]
  wire  _GEN_6308 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6001; // @[lut_35.scala 1910:74 lut_35.scala 1921:39]
  wire  _GEN_6309 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6002; // @[lut_35.scala 1910:74 lut_35.scala 1922:39]
  wire  _GEN_6310 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6003; // @[lut_35.scala 1910:74 lut_35.scala 1923:39]
  wire  _GEN_6311 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6004; // @[lut_35.scala 1910:74 lut_35.scala 1924:39]
  wire  _GEN_6312 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6005; // @[lut_35.scala 1910:74 lut_35.scala 1925:39]
  wire  _GEN_6313 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6006; // @[lut_35.scala 1910:74 lut_35.scala 1926:39]
  wire  _GEN_6314 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6007; // @[lut_35.scala 1910:74 lut_35.scala 1927:39]
  wire  _GEN_6315 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6008; // @[lut_35.scala 1910:74 lut_35.scala 1928:39]
  wire  _GEN_6316 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6009; // @[lut_35.scala 1910:74 lut_35.scala 1929:39]
  wire  _GEN_6317 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6010; // @[lut_35.scala 1910:74 lut_35.scala 1930:39]
  wire  _GEN_6318 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6011; // @[lut_35.scala 1910:74 lut_35.scala 1931:39]
  wire  _GEN_6319 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6012; // @[lut_35.scala 1910:74 lut_35.scala 1932:39]
  wire  _GEN_6320 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6013; // @[lut_35.scala 1910:74 lut_35.scala 1933:39]
  wire  _GEN_6321 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6014; // @[lut_35.scala 1910:74 lut_35.scala 1934:39]
  wire  _GEN_6322 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6015; // @[lut_35.scala 1910:74 lut_35.scala 1935:39]
  wire  _GEN_6323 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6016; // @[lut_35.scala 1910:74 lut_35.scala 1936:39]
  wire  _GEN_6324 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6017; // @[lut_35.scala 1910:74 lut_35.scala 1937:39]
  wire  _GEN_6325 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6018; // @[lut_35.scala 1910:74 lut_35.scala 1938:39]
  wire  _GEN_6326 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6019; // @[lut_35.scala 1910:74 lut_35.scala 1939:39]
  wire  _GEN_6327 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6020; // @[lut_35.scala 1910:74 lut_35.scala 1940:39]
  wire  _GEN_6328 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6021; // @[lut_35.scala 1910:74 lut_35.scala 1941:39]
  wire  _GEN_6329 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6022; // @[lut_35.scala 1910:74 lut_35.scala 1942:39]
  wire  _GEN_6330 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6023; // @[lut_35.scala 1910:74 lut_35.scala 1943:39]
  wire  _GEN_6331 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6024; // @[lut_35.scala 1910:74 lut_35.scala 1944:39]
  wire  _GEN_6332 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid | _GEN_6025; // @[lut_35.scala 1910:74 lut_35.scala 1945:39]
  wire  _GEN_6333 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid | _GEN_6026; // @[lut_35.scala 1910:74 lut_35.scala 1946:34]
  wire  _GEN_6337 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _T_320; // @[lut_35.scala 1910:74 lut_35.scala 177:26]
  wire  _GEN_6345 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6030; // @[lut_35.scala 1910:74 lut_35.scala 177:26]
  wire  _GEN_6352 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6037; // @[lut_35.scala 1910:74 lut_35.scala 177:26]
  wire  _GEN_6360 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6045; // @[lut_35.scala 1910:74 lut_35.scala 177:26]
  wire  _GEN_6368 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6053; // @[lut_35.scala 1910:74 lut_35.scala 177:26]
  wire  _GEN_6376 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6061; // @[lut_35.scala 1910:74 lut_35.scala 177:26]
  wire  _GEN_6384 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6069; // @[lut_35.scala 1910:74 lut_35.scala 177:26]
  wire  _GEN_6392 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6077; // @[lut_35.scala 1910:74 lut_35.scala 177:26]
  wire  _GEN_6400 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6085; // @[lut_35.scala 1910:74 lut_35.scala 177:26]
  wire  _GEN_6408 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6093; // @[lut_35.scala 1910:74 lut_35.scala 177:26]
  wire  _GEN_6416 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6101; // @[lut_35.scala 1910:74 lut_35.scala 177:26]
  wire  _GEN_6424 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6109; // @[lut_35.scala 1910:74 lut_35.scala 177:26]
  wire  _GEN_6432 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6117; // @[lut_35.scala 1910:74 lut_35.scala 177:26]
  wire  _GEN_6440 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6125; // @[lut_35.scala 1910:74 lut_35.scala 177:26]
  wire  _GEN_6448 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6133; // @[lut_35.scala 1910:74 lut_35.scala 177:26]
  wire  _GEN_6456 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6141; // @[lut_35.scala 1910:74 lut_35.scala 177:26]
  wire  _GEN_6464 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6149; // @[lut_35.scala 1910:74 lut_35.scala 177:26]
  wire  _GEN_6472 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6157; // @[lut_35.scala 1910:74 lut_35.scala 177:26]
  wire  _GEN_6480 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6165; // @[lut_35.scala 1910:74 lut_35.scala 177:26]
  wire  _GEN_6488 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6173; // @[lut_35.scala 1910:74 lut_35.scala 177:26]
  wire  _GEN_6496 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6181; // @[lut_35.scala 1910:74 lut_35.scala 177:26]
  wire  _GEN_6504 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6189; // @[lut_35.scala 1910:74 lut_35.scala 177:26]
  wire  _GEN_6512 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6197; // @[lut_35.scala 1910:74 lut_35.scala 177:26]
  wire  _GEN_6520 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6205; // @[lut_35.scala 1910:74 lut_35.scala 177:26]
  wire  _GEN_6528 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6213; // @[lut_35.scala 1910:74 lut_35.scala 177:26]
  wire  _GEN_6536 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6221; // @[lut_35.scala 1910:74 lut_35.scala 177:26]
  wire  _GEN_6544 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6229; // @[lut_35.scala 1910:74 lut_35.scala 177:26]
  wire  _GEN_6552 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6237; // @[lut_35.scala 1910:74 lut_35.scala 177:26]
  wire  _GEN_6560 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6245; // @[lut_35.scala 1910:74 lut_35.scala 177:26]
  wire  _GEN_6568 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6253; // @[lut_35.scala 1910:74 lut_35.scala 177:26]
  wire  _GEN_6576 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6261; // @[lut_35.scala 1910:74 lut_35.scala 177:26]
  wire  _GEN_6584 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6269; // @[lut_35.scala 1910:74 lut_35.scala 177:26]
  wire  _GEN_6592 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6277; // @[lut_35.scala 1910:74 lut_35.scala 177:26]
  wire  _GEN_6600 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6285; // @[lut_35.scala 1910:74 lut_35.scala 177:26]
  wire  _GEN_6608 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6293; // @[lut_35.scala 1910:74 lut_35.scala 177:26]
  wire  _GEN_6611 = LUT_mem_MPORT_209_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6025; // @[lut_35.scala 1910:74 lut_35.scala 177:26]
  wire  _GEN_6614 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6298; // @[lut_35.scala 1872:74 lut_35.scala 1873:38]
  wire  _GEN_6615 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6299; // @[lut_35.scala 1872:74 lut_35.scala 1874:38]
  wire  _GEN_6616 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6300; // @[lut_35.scala 1872:74 lut_35.scala 1875:38]
  wire  _GEN_6617 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6301; // @[lut_35.scala 1872:74 lut_35.scala 1876:38]
  wire  _GEN_6618 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6302; // @[lut_35.scala 1872:74 lut_35.scala 1877:38]
  wire  _GEN_6619 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6303; // @[lut_35.scala 1872:74 lut_35.scala 1878:38]
  wire  _GEN_6620 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6304; // @[lut_35.scala 1872:74 lut_35.scala 1879:38]
  wire  _GEN_6621 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6305; // @[lut_35.scala 1872:74 lut_35.scala 1880:38]
  wire  _GEN_6622 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6306; // @[lut_35.scala 1872:74 lut_35.scala 1881:38]
  wire  _GEN_6623 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6307; // @[lut_35.scala 1872:74 lut_35.scala 1882:38]
  wire  _GEN_6624 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6308; // @[lut_35.scala 1872:74 lut_35.scala 1883:39]
  wire  _GEN_6625 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6309; // @[lut_35.scala 1872:74 lut_35.scala 1884:39]
  wire  _GEN_6626 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6310; // @[lut_35.scala 1872:74 lut_35.scala 1885:39]
  wire  _GEN_6627 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6311; // @[lut_35.scala 1872:74 lut_35.scala 1886:39]
  wire  _GEN_6628 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6312; // @[lut_35.scala 1872:74 lut_35.scala 1887:39]
  wire  _GEN_6629 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6313; // @[lut_35.scala 1872:74 lut_35.scala 1888:39]
  wire  _GEN_6630 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6314; // @[lut_35.scala 1872:74 lut_35.scala 1889:39]
  wire  _GEN_6631 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6315; // @[lut_35.scala 1872:74 lut_35.scala 1890:39]
  wire  _GEN_6632 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6316; // @[lut_35.scala 1872:74 lut_35.scala 1891:39]
  wire  _GEN_6633 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6317; // @[lut_35.scala 1872:74 lut_35.scala 1892:39]
  wire  _GEN_6634 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6318; // @[lut_35.scala 1872:74 lut_35.scala 1893:39]
  wire  _GEN_6635 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6319; // @[lut_35.scala 1872:74 lut_35.scala 1894:39]
  wire  _GEN_6636 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6320; // @[lut_35.scala 1872:74 lut_35.scala 1895:39]
  wire  _GEN_6637 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6321; // @[lut_35.scala 1872:74 lut_35.scala 1896:39]
  wire  _GEN_6638 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6322; // @[lut_35.scala 1872:74 lut_35.scala 1897:39]
  wire  _GEN_6639 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6323; // @[lut_35.scala 1872:74 lut_35.scala 1898:39]
  wire  _GEN_6640 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6324; // @[lut_35.scala 1872:74 lut_35.scala 1899:39]
  wire  _GEN_6641 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6325; // @[lut_35.scala 1872:74 lut_35.scala 1900:39]
  wire  _GEN_6642 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6326; // @[lut_35.scala 1872:74 lut_35.scala 1901:39]
  wire  _GEN_6643 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6327; // @[lut_35.scala 1872:74 lut_35.scala 1902:39]
  wire  _GEN_6644 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6328; // @[lut_35.scala 1872:74 lut_35.scala 1903:39]
  wire  _GEN_6645 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6329; // @[lut_35.scala 1872:74 lut_35.scala 1904:39]
  wire  _GEN_6646 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6330; // @[lut_35.scala 1872:74 lut_35.scala 1905:39]
  wire  _GEN_6647 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid | _GEN_6331; // @[lut_35.scala 1872:74 lut_35.scala 1906:39]
  wire  _GEN_6648 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6332; // @[lut_35.scala 1872:74 lut_35.scala 1907:39]
  wire  _GEN_6649 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid | _GEN_6333; // @[lut_35.scala 1872:74 lut_35.scala 1908:34]
  wire  _GEN_6653 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1872:74 lut_35.scala 177:26 lut_35.scala 1910:27]
  wire  _GEN_6656 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6337; // @[lut_35.scala 1872:74 lut_35.scala 177:26]
  wire  _GEN_6664 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6345; // @[lut_35.scala 1872:74 lut_35.scala 177:26]
  wire  _GEN_6671 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6352; // @[lut_35.scala 1872:74 lut_35.scala 177:26]
  wire  _GEN_6679 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6360; // @[lut_35.scala 1872:74 lut_35.scala 177:26]
  wire  _GEN_6687 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6368; // @[lut_35.scala 1872:74 lut_35.scala 177:26]
  wire  _GEN_6695 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6376; // @[lut_35.scala 1872:74 lut_35.scala 177:26]
  wire  _GEN_6703 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6384; // @[lut_35.scala 1872:74 lut_35.scala 177:26]
  wire  _GEN_6711 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6392; // @[lut_35.scala 1872:74 lut_35.scala 177:26]
  wire  _GEN_6719 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6400; // @[lut_35.scala 1872:74 lut_35.scala 177:26]
  wire  _GEN_6727 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6408; // @[lut_35.scala 1872:74 lut_35.scala 177:26]
  wire  _GEN_6735 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6416; // @[lut_35.scala 1872:74 lut_35.scala 177:26]
  wire  _GEN_6743 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6424; // @[lut_35.scala 1872:74 lut_35.scala 177:26]
  wire  _GEN_6751 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6432; // @[lut_35.scala 1872:74 lut_35.scala 177:26]
  wire  _GEN_6759 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6440; // @[lut_35.scala 1872:74 lut_35.scala 177:26]
  wire  _GEN_6767 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6448; // @[lut_35.scala 1872:74 lut_35.scala 177:26]
  wire  _GEN_6775 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6456; // @[lut_35.scala 1872:74 lut_35.scala 177:26]
  wire  _GEN_6783 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6464; // @[lut_35.scala 1872:74 lut_35.scala 177:26]
  wire  _GEN_6791 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6472; // @[lut_35.scala 1872:74 lut_35.scala 177:26]
  wire  _GEN_6799 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6480; // @[lut_35.scala 1872:74 lut_35.scala 177:26]
  wire  _GEN_6807 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6488; // @[lut_35.scala 1872:74 lut_35.scala 177:26]
  wire  _GEN_6815 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6496; // @[lut_35.scala 1872:74 lut_35.scala 177:26]
  wire  _GEN_6823 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6504; // @[lut_35.scala 1872:74 lut_35.scala 177:26]
  wire  _GEN_6831 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6512; // @[lut_35.scala 1872:74 lut_35.scala 177:26]
  wire  _GEN_6839 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6520; // @[lut_35.scala 1872:74 lut_35.scala 177:26]
  wire  _GEN_6847 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6528; // @[lut_35.scala 1872:74 lut_35.scala 177:26]
  wire  _GEN_6855 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6536; // @[lut_35.scala 1872:74 lut_35.scala 177:26]
  wire  _GEN_6863 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6544; // @[lut_35.scala 1872:74 lut_35.scala 177:26]
  wire  _GEN_6871 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6552; // @[lut_35.scala 1872:74 lut_35.scala 177:26]
  wire  _GEN_6879 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6560; // @[lut_35.scala 1872:74 lut_35.scala 177:26]
  wire  _GEN_6887 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6568; // @[lut_35.scala 1872:74 lut_35.scala 177:26]
  wire  _GEN_6895 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6576; // @[lut_35.scala 1872:74 lut_35.scala 177:26]
  wire  _GEN_6903 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6584; // @[lut_35.scala 1872:74 lut_35.scala 177:26]
  wire  _GEN_6911 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6592; // @[lut_35.scala 1872:74 lut_35.scala 177:26]
  wire  _GEN_6919 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6600; // @[lut_35.scala 1872:74 lut_35.scala 177:26]
  wire  _GEN_6922 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6331; // @[lut_35.scala 1872:74 lut_35.scala 177:26]
  wire  _GEN_6927 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6608; // @[lut_35.scala 1872:74 lut_35.scala 177:26]
  wire  _GEN_6930 = LUT_mem_MPORT_208_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6611; // @[lut_35.scala 1872:74 lut_35.scala 177:26]
  wire  _GEN_6933 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6614; // @[lut_35.scala 1834:74 lut_35.scala 1835:38]
  wire  _GEN_6934 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6615; // @[lut_35.scala 1834:74 lut_35.scala 1836:38]
  wire  _GEN_6935 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6616; // @[lut_35.scala 1834:74 lut_35.scala 1837:38]
  wire  _GEN_6936 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6617; // @[lut_35.scala 1834:74 lut_35.scala 1838:38]
  wire  _GEN_6937 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6618; // @[lut_35.scala 1834:74 lut_35.scala 1839:38]
  wire  _GEN_6938 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6619; // @[lut_35.scala 1834:74 lut_35.scala 1840:38]
  wire  _GEN_6939 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6620; // @[lut_35.scala 1834:74 lut_35.scala 1841:38]
  wire  _GEN_6940 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6621; // @[lut_35.scala 1834:74 lut_35.scala 1842:38]
  wire  _GEN_6941 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6622; // @[lut_35.scala 1834:74 lut_35.scala 1843:38]
  wire  _GEN_6942 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6623; // @[lut_35.scala 1834:74 lut_35.scala 1844:38]
  wire  _GEN_6943 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6624; // @[lut_35.scala 1834:74 lut_35.scala 1845:39]
  wire  _GEN_6944 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6625; // @[lut_35.scala 1834:74 lut_35.scala 1846:39]
  wire  _GEN_6945 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6626; // @[lut_35.scala 1834:74 lut_35.scala 1847:39]
  wire  _GEN_6946 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6627; // @[lut_35.scala 1834:74 lut_35.scala 1848:39]
  wire  _GEN_6947 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6628; // @[lut_35.scala 1834:74 lut_35.scala 1849:39]
  wire  _GEN_6948 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6629; // @[lut_35.scala 1834:74 lut_35.scala 1850:39]
  wire  _GEN_6949 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6630; // @[lut_35.scala 1834:74 lut_35.scala 1851:39]
  wire  _GEN_6950 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6631; // @[lut_35.scala 1834:74 lut_35.scala 1852:39]
  wire  _GEN_6951 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6632; // @[lut_35.scala 1834:74 lut_35.scala 1853:39]
  wire  _GEN_6952 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6633; // @[lut_35.scala 1834:74 lut_35.scala 1854:39]
  wire  _GEN_6953 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6634; // @[lut_35.scala 1834:74 lut_35.scala 1855:39]
  wire  _GEN_6954 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6635; // @[lut_35.scala 1834:74 lut_35.scala 1856:39]
  wire  _GEN_6955 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6636; // @[lut_35.scala 1834:74 lut_35.scala 1857:39]
  wire  _GEN_6956 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6637; // @[lut_35.scala 1834:74 lut_35.scala 1858:39]
  wire  _GEN_6957 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6638; // @[lut_35.scala 1834:74 lut_35.scala 1859:39]
  wire  _GEN_6958 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6639; // @[lut_35.scala 1834:74 lut_35.scala 1860:39]
  wire  _GEN_6959 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6640; // @[lut_35.scala 1834:74 lut_35.scala 1861:39]
  wire  _GEN_6960 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6641; // @[lut_35.scala 1834:74 lut_35.scala 1862:39]
  wire  _GEN_6961 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6642; // @[lut_35.scala 1834:74 lut_35.scala 1863:39]
  wire  _GEN_6962 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6643; // @[lut_35.scala 1834:74 lut_35.scala 1864:39]
  wire  _GEN_6963 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6644; // @[lut_35.scala 1834:74 lut_35.scala 1865:39]
  wire  _GEN_6964 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6645; // @[lut_35.scala 1834:74 lut_35.scala 1866:39]
  wire  _GEN_6965 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid | _GEN_6646; // @[lut_35.scala 1834:74 lut_35.scala 1867:39]
  wire  _GEN_6966 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6647; // @[lut_35.scala 1834:74 lut_35.scala 1868:39]
  wire  _GEN_6967 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6648; // @[lut_35.scala 1834:74 lut_35.scala 1869:39]
  wire  _GEN_6968 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid | _GEN_6649; // @[lut_35.scala 1834:74 lut_35.scala 1870:34]
  wire  _GEN_6972 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1834:74 lut_35.scala 177:26 lut_35.scala 1872:27]
  wire  _GEN_6975 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6653; // @[lut_35.scala 1834:74 lut_35.scala 177:26]
  wire  _GEN_6978 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6656; // @[lut_35.scala 1834:74 lut_35.scala 177:26]
  wire  _GEN_6986 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6664; // @[lut_35.scala 1834:74 lut_35.scala 177:26]
  wire  _GEN_6993 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6671; // @[lut_35.scala 1834:74 lut_35.scala 177:26]
  wire  _GEN_7001 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6679; // @[lut_35.scala 1834:74 lut_35.scala 177:26]
  wire  _GEN_7009 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6687; // @[lut_35.scala 1834:74 lut_35.scala 177:26]
  wire  _GEN_7017 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6695; // @[lut_35.scala 1834:74 lut_35.scala 177:26]
  wire  _GEN_7025 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6703; // @[lut_35.scala 1834:74 lut_35.scala 177:26]
  wire  _GEN_7033 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6711; // @[lut_35.scala 1834:74 lut_35.scala 177:26]
  wire  _GEN_7041 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6719; // @[lut_35.scala 1834:74 lut_35.scala 177:26]
  wire  _GEN_7049 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6727; // @[lut_35.scala 1834:74 lut_35.scala 177:26]
  wire  _GEN_7057 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6735; // @[lut_35.scala 1834:74 lut_35.scala 177:26]
  wire  _GEN_7065 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6743; // @[lut_35.scala 1834:74 lut_35.scala 177:26]
  wire  _GEN_7073 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6751; // @[lut_35.scala 1834:74 lut_35.scala 177:26]
  wire  _GEN_7081 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6759; // @[lut_35.scala 1834:74 lut_35.scala 177:26]
  wire  _GEN_7089 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6767; // @[lut_35.scala 1834:74 lut_35.scala 177:26]
  wire  _GEN_7097 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6775; // @[lut_35.scala 1834:74 lut_35.scala 177:26]
  wire  _GEN_7105 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6783; // @[lut_35.scala 1834:74 lut_35.scala 177:26]
  wire  _GEN_7113 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6791; // @[lut_35.scala 1834:74 lut_35.scala 177:26]
  wire  _GEN_7121 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6799; // @[lut_35.scala 1834:74 lut_35.scala 177:26]
  wire  _GEN_7129 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6807; // @[lut_35.scala 1834:74 lut_35.scala 177:26]
  wire  _GEN_7137 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6815; // @[lut_35.scala 1834:74 lut_35.scala 177:26]
  wire  _GEN_7145 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6823; // @[lut_35.scala 1834:74 lut_35.scala 177:26]
  wire  _GEN_7153 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6831; // @[lut_35.scala 1834:74 lut_35.scala 177:26]
  wire  _GEN_7161 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6839; // @[lut_35.scala 1834:74 lut_35.scala 177:26]
  wire  _GEN_7169 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6847; // @[lut_35.scala 1834:74 lut_35.scala 177:26]
  wire  _GEN_7177 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6855; // @[lut_35.scala 1834:74 lut_35.scala 177:26]
  wire  _GEN_7185 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6863; // @[lut_35.scala 1834:74 lut_35.scala 177:26]
  wire  _GEN_7193 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6871; // @[lut_35.scala 1834:74 lut_35.scala 177:26]
  wire  _GEN_7201 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6879; // @[lut_35.scala 1834:74 lut_35.scala 177:26]
  wire  _GEN_7209 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6887; // @[lut_35.scala 1834:74 lut_35.scala 177:26]
  wire  _GEN_7217 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6895; // @[lut_35.scala 1834:74 lut_35.scala 177:26]
  wire  _GEN_7225 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6903; // @[lut_35.scala 1834:74 lut_35.scala 177:26]
  wire  _GEN_7233 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6911; // @[lut_35.scala 1834:74 lut_35.scala 177:26]
  wire  _GEN_7236 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6646; // @[lut_35.scala 1834:74 lut_35.scala 177:26]
  wire  _GEN_7241 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6919; // @[lut_35.scala 1834:74 lut_35.scala 177:26]
  wire  _GEN_7244 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6922; // @[lut_35.scala 1834:74 lut_35.scala 177:26]
  wire  _GEN_7249 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6927; // @[lut_35.scala 1834:74 lut_35.scala 177:26]
  wire  _GEN_7252 = LUT_mem_MPORT_207_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6930; // @[lut_35.scala 1834:74 lut_35.scala 177:26]
  wire  _GEN_7255 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6933; // @[lut_35.scala 1796:74 lut_35.scala 1797:38]
  wire  _GEN_7256 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6934; // @[lut_35.scala 1796:74 lut_35.scala 1798:38]
  wire  _GEN_7257 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6935; // @[lut_35.scala 1796:74 lut_35.scala 1799:38]
  wire  _GEN_7258 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6936; // @[lut_35.scala 1796:74 lut_35.scala 1800:38]
  wire  _GEN_7259 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6937; // @[lut_35.scala 1796:74 lut_35.scala 1801:38]
  wire  _GEN_7260 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6938; // @[lut_35.scala 1796:74 lut_35.scala 1802:38]
  wire  _GEN_7261 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6939; // @[lut_35.scala 1796:74 lut_35.scala 1803:38]
  wire  _GEN_7262 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6940; // @[lut_35.scala 1796:74 lut_35.scala 1804:38]
  wire  _GEN_7263 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6941; // @[lut_35.scala 1796:74 lut_35.scala 1805:38]
  wire  _GEN_7264 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6942; // @[lut_35.scala 1796:74 lut_35.scala 1806:38]
  wire  _GEN_7265 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6943; // @[lut_35.scala 1796:74 lut_35.scala 1807:39]
  wire  _GEN_7266 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6944; // @[lut_35.scala 1796:74 lut_35.scala 1808:39]
  wire  _GEN_7267 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6945; // @[lut_35.scala 1796:74 lut_35.scala 1809:39]
  wire  _GEN_7268 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6946; // @[lut_35.scala 1796:74 lut_35.scala 1810:39]
  wire  _GEN_7269 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6947; // @[lut_35.scala 1796:74 lut_35.scala 1811:39]
  wire  _GEN_7270 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6948; // @[lut_35.scala 1796:74 lut_35.scala 1812:39]
  wire  _GEN_7271 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6949; // @[lut_35.scala 1796:74 lut_35.scala 1813:39]
  wire  _GEN_7272 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6950; // @[lut_35.scala 1796:74 lut_35.scala 1814:39]
  wire  _GEN_7273 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6951; // @[lut_35.scala 1796:74 lut_35.scala 1815:39]
  wire  _GEN_7274 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6952; // @[lut_35.scala 1796:74 lut_35.scala 1816:39]
  wire  _GEN_7275 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6953; // @[lut_35.scala 1796:74 lut_35.scala 1817:39]
  wire  _GEN_7276 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6954; // @[lut_35.scala 1796:74 lut_35.scala 1818:39]
  wire  _GEN_7277 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6955; // @[lut_35.scala 1796:74 lut_35.scala 1819:39]
  wire  _GEN_7278 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6956; // @[lut_35.scala 1796:74 lut_35.scala 1820:39]
  wire  _GEN_7279 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6957; // @[lut_35.scala 1796:74 lut_35.scala 1821:39]
  wire  _GEN_7280 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6958; // @[lut_35.scala 1796:74 lut_35.scala 1822:39]
  wire  _GEN_7281 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6959; // @[lut_35.scala 1796:74 lut_35.scala 1823:39]
  wire  _GEN_7282 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6960; // @[lut_35.scala 1796:74 lut_35.scala 1824:39]
  wire  _GEN_7283 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6961; // @[lut_35.scala 1796:74 lut_35.scala 1825:39]
  wire  _GEN_7284 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6962; // @[lut_35.scala 1796:74 lut_35.scala 1826:39]
  wire  _GEN_7285 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6963; // @[lut_35.scala 1796:74 lut_35.scala 1827:39]
  wire  _GEN_7286 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid | _GEN_6964; // @[lut_35.scala 1796:74 lut_35.scala 1828:39]
  wire  _GEN_7287 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6965; // @[lut_35.scala 1796:74 lut_35.scala 1829:39]
  wire  _GEN_7288 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6966; // @[lut_35.scala 1796:74 lut_35.scala 1830:39]
  wire  _GEN_7289 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6967; // @[lut_35.scala 1796:74 lut_35.scala 1831:39]
  wire  _GEN_7290 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid | _GEN_6968; // @[lut_35.scala 1796:74 lut_35.scala 1832:34]
  wire  _GEN_7294 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1796:74 lut_35.scala 177:26 lut_35.scala 1834:27]
  wire  _GEN_7297 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6972; // @[lut_35.scala 1796:74 lut_35.scala 177:26]
  wire  _GEN_7300 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6975; // @[lut_35.scala 1796:74 lut_35.scala 177:26]
  wire  _GEN_7303 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6978; // @[lut_35.scala 1796:74 lut_35.scala 177:26]
  wire  _GEN_7311 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6986; // @[lut_35.scala 1796:74 lut_35.scala 177:26]
  wire  _GEN_7318 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6993; // @[lut_35.scala 1796:74 lut_35.scala 177:26]
  wire  _GEN_7326 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7001; // @[lut_35.scala 1796:74 lut_35.scala 177:26]
  wire  _GEN_7334 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7009; // @[lut_35.scala 1796:74 lut_35.scala 177:26]
  wire  _GEN_7342 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7017; // @[lut_35.scala 1796:74 lut_35.scala 177:26]
  wire  _GEN_7350 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7025; // @[lut_35.scala 1796:74 lut_35.scala 177:26]
  wire  _GEN_7358 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7033; // @[lut_35.scala 1796:74 lut_35.scala 177:26]
  wire  _GEN_7366 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7041; // @[lut_35.scala 1796:74 lut_35.scala 177:26]
  wire  _GEN_7374 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7049; // @[lut_35.scala 1796:74 lut_35.scala 177:26]
  wire  _GEN_7382 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7057; // @[lut_35.scala 1796:74 lut_35.scala 177:26]
  wire  _GEN_7390 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7065; // @[lut_35.scala 1796:74 lut_35.scala 177:26]
  wire  _GEN_7398 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7073; // @[lut_35.scala 1796:74 lut_35.scala 177:26]
  wire  _GEN_7406 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7081; // @[lut_35.scala 1796:74 lut_35.scala 177:26]
  wire  _GEN_7414 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7089; // @[lut_35.scala 1796:74 lut_35.scala 177:26]
  wire  _GEN_7422 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7097; // @[lut_35.scala 1796:74 lut_35.scala 177:26]
  wire  _GEN_7430 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7105; // @[lut_35.scala 1796:74 lut_35.scala 177:26]
  wire  _GEN_7438 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7113; // @[lut_35.scala 1796:74 lut_35.scala 177:26]
  wire  _GEN_7446 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7121; // @[lut_35.scala 1796:74 lut_35.scala 177:26]
  wire  _GEN_7454 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7129; // @[lut_35.scala 1796:74 lut_35.scala 177:26]
  wire  _GEN_7462 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7137; // @[lut_35.scala 1796:74 lut_35.scala 177:26]
  wire  _GEN_7470 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7145; // @[lut_35.scala 1796:74 lut_35.scala 177:26]
  wire  _GEN_7478 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7153; // @[lut_35.scala 1796:74 lut_35.scala 177:26]
  wire  _GEN_7486 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7161; // @[lut_35.scala 1796:74 lut_35.scala 177:26]
  wire  _GEN_7494 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7169; // @[lut_35.scala 1796:74 lut_35.scala 177:26]
  wire  _GEN_7502 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7177; // @[lut_35.scala 1796:74 lut_35.scala 177:26]
  wire  _GEN_7510 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7185; // @[lut_35.scala 1796:74 lut_35.scala 177:26]
  wire  _GEN_7518 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7193; // @[lut_35.scala 1796:74 lut_35.scala 177:26]
  wire  _GEN_7526 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7201; // @[lut_35.scala 1796:74 lut_35.scala 177:26]
  wire  _GEN_7534 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7209; // @[lut_35.scala 1796:74 lut_35.scala 177:26]
  wire  _GEN_7542 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7217; // @[lut_35.scala 1796:74 lut_35.scala 177:26]
  wire  _GEN_7550 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7225; // @[lut_35.scala 1796:74 lut_35.scala 177:26]
  wire  _GEN_7553 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_6964; // @[lut_35.scala 1796:74 lut_35.scala 177:26]
  wire  _GEN_7558 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7233; // @[lut_35.scala 1796:74 lut_35.scala 177:26]
  wire  _GEN_7561 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7236; // @[lut_35.scala 1796:74 lut_35.scala 177:26]
  wire  _GEN_7566 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7241; // @[lut_35.scala 1796:74 lut_35.scala 177:26]
  wire  _GEN_7569 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7244; // @[lut_35.scala 1796:74 lut_35.scala 177:26]
  wire  _GEN_7574 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7249; // @[lut_35.scala 1796:74 lut_35.scala 177:26]
  wire  _GEN_7577 = LUT_mem_MPORT_206_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7252; // @[lut_35.scala 1796:74 lut_35.scala 177:26]
  wire  _GEN_7580 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7255; // @[lut_35.scala 1758:74 lut_35.scala 1759:38]
  wire  _GEN_7581 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7256; // @[lut_35.scala 1758:74 lut_35.scala 1760:38]
  wire  _GEN_7582 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7257; // @[lut_35.scala 1758:74 lut_35.scala 1761:38]
  wire  _GEN_7583 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7258; // @[lut_35.scala 1758:74 lut_35.scala 1762:38]
  wire  _GEN_7584 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7259; // @[lut_35.scala 1758:74 lut_35.scala 1763:38]
  wire  _GEN_7585 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7260; // @[lut_35.scala 1758:74 lut_35.scala 1764:38]
  wire  _GEN_7586 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7261; // @[lut_35.scala 1758:74 lut_35.scala 1765:38]
  wire  _GEN_7587 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7262; // @[lut_35.scala 1758:74 lut_35.scala 1766:38]
  wire  _GEN_7588 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7263; // @[lut_35.scala 1758:74 lut_35.scala 1767:38]
  wire  _GEN_7589 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7264; // @[lut_35.scala 1758:74 lut_35.scala 1768:38]
  wire  _GEN_7590 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7265; // @[lut_35.scala 1758:74 lut_35.scala 1769:39]
  wire  _GEN_7591 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7266; // @[lut_35.scala 1758:74 lut_35.scala 1770:39]
  wire  _GEN_7592 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7267; // @[lut_35.scala 1758:74 lut_35.scala 1771:39]
  wire  _GEN_7593 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7268; // @[lut_35.scala 1758:74 lut_35.scala 1772:39]
  wire  _GEN_7594 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7269; // @[lut_35.scala 1758:74 lut_35.scala 1773:39]
  wire  _GEN_7595 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7270; // @[lut_35.scala 1758:74 lut_35.scala 1774:39]
  wire  _GEN_7596 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7271; // @[lut_35.scala 1758:74 lut_35.scala 1775:39]
  wire  _GEN_7597 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7272; // @[lut_35.scala 1758:74 lut_35.scala 1776:39]
  wire  _GEN_7598 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7273; // @[lut_35.scala 1758:74 lut_35.scala 1777:39]
  wire  _GEN_7599 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7274; // @[lut_35.scala 1758:74 lut_35.scala 1778:39]
  wire  _GEN_7600 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7275; // @[lut_35.scala 1758:74 lut_35.scala 1779:39]
  wire  _GEN_7601 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7276; // @[lut_35.scala 1758:74 lut_35.scala 1780:39]
  wire  _GEN_7602 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7277; // @[lut_35.scala 1758:74 lut_35.scala 1781:39]
  wire  _GEN_7603 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7278; // @[lut_35.scala 1758:74 lut_35.scala 1782:39]
  wire  _GEN_7604 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7279; // @[lut_35.scala 1758:74 lut_35.scala 1783:39]
  wire  _GEN_7605 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7280; // @[lut_35.scala 1758:74 lut_35.scala 1784:39]
  wire  _GEN_7606 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7281; // @[lut_35.scala 1758:74 lut_35.scala 1785:39]
  wire  _GEN_7607 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7282; // @[lut_35.scala 1758:74 lut_35.scala 1786:39]
  wire  _GEN_7608 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7283; // @[lut_35.scala 1758:74 lut_35.scala 1787:39]
  wire  _GEN_7609 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7284; // @[lut_35.scala 1758:74 lut_35.scala 1788:39]
  wire  _GEN_7610 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid | _GEN_7285; // @[lut_35.scala 1758:74 lut_35.scala 1789:39]
  wire  _GEN_7611 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7286; // @[lut_35.scala 1758:74 lut_35.scala 1790:39]
  wire  _GEN_7612 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7287; // @[lut_35.scala 1758:74 lut_35.scala 1791:39]
  wire  _GEN_7613 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7288; // @[lut_35.scala 1758:74 lut_35.scala 1792:39]
  wire  _GEN_7614 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7289; // @[lut_35.scala 1758:74 lut_35.scala 1793:39]
  wire  _GEN_7615 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid | _GEN_7290; // @[lut_35.scala 1758:74 lut_35.scala 1794:34]
  wire  _GEN_7619 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1758:74 lut_35.scala 177:26 lut_35.scala 1796:27]
  wire  _GEN_7622 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7294; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7625 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7297; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7628 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7300; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7631 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7303; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7639 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7311; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7646 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7318; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7654 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7326; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7662 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7334; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7670 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7342; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7678 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7350; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7686 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7358; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7694 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7366; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7702 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7374; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7710 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7382; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7718 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7390; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7726 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7398; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7734 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7406; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7742 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7414; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7750 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7422; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7758 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7430; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7766 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7438; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7774 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7446; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7782 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7454; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7790 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7462; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7798 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7470; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7806 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7478; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7814 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7486; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7822 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7494; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7830 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7502; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7838 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7510; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7846 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7518; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7854 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7526; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7862 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7534; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7870 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7542; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7873 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7285; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7878 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7550; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7881 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7553; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7886 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7558; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7889 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7561; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7894 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7566; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7897 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7569; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7902 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7574; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7905 = LUT_mem_MPORT_205_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7577; // @[lut_35.scala 1758:74 lut_35.scala 177:26]
  wire  _GEN_7908 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7580; // @[lut_35.scala 1720:74 lut_35.scala 1721:38]
  wire  _GEN_7909 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7581; // @[lut_35.scala 1720:74 lut_35.scala 1722:38]
  wire  _GEN_7910 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7582; // @[lut_35.scala 1720:74 lut_35.scala 1723:38]
  wire  _GEN_7911 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7583; // @[lut_35.scala 1720:74 lut_35.scala 1724:38]
  wire  _GEN_7912 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7584; // @[lut_35.scala 1720:74 lut_35.scala 1725:38]
  wire  _GEN_7913 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7585; // @[lut_35.scala 1720:74 lut_35.scala 1726:38]
  wire  _GEN_7914 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7586; // @[lut_35.scala 1720:74 lut_35.scala 1727:38]
  wire  _GEN_7915 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7587; // @[lut_35.scala 1720:74 lut_35.scala 1728:38]
  wire  _GEN_7916 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7588; // @[lut_35.scala 1720:74 lut_35.scala 1729:38]
  wire  _GEN_7917 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7589; // @[lut_35.scala 1720:74 lut_35.scala 1730:38]
  wire  _GEN_7918 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7590; // @[lut_35.scala 1720:74 lut_35.scala 1731:39]
  wire  _GEN_7919 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7591; // @[lut_35.scala 1720:74 lut_35.scala 1732:39]
  wire  _GEN_7920 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7592; // @[lut_35.scala 1720:74 lut_35.scala 1733:39]
  wire  _GEN_7921 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7593; // @[lut_35.scala 1720:74 lut_35.scala 1734:39]
  wire  _GEN_7922 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7594; // @[lut_35.scala 1720:74 lut_35.scala 1735:39]
  wire  _GEN_7923 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7595; // @[lut_35.scala 1720:74 lut_35.scala 1736:39]
  wire  _GEN_7924 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7596; // @[lut_35.scala 1720:74 lut_35.scala 1737:39]
  wire  _GEN_7925 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7597; // @[lut_35.scala 1720:74 lut_35.scala 1738:39]
  wire  _GEN_7926 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7598; // @[lut_35.scala 1720:74 lut_35.scala 1739:39]
  wire  _GEN_7927 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7599; // @[lut_35.scala 1720:74 lut_35.scala 1740:39]
  wire  _GEN_7928 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7600; // @[lut_35.scala 1720:74 lut_35.scala 1741:39]
  wire  _GEN_7929 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7601; // @[lut_35.scala 1720:74 lut_35.scala 1742:39]
  wire  _GEN_7930 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7602; // @[lut_35.scala 1720:74 lut_35.scala 1743:39]
  wire  _GEN_7931 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7603; // @[lut_35.scala 1720:74 lut_35.scala 1744:39]
  wire  _GEN_7932 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7604; // @[lut_35.scala 1720:74 lut_35.scala 1745:39]
  wire  _GEN_7933 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7605; // @[lut_35.scala 1720:74 lut_35.scala 1746:39]
  wire  _GEN_7934 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7606; // @[lut_35.scala 1720:74 lut_35.scala 1747:39]
  wire  _GEN_7935 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7607; // @[lut_35.scala 1720:74 lut_35.scala 1748:39]
  wire  _GEN_7936 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7608; // @[lut_35.scala 1720:74 lut_35.scala 1749:39]
  wire  _GEN_7937 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid | _GEN_7609; // @[lut_35.scala 1720:74 lut_35.scala 1750:39]
  wire  _GEN_7938 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7610; // @[lut_35.scala 1720:74 lut_35.scala 1751:39]
  wire  _GEN_7939 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7611; // @[lut_35.scala 1720:74 lut_35.scala 1752:39]
  wire  _GEN_7940 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7612; // @[lut_35.scala 1720:74 lut_35.scala 1753:39]
  wire  _GEN_7941 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7613; // @[lut_35.scala 1720:74 lut_35.scala 1754:39]
  wire  _GEN_7942 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7614; // @[lut_35.scala 1720:74 lut_35.scala 1755:39]
  wire  _GEN_7943 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid | _GEN_7615; // @[lut_35.scala 1720:74 lut_35.scala 1756:34]
  wire  _GEN_7947 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1720:74 lut_35.scala 177:26 lut_35.scala 1758:27]
  wire  _GEN_7950 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7619; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_7953 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7622; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_7956 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7625; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_7959 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7628; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_7962 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7631; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_7970 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7639; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_7977 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7646; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_7985 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7654; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_7993 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7662; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_8001 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7670; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_8009 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7678; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_8017 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7686; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_8025 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7694; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_8033 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7702; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_8041 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7710; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_8049 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7718; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_8057 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7726; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_8065 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7734; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_8073 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7742; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_8081 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7750; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_8089 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7758; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_8097 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7766; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_8105 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7774; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_8113 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7782; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_8121 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7790; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_8129 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7798; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_8137 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7806; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_8145 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7814; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_8153 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7822; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_8161 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7830; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_8169 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7838; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_8177 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7846; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_8185 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7854; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_8193 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7862; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_8196 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7609; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_8201 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7870; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_8204 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7873; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_8209 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7878; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_8212 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7881; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_8217 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7886; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_8220 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7889; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_8225 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7894; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_8228 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7897; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_8233 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7902; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_8236 = LUT_mem_MPORT_204_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7905; // @[lut_35.scala 1720:74 lut_35.scala 177:26]
  wire  _GEN_8239 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7908; // @[lut_35.scala 1682:74 lut_35.scala 1683:38]
  wire  _GEN_8240 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7909; // @[lut_35.scala 1682:74 lut_35.scala 1684:38]
  wire  _GEN_8241 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7910; // @[lut_35.scala 1682:74 lut_35.scala 1685:38]
  wire  _GEN_8242 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7911; // @[lut_35.scala 1682:74 lut_35.scala 1686:38]
  wire  _GEN_8243 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7912; // @[lut_35.scala 1682:74 lut_35.scala 1687:38]
  wire  _GEN_8244 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7913; // @[lut_35.scala 1682:74 lut_35.scala 1688:38]
  wire  _GEN_8245 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7914; // @[lut_35.scala 1682:74 lut_35.scala 1689:38]
  wire  _GEN_8246 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7915; // @[lut_35.scala 1682:74 lut_35.scala 1690:38]
  wire  _GEN_8247 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7916; // @[lut_35.scala 1682:74 lut_35.scala 1691:38]
  wire  _GEN_8248 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7917; // @[lut_35.scala 1682:74 lut_35.scala 1692:38]
  wire  _GEN_8249 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7918; // @[lut_35.scala 1682:74 lut_35.scala 1693:39]
  wire  _GEN_8250 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7919; // @[lut_35.scala 1682:74 lut_35.scala 1694:39]
  wire  _GEN_8251 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7920; // @[lut_35.scala 1682:74 lut_35.scala 1695:39]
  wire  _GEN_8252 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7921; // @[lut_35.scala 1682:74 lut_35.scala 1696:39]
  wire  _GEN_8253 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7922; // @[lut_35.scala 1682:74 lut_35.scala 1697:39]
  wire  _GEN_8254 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7923; // @[lut_35.scala 1682:74 lut_35.scala 1698:39]
  wire  _GEN_8255 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7924; // @[lut_35.scala 1682:74 lut_35.scala 1699:39]
  wire  _GEN_8256 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7925; // @[lut_35.scala 1682:74 lut_35.scala 1700:39]
  wire  _GEN_8257 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7926; // @[lut_35.scala 1682:74 lut_35.scala 1701:39]
  wire  _GEN_8258 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7927; // @[lut_35.scala 1682:74 lut_35.scala 1702:39]
  wire  _GEN_8259 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7928; // @[lut_35.scala 1682:74 lut_35.scala 1703:39]
  wire  _GEN_8260 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7929; // @[lut_35.scala 1682:74 lut_35.scala 1704:39]
  wire  _GEN_8261 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7930; // @[lut_35.scala 1682:74 lut_35.scala 1705:39]
  wire  _GEN_8262 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7931; // @[lut_35.scala 1682:74 lut_35.scala 1706:39]
  wire  _GEN_8263 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7932; // @[lut_35.scala 1682:74 lut_35.scala 1707:39]
  wire  _GEN_8264 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7933; // @[lut_35.scala 1682:74 lut_35.scala 1708:39]
  wire  _GEN_8265 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7934; // @[lut_35.scala 1682:74 lut_35.scala 1709:39]
  wire  _GEN_8266 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7935; // @[lut_35.scala 1682:74 lut_35.scala 1710:39]
  wire  _GEN_8267 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid | _GEN_7936; // @[lut_35.scala 1682:74 lut_35.scala 1711:39]
  wire  _GEN_8268 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7937; // @[lut_35.scala 1682:74 lut_35.scala 1712:39]
  wire  _GEN_8269 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7938; // @[lut_35.scala 1682:74 lut_35.scala 1713:39]
  wire  _GEN_8270 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7939; // @[lut_35.scala 1682:74 lut_35.scala 1714:39]
  wire  _GEN_8271 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7940; // @[lut_35.scala 1682:74 lut_35.scala 1715:39]
  wire  _GEN_8272 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7941; // @[lut_35.scala 1682:74 lut_35.scala 1716:39]
  wire  _GEN_8273 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7942; // @[lut_35.scala 1682:74 lut_35.scala 1717:39]
  wire  _GEN_8274 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid | _GEN_7943; // @[lut_35.scala 1682:74 lut_35.scala 1718:34]
  wire  _GEN_8278 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1682:74 lut_35.scala 177:26 lut_35.scala 1720:27]
  wire  _GEN_8281 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7947; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8284 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7950; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8287 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7953; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8290 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7956; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8293 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7959; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8296 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7962; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8304 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7970; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8311 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7977; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8319 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7985; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8327 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7993; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8335 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8001; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8343 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8009; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8351 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8017; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8359 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8025; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8367 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8033; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8375 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8041; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8383 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8049; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8391 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8057; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8399 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8065; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8407 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8073; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8415 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8081; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8423 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8089; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8431 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8097; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8439 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8105; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8447 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8113; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8455 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8121; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8463 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8129; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8471 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8137; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8479 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8145; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8487 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8153; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8495 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8161; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8503 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8169; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8511 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8177; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8519 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8185; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8522 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_7936; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8527 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8193; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8530 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8196; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8535 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8201; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8538 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8204; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8543 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8209; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8546 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8212; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8551 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8217; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8554 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8220; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8559 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8225; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8562 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8228; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8567 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8233; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8570 = LUT_mem_MPORT_203_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8236; // @[lut_35.scala 1682:74 lut_35.scala 177:26]
  wire  _GEN_8573 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8239; // @[lut_35.scala 1644:74 lut_35.scala 1645:38]
  wire  _GEN_8574 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8240; // @[lut_35.scala 1644:74 lut_35.scala 1646:38]
  wire  _GEN_8575 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8241; // @[lut_35.scala 1644:74 lut_35.scala 1647:38]
  wire  _GEN_8576 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8242; // @[lut_35.scala 1644:74 lut_35.scala 1648:38]
  wire  _GEN_8577 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8243; // @[lut_35.scala 1644:74 lut_35.scala 1649:38]
  wire  _GEN_8578 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8244; // @[lut_35.scala 1644:74 lut_35.scala 1650:38]
  wire  _GEN_8579 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8245; // @[lut_35.scala 1644:74 lut_35.scala 1651:38]
  wire  _GEN_8580 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8246; // @[lut_35.scala 1644:74 lut_35.scala 1652:38]
  wire  _GEN_8581 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8247; // @[lut_35.scala 1644:74 lut_35.scala 1653:38]
  wire  _GEN_8582 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8248; // @[lut_35.scala 1644:74 lut_35.scala 1654:38]
  wire  _GEN_8583 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8249; // @[lut_35.scala 1644:74 lut_35.scala 1655:39]
  wire  _GEN_8584 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8250; // @[lut_35.scala 1644:74 lut_35.scala 1656:39]
  wire  _GEN_8585 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8251; // @[lut_35.scala 1644:74 lut_35.scala 1657:39]
  wire  _GEN_8586 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8252; // @[lut_35.scala 1644:74 lut_35.scala 1658:39]
  wire  _GEN_8587 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8253; // @[lut_35.scala 1644:74 lut_35.scala 1659:39]
  wire  _GEN_8588 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8254; // @[lut_35.scala 1644:74 lut_35.scala 1660:39]
  wire  _GEN_8589 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8255; // @[lut_35.scala 1644:74 lut_35.scala 1661:39]
  wire  _GEN_8590 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8256; // @[lut_35.scala 1644:74 lut_35.scala 1662:39]
  wire  _GEN_8591 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8257; // @[lut_35.scala 1644:74 lut_35.scala 1663:39]
  wire  _GEN_8592 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8258; // @[lut_35.scala 1644:74 lut_35.scala 1664:39]
  wire  _GEN_8593 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8259; // @[lut_35.scala 1644:74 lut_35.scala 1665:39]
  wire  _GEN_8594 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8260; // @[lut_35.scala 1644:74 lut_35.scala 1666:39]
  wire  _GEN_8595 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8261; // @[lut_35.scala 1644:74 lut_35.scala 1667:39]
  wire  _GEN_8596 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8262; // @[lut_35.scala 1644:74 lut_35.scala 1668:39]
  wire  _GEN_8597 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8263; // @[lut_35.scala 1644:74 lut_35.scala 1669:39]
  wire  _GEN_8598 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8264; // @[lut_35.scala 1644:74 lut_35.scala 1670:39]
  wire  _GEN_8599 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8265; // @[lut_35.scala 1644:74 lut_35.scala 1671:39]
  wire  _GEN_8600 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid | _GEN_8266; // @[lut_35.scala 1644:74 lut_35.scala 1672:39]
  wire  _GEN_8601 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8267; // @[lut_35.scala 1644:74 lut_35.scala 1673:39]
  wire  _GEN_8602 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8268; // @[lut_35.scala 1644:74 lut_35.scala 1674:39]
  wire  _GEN_8603 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8269; // @[lut_35.scala 1644:74 lut_35.scala 1675:39]
  wire  _GEN_8604 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8270; // @[lut_35.scala 1644:74 lut_35.scala 1676:39]
  wire  _GEN_8605 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8271; // @[lut_35.scala 1644:74 lut_35.scala 1677:39]
  wire  _GEN_8606 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8272; // @[lut_35.scala 1644:74 lut_35.scala 1678:39]
  wire  _GEN_8607 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8273; // @[lut_35.scala 1644:74 lut_35.scala 1679:39]
  wire  _GEN_8608 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid | _GEN_8274; // @[lut_35.scala 1644:74 lut_35.scala 1680:34]
  wire  _GEN_8612 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1644:74 lut_35.scala 177:26 lut_35.scala 1682:27]
  wire  _GEN_8615 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8278; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8618 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8281; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8621 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8284; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8624 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8287; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8627 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8290; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8630 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8293; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8633 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8296; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8641 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8304; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8648 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8311; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8656 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8319; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8664 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8327; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8672 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8335; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8680 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8343; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8688 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8351; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8696 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8359; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8704 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8367; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8712 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8375; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8720 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8383; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8728 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8391; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8736 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8399; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8744 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8407; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8752 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8415; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8760 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8423; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8768 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8431; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8776 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8439; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8784 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8447; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8792 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8455; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8800 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8463; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8808 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8471; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8816 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8479; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8824 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8487; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8832 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8495; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8840 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8503; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8848 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8511; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8851 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8266; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8856 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8519; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8859 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8522; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8864 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8527; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8867 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8530; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8872 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8535; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8875 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8538; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8880 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8543; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8883 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8546; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8888 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8551; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8891 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8554; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8896 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8559; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8899 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8562; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8904 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8567; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8907 = LUT_mem_MPORT_202_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8570; // @[lut_35.scala 1644:74 lut_35.scala 177:26]
  wire  _GEN_8910 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8573; // @[lut_35.scala 1606:74 lut_35.scala 1607:38]
  wire  _GEN_8911 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8574; // @[lut_35.scala 1606:74 lut_35.scala 1608:38]
  wire  _GEN_8912 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8575; // @[lut_35.scala 1606:74 lut_35.scala 1609:38]
  wire  _GEN_8913 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8576; // @[lut_35.scala 1606:74 lut_35.scala 1610:38]
  wire  _GEN_8914 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8577; // @[lut_35.scala 1606:74 lut_35.scala 1611:38]
  wire  _GEN_8915 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8578; // @[lut_35.scala 1606:74 lut_35.scala 1612:38]
  wire  _GEN_8916 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8579; // @[lut_35.scala 1606:74 lut_35.scala 1613:38]
  wire  _GEN_8917 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8580; // @[lut_35.scala 1606:74 lut_35.scala 1614:38]
  wire  _GEN_8918 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8581; // @[lut_35.scala 1606:74 lut_35.scala 1615:38]
  wire  _GEN_8919 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8582; // @[lut_35.scala 1606:74 lut_35.scala 1616:38]
  wire  _GEN_8920 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8583; // @[lut_35.scala 1606:74 lut_35.scala 1617:39]
  wire  _GEN_8921 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8584; // @[lut_35.scala 1606:74 lut_35.scala 1618:39]
  wire  _GEN_8922 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8585; // @[lut_35.scala 1606:74 lut_35.scala 1619:39]
  wire  _GEN_8923 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8586; // @[lut_35.scala 1606:74 lut_35.scala 1620:39]
  wire  _GEN_8924 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8587; // @[lut_35.scala 1606:74 lut_35.scala 1621:39]
  wire  _GEN_8925 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8588; // @[lut_35.scala 1606:74 lut_35.scala 1622:39]
  wire  _GEN_8926 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8589; // @[lut_35.scala 1606:74 lut_35.scala 1623:39]
  wire  _GEN_8927 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8590; // @[lut_35.scala 1606:74 lut_35.scala 1624:39]
  wire  _GEN_8928 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8591; // @[lut_35.scala 1606:74 lut_35.scala 1625:39]
  wire  _GEN_8929 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8592; // @[lut_35.scala 1606:74 lut_35.scala 1626:39]
  wire  _GEN_8930 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8593; // @[lut_35.scala 1606:74 lut_35.scala 1627:39]
  wire  _GEN_8931 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8594; // @[lut_35.scala 1606:74 lut_35.scala 1628:39]
  wire  _GEN_8932 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8595; // @[lut_35.scala 1606:74 lut_35.scala 1629:39]
  wire  _GEN_8933 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8596; // @[lut_35.scala 1606:74 lut_35.scala 1630:39]
  wire  _GEN_8934 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8597; // @[lut_35.scala 1606:74 lut_35.scala 1631:39]
  wire  _GEN_8935 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8598; // @[lut_35.scala 1606:74 lut_35.scala 1632:39]
  wire  _GEN_8936 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid | _GEN_8599; // @[lut_35.scala 1606:74 lut_35.scala 1633:39]
  wire  _GEN_8937 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8600; // @[lut_35.scala 1606:74 lut_35.scala 1634:39]
  wire  _GEN_8938 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8601; // @[lut_35.scala 1606:74 lut_35.scala 1635:39]
  wire  _GEN_8939 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8602; // @[lut_35.scala 1606:74 lut_35.scala 1636:39]
  wire  _GEN_8940 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8603; // @[lut_35.scala 1606:74 lut_35.scala 1637:39]
  wire  _GEN_8941 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8604; // @[lut_35.scala 1606:74 lut_35.scala 1638:39]
  wire  _GEN_8942 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8605; // @[lut_35.scala 1606:74 lut_35.scala 1639:39]
  wire  _GEN_8943 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8606; // @[lut_35.scala 1606:74 lut_35.scala 1640:39]
  wire  _GEN_8944 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8607; // @[lut_35.scala 1606:74 lut_35.scala 1641:39]
  wire  _GEN_8945 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid | _GEN_8608; // @[lut_35.scala 1606:74 lut_35.scala 1642:34]
  wire  _GEN_8949 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1606:74 lut_35.scala 177:26 lut_35.scala 1644:27]
  wire  _GEN_8952 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8612; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_8955 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8615; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_8958 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8618; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_8961 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8621; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_8964 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8624; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_8967 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8627; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_8970 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8630; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_8973 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8633; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_8981 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8641; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_8988 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8648; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_8996 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8656; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_9004 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8664; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_9012 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8672; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_9020 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8680; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_9028 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8688; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_9036 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8696; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_9044 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8704; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_9052 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8712; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_9060 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8720; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_9068 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8728; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_9076 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8736; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_9084 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8744; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_9092 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8752; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_9100 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8760; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_9108 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8768; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_9116 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8776; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_9124 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8784; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_9132 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8792; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_9140 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8800; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_9148 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8808; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_9156 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8816; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_9164 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8824; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_9172 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8832; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_9180 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8840; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_9183 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8599; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_9188 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8848; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_9191 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8851; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_9196 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8856; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_9199 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8859; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_9204 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8864; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_9207 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8867; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_9212 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8872; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_9215 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8875; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_9220 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8880; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_9223 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8883; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_9228 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8888; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_9231 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8891; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_9236 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8896; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_9239 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8899; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_9244 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8904; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_9247 = LUT_mem_MPORT_201_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8907; // @[lut_35.scala 1606:74 lut_35.scala 177:26]
  wire  _GEN_9250 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8910; // @[lut_35.scala 1568:74 lut_35.scala 1569:38]
  wire  _GEN_9251 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8911; // @[lut_35.scala 1568:74 lut_35.scala 1570:38]
  wire  _GEN_9252 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8912; // @[lut_35.scala 1568:74 lut_35.scala 1571:38]
  wire  _GEN_9253 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8913; // @[lut_35.scala 1568:74 lut_35.scala 1572:38]
  wire  _GEN_9254 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8914; // @[lut_35.scala 1568:74 lut_35.scala 1573:38]
  wire  _GEN_9255 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8915; // @[lut_35.scala 1568:74 lut_35.scala 1574:38]
  wire  _GEN_9256 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8916; // @[lut_35.scala 1568:74 lut_35.scala 1575:38]
  wire  _GEN_9257 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8917; // @[lut_35.scala 1568:74 lut_35.scala 1576:38]
  wire  _GEN_9258 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8918; // @[lut_35.scala 1568:74 lut_35.scala 1577:38]
  wire  _GEN_9259 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8919; // @[lut_35.scala 1568:74 lut_35.scala 1578:38]
  wire  _GEN_9260 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8920; // @[lut_35.scala 1568:74 lut_35.scala 1579:39]
  wire  _GEN_9261 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8921; // @[lut_35.scala 1568:74 lut_35.scala 1580:39]
  wire  _GEN_9262 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8922; // @[lut_35.scala 1568:74 lut_35.scala 1581:39]
  wire  _GEN_9263 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8923; // @[lut_35.scala 1568:74 lut_35.scala 1582:39]
  wire  _GEN_9264 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8924; // @[lut_35.scala 1568:74 lut_35.scala 1583:39]
  wire  _GEN_9265 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8925; // @[lut_35.scala 1568:74 lut_35.scala 1584:39]
  wire  _GEN_9266 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8926; // @[lut_35.scala 1568:74 lut_35.scala 1585:39]
  wire  _GEN_9267 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8927; // @[lut_35.scala 1568:74 lut_35.scala 1586:39]
  wire  _GEN_9268 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8928; // @[lut_35.scala 1568:74 lut_35.scala 1587:39]
  wire  _GEN_9269 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8929; // @[lut_35.scala 1568:74 lut_35.scala 1588:39]
  wire  _GEN_9270 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8930; // @[lut_35.scala 1568:74 lut_35.scala 1589:39]
  wire  _GEN_9271 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8931; // @[lut_35.scala 1568:74 lut_35.scala 1590:39]
  wire  _GEN_9272 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8932; // @[lut_35.scala 1568:74 lut_35.scala 1591:39]
  wire  _GEN_9273 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8933; // @[lut_35.scala 1568:74 lut_35.scala 1592:39]
  wire  _GEN_9274 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8934; // @[lut_35.scala 1568:74 lut_35.scala 1593:39]
  wire  _GEN_9275 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid | _GEN_8935; // @[lut_35.scala 1568:74 lut_35.scala 1594:39]
  wire  _GEN_9276 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8936; // @[lut_35.scala 1568:74 lut_35.scala 1595:39]
  wire  _GEN_9277 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8937; // @[lut_35.scala 1568:74 lut_35.scala 1596:39]
  wire  _GEN_9278 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8938; // @[lut_35.scala 1568:74 lut_35.scala 1597:39]
  wire  _GEN_9279 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8939; // @[lut_35.scala 1568:74 lut_35.scala 1598:39]
  wire  _GEN_9280 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8940; // @[lut_35.scala 1568:74 lut_35.scala 1599:39]
  wire  _GEN_9281 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8941; // @[lut_35.scala 1568:74 lut_35.scala 1600:39]
  wire  _GEN_9282 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8942; // @[lut_35.scala 1568:74 lut_35.scala 1601:39]
  wire  _GEN_9283 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8943; // @[lut_35.scala 1568:74 lut_35.scala 1602:39]
  wire  _GEN_9284 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8944; // @[lut_35.scala 1568:74 lut_35.scala 1603:39]
  wire  _GEN_9285 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid | _GEN_8945; // @[lut_35.scala 1568:74 lut_35.scala 1604:34]
  wire  _GEN_9289 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1568:74 lut_35.scala 177:26 lut_35.scala 1606:27]
  wire  _GEN_9292 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8949; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9295 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8952; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9298 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8955; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9301 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8958; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9304 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8961; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9307 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8964; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9310 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8967; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9313 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8970; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9316 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8973; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9324 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8981; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9331 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8988; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9339 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8996; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9347 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9004; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9355 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9012; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9363 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9020; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9371 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9028; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9379 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9036; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9387 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9044; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9395 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9052; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9403 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9060; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9411 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9068; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9419 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9076; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9427 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9084; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9435 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9092; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9443 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9100; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9451 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9108; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9459 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9116; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9467 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9124; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9475 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9132; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9483 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9140; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9491 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9148; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9499 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9156; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9507 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9164; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9515 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9172; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9518 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_8935; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9523 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9180; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9526 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9183; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9531 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9188; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9534 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9191; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9539 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9196; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9542 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9199; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9547 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9204; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9550 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9207; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9555 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9212; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9558 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9215; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9563 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9220; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9566 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9223; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9571 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9228; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9574 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9231; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9579 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9236; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9582 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9239; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9587 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9244; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9590 = LUT_mem_MPORT_200_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9247; // @[lut_35.scala 1568:74 lut_35.scala 177:26]
  wire  _GEN_9593 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9250; // @[lut_35.scala 1530:74 lut_35.scala 1531:38]
  wire  _GEN_9594 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9251; // @[lut_35.scala 1530:74 lut_35.scala 1532:38]
  wire  _GEN_9595 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9252; // @[lut_35.scala 1530:74 lut_35.scala 1533:38]
  wire  _GEN_9596 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9253; // @[lut_35.scala 1530:74 lut_35.scala 1534:38]
  wire  _GEN_9597 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9254; // @[lut_35.scala 1530:74 lut_35.scala 1535:38]
  wire  _GEN_9598 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9255; // @[lut_35.scala 1530:74 lut_35.scala 1536:38]
  wire  _GEN_9599 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9256; // @[lut_35.scala 1530:74 lut_35.scala 1537:38]
  wire  _GEN_9600 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9257; // @[lut_35.scala 1530:74 lut_35.scala 1538:38]
  wire  _GEN_9601 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9258; // @[lut_35.scala 1530:74 lut_35.scala 1539:38]
  wire  _GEN_9602 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9259; // @[lut_35.scala 1530:74 lut_35.scala 1540:38]
  wire  _GEN_9603 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9260; // @[lut_35.scala 1530:74 lut_35.scala 1541:39]
  wire  _GEN_9604 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9261; // @[lut_35.scala 1530:74 lut_35.scala 1542:39]
  wire  _GEN_9605 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9262; // @[lut_35.scala 1530:74 lut_35.scala 1543:39]
  wire  _GEN_9606 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9263; // @[lut_35.scala 1530:74 lut_35.scala 1544:39]
  wire  _GEN_9607 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9264; // @[lut_35.scala 1530:74 lut_35.scala 1545:39]
  wire  _GEN_9608 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9265; // @[lut_35.scala 1530:74 lut_35.scala 1546:39]
  wire  _GEN_9609 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9266; // @[lut_35.scala 1530:74 lut_35.scala 1547:39]
  wire  _GEN_9610 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9267; // @[lut_35.scala 1530:74 lut_35.scala 1548:39]
  wire  _GEN_9611 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9268; // @[lut_35.scala 1530:74 lut_35.scala 1549:39]
  wire  _GEN_9612 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9269; // @[lut_35.scala 1530:74 lut_35.scala 1550:39]
  wire  _GEN_9613 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9270; // @[lut_35.scala 1530:74 lut_35.scala 1551:39]
  wire  _GEN_9614 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9271; // @[lut_35.scala 1530:74 lut_35.scala 1552:39]
  wire  _GEN_9615 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9272; // @[lut_35.scala 1530:74 lut_35.scala 1553:39]
  wire  _GEN_9616 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9273; // @[lut_35.scala 1530:74 lut_35.scala 1554:39]
  wire  _GEN_9617 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid | _GEN_9274; // @[lut_35.scala 1530:74 lut_35.scala 1555:39]
  wire  _GEN_9618 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9275; // @[lut_35.scala 1530:74 lut_35.scala 1556:39]
  wire  _GEN_9619 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9276; // @[lut_35.scala 1530:74 lut_35.scala 1557:39]
  wire  _GEN_9620 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9277; // @[lut_35.scala 1530:74 lut_35.scala 1558:39]
  wire  _GEN_9621 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9278; // @[lut_35.scala 1530:74 lut_35.scala 1559:39]
  wire  _GEN_9622 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9279; // @[lut_35.scala 1530:74 lut_35.scala 1560:39]
  wire  _GEN_9623 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9280; // @[lut_35.scala 1530:74 lut_35.scala 1561:39]
  wire  _GEN_9624 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9281; // @[lut_35.scala 1530:74 lut_35.scala 1562:39]
  wire  _GEN_9625 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9282; // @[lut_35.scala 1530:74 lut_35.scala 1563:39]
  wire  _GEN_9626 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9283; // @[lut_35.scala 1530:74 lut_35.scala 1564:39]
  wire  _GEN_9627 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9284; // @[lut_35.scala 1530:74 lut_35.scala 1565:39]
  wire  _GEN_9628 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid | _GEN_9285; // @[lut_35.scala 1530:74 lut_35.scala 1566:34]
  wire  _GEN_9632 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1530:74 lut_35.scala 177:26 lut_35.scala 1568:27]
  wire  _GEN_9635 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9289; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9638 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9292; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9641 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9295; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9644 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9298; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9647 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9301; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9650 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9304; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9653 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9307; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9656 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9310; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9659 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9313; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9662 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9316; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9670 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9324; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9677 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9331; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9685 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9339; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9693 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9347; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9701 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9355; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9709 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9363; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9717 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9371; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9725 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9379; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9733 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9387; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9741 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9395; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9749 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9403; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9757 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9411; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9765 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9419; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9773 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9427; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9781 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9435; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9789 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9443; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9797 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9451; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9805 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9459; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9813 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9467; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9821 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9475; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9829 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9483; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9837 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9491; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9845 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9499; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9853 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9507; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9856 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9274; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9861 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9515; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9864 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9518; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9869 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9523; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9872 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9526; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9877 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9531; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9880 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9534; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9885 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9539; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9888 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9542; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9893 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9547; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9896 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9550; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9901 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9555; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9904 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9558; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9909 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9563; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9912 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9566; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9917 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9571; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9920 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9574; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9925 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9579; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9928 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9582; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9933 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9587; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9936 = LUT_mem_MPORT_199_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9590; // @[lut_35.scala 1530:74 lut_35.scala 177:26]
  wire  _GEN_9939 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9593; // @[lut_35.scala 1492:74 lut_35.scala 1493:38]
  wire  _GEN_9940 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9594; // @[lut_35.scala 1492:74 lut_35.scala 1494:38]
  wire  _GEN_9941 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9595; // @[lut_35.scala 1492:74 lut_35.scala 1495:38]
  wire  _GEN_9942 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9596; // @[lut_35.scala 1492:74 lut_35.scala 1496:38]
  wire  _GEN_9943 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9597; // @[lut_35.scala 1492:74 lut_35.scala 1497:38]
  wire  _GEN_9944 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9598; // @[lut_35.scala 1492:74 lut_35.scala 1498:38]
  wire  _GEN_9945 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9599; // @[lut_35.scala 1492:74 lut_35.scala 1499:38]
  wire  _GEN_9946 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9600; // @[lut_35.scala 1492:74 lut_35.scala 1500:38]
  wire  _GEN_9947 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9601; // @[lut_35.scala 1492:74 lut_35.scala 1501:38]
  wire  _GEN_9948 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9602; // @[lut_35.scala 1492:74 lut_35.scala 1502:38]
  wire  _GEN_9949 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9603; // @[lut_35.scala 1492:74 lut_35.scala 1503:39]
  wire  _GEN_9950 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9604; // @[lut_35.scala 1492:74 lut_35.scala 1504:39]
  wire  _GEN_9951 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9605; // @[lut_35.scala 1492:74 lut_35.scala 1505:39]
  wire  _GEN_9952 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9606; // @[lut_35.scala 1492:74 lut_35.scala 1506:39]
  wire  _GEN_9953 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9607; // @[lut_35.scala 1492:74 lut_35.scala 1507:39]
  wire  _GEN_9954 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9608; // @[lut_35.scala 1492:74 lut_35.scala 1508:39]
  wire  _GEN_9955 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9609; // @[lut_35.scala 1492:74 lut_35.scala 1509:39]
  wire  _GEN_9956 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9610; // @[lut_35.scala 1492:74 lut_35.scala 1510:39]
  wire  _GEN_9957 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9611; // @[lut_35.scala 1492:74 lut_35.scala 1511:39]
  wire  _GEN_9958 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9612; // @[lut_35.scala 1492:74 lut_35.scala 1512:39]
  wire  _GEN_9959 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9613; // @[lut_35.scala 1492:74 lut_35.scala 1513:39]
  wire  _GEN_9960 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9614; // @[lut_35.scala 1492:74 lut_35.scala 1514:39]
  wire  _GEN_9961 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9615; // @[lut_35.scala 1492:74 lut_35.scala 1515:39]
  wire  _GEN_9962 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid | _GEN_9616; // @[lut_35.scala 1492:74 lut_35.scala 1516:39]
  wire  _GEN_9963 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9617; // @[lut_35.scala 1492:74 lut_35.scala 1517:39]
  wire  _GEN_9964 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9618; // @[lut_35.scala 1492:74 lut_35.scala 1518:39]
  wire  _GEN_9965 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9619; // @[lut_35.scala 1492:74 lut_35.scala 1519:39]
  wire  _GEN_9966 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9620; // @[lut_35.scala 1492:74 lut_35.scala 1520:39]
  wire  _GEN_9967 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9621; // @[lut_35.scala 1492:74 lut_35.scala 1521:39]
  wire  _GEN_9968 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9622; // @[lut_35.scala 1492:74 lut_35.scala 1522:39]
  wire  _GEN_9969 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9623; // @[lut_35.scala 1492:74 lut_35.scala 1523:39]
  wire  _GEN_9970 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9624; // @[lut_35.scala 1492:74 lut_35.scala 1524:39]
  wire  _GEN_9971 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9625; // @[lut_35.scala 1492:74 lut_35.scala 1525:39]
  wire  _GEN_9972 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9626; // @[lut_35.scala 1492:74 lut_35.scala 1526:39]
  wire  _GEN_9973 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9627; // @[lut_35.scala 1492:74 lut_35.scala 1527:39]
  wire  _GEN_9974 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid | _GEN_9628; // @[lut_35.scala 1492:74 lut_35.scala 1528:34]
  wire  _GEN_9978 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1492:74 lut_35.scala 177:26 lut_35.scala 1530:27]
  wire  _GEN_9981 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9632; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_9984 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9635; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_9987 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9638; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_9990 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9641; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_9993 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9644; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_9996 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9647; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_9999 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9650; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10002 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9653; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10005 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9656; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10008 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9659; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10011 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9662; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10019 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9670; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10026 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9677; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10034 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9685; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10042 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9693; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10050 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9701; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10058 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9709; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10066 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9717; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10074 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9725; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10082 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9733; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10090 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9741; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10098 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9749; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10106 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9757; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10114 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9765; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10122 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9773; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10130 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9781; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10138 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9789; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10146 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9797; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10154 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9805; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10162 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9813; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10170 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9821; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10178 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9829; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10186 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9837; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10194 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9845; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10197 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9616; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10202 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9853; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10205 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9856; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10210 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9861; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10213 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9864; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10218 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9869; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10221 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9872; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10226 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9877; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10229 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9880; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10234 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9885; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10237 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9888; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10242 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9893; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10245 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9896; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10250 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9901; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10253 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9904; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10258 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9909; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10261 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9912; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10266 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9917; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10269 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9920; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10274 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9925; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10277 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9928; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10282 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9933; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10285 = LUT_mem_MPORT_198_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9936; // @[lut_35.scala 1492:74 lut_35.scala 177:26]
  wire  _GEN_10288 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9939; // @[lut_35.scala 1454:75 lut_35.scala 1455:38]
  wire  _GEN_10289 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9940; // @[lut_35.scala 1454:75 lut_35.scala 1456:38]
  wire  _GEN_10290 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9941; // @[lut_35.scala 1454:75 lut_35.scala 1457:38]
  wire  _GEN_10291 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9942; // @[lut_35.scala 1454:75 lut_35.scala 1458:38]
  wire  _GEN_10292 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9943; // @[lut_35.scala 1454:75 lut_35.scala 1459:38]
  wire  _GEN_10293 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9944; // @[lut_35.scala 1454:75 lut_35.scala 1460:38]
  wire  _GEN_10294 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9945; // @[lut_35.scala 1454:75 lut_35.scala 1461:38]
  wire  _GEN_10295 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9946; // @[lut_35.scala 1454:75 lut_35.scala 1462:38]
  wire  _GEN_10296 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9947; // @[lut_35.scala 1454:75 lut_35.scala 1463:38]
  wire  _GEN_10297 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9948; // @[lut_35.scala 1454:75 lut_35.scala 1464:38]
  wire  _GEN_10298 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9949; // @[lut_35.scala 1454:75 lut_35.scala 1465:39]
  wire  _GEN_10299 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9950; // @[lut_35.scala 1454:75 lut_35.scala 1466:39]
  wire  _GEN_10300 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9951; // @[lut_35.scala 1454:75 lut_35.scala 1467:39]
  wire  _GEN_10301 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9952; // @[lut_35.scala 1454:75 lut_35.scala 1468:39]
  wire  _GEN_10302 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9953; // @[lut_35.scala 1454:75 lut_35.scala 1469:39]
  wire  _GEN_10303 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9954; // @[lut_35.scala 1454:75 lut_35.scala 1470:39]
  wire  _GEN_10304 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9955; // @[lut_35.scala 1454:75 lut_35.scala 1471:39]
  wire  _GEN_10305 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9956; // @[lut_35.scala 1454:75 lut_35.scala 1472:39]
  wire  _GEN_10306 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9957; // @[lut_35.scala 1454:75 lut_35.scala 1473:39]
  wire  _GEN_10307 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9958; // @[lut_35.scala 1454:75 lut_35.scala 1474:39]
  wire  _GEN_10308 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9959; // @[lut_35.scala 1454:75 lut_35.scala 1475:39]
  wire  _GEN_10309 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9960; // @[lut_35.scala 1454:75 lut_35.scala 1476:39]
  wire  _GEN_10310 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid | _GEN_9961; // @[lut_35.scala 1454:75 lut_35.scala 1477:39]
  wire  _GEN_10311 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9962; // @[lut_35.scala 1454:75 lut_35.scala 1478:39]
  wire  _GEN_10312 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9963; // @[lut_35.scala 1454:75 lut_35.scala 1479:39]
  wire  _GEN_10313 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9964; // @[lut_35.scala 1454:75 lut_35.scala 1480:39]
  wire  _GEN_10314 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9965; // @[lut_35.scala 1454:75 lut_35.scala 1481:39]
  wire  _GEN_10315 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9966; // @[lut_35.scala 1454:75 lut_35.scala 1482:39]
  wire  _GEN_10316 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9967; // @[lut_35.scala 1454:75 lut_35.scala 1483:39]
  wire  _GEN_10317 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9968; // @[lut_35.scala 1454:75 lut_35.scala 1484:39]
  wire  _GEN_10318 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9969; // @[lut_35.scala 1454:75 lut_35.scala 1485:39]
  wire  _GEN_10319 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9970; // @[lut_35.scala 1454:75 lut_35.scala 1486:39]
  wire  _GEN_10320 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9971; // @[lut_35.scala 1454:75 lut_35.scala 1487:39]
  wire  _GEN_10321 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9972; // @[lut_35.scala 1454:75 lut_35.scala 1488:39]
  wire  _GEN_10322 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9973; // @[lut_35.scala 1454:75 lut_35.scala 1489:39]
  wire  _GEN_10323 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid | _GEN_9974; // @[lut_35.scala 1454:75 lut_35.scala 1490:34]
  wire  _GEN_10327 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1454:75 lut_35.scala 177:26 lut_35.scala 1492:27]
  wire  _GEN_10330 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9978; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10333 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9981; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10336 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9984; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10339 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9987; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10342 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9990; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10345 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9993; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10348 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9996; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10351 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9999; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10354 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10002; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10357 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10005; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10360 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10008; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10363 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10011; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10371 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10019; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10378 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10026; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10386 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10034; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10394 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10042; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10402 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10050; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10410 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10058; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10418 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10066; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10426 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10074; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10434 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10082; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10442 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10090; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10450 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10098; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10458 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10106; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10466 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10114; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10474 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10122; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10482 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10130; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10490 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10138; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10498 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10146; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10506 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10154; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10514 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10162; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10522 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10170; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10530 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10178; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10538 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10186; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10541 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_9961; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10546 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10194; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10549 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10197; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10554 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10202; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10557 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10205; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10562 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10210; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10565 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10213; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10570 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10218; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10573 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10221; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10578 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10226; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10581 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10229; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10586 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10234; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10589 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10237; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10594 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10242; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10597 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10245; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10602 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10250; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10605 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10253; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10610 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10258; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10613 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10261; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10618 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10266; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10621 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10269; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10626 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10274; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10629 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10277; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10634 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10282; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10637 = LUT_mem_MPORT_197_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10285; // @[lut_35.scala 1454:75 lut_35.scala 177:26]
  wire  _GEN_10640 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10288; // @[lut_35.scala 1416:74 lut_35.scala 1417:38]
  wire  _GEN_10641 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10289; // @[lut_35.scala 1416:74 lut_35.scala 1418:38]
  wire  _GEN_10642 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10290; // @[lut_35.scala 1416:74 lut_35.scala 1419:38]
  wire  _GEN_10643 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10291; // @[lut_35.scala 1416:74 lut_35.scala 1420:38]
  wire  _GEN_10644 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10292; // @[lut_35.scala 1416:74 lut_35.scala 1421:38]
  wire  _GEN_10645 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10293; // @[lut_35.scala 1416:74 lut_35.scala 1422:38]
  wire  _GEN_10646 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10294; // @[lut_35.scala 1416:74 lut_35.scala 1423:38]
  wire  _GEN_10647 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10295; // @[lut_35.scala 1416:74 lut_35.scala 1424:38]
  wire  _GEN_10648 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10296; // @[lut_35.scala 1416:74 lut_35.scala 1425:38]
  wire  _GEN_10649 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10297; // @[lut_35.scala 1416:74 lut_35.scala 1426:38]
  wire  _GEN_10650 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10298; // @[lut_35.scala 1416:74 lut_35.scala 1427:39]
  wire  _GEN_10651 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10299; // @[lut_35.scala 1416:74 lut_35.scala 1428:39]
  wire  _GEN_10652 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10300; // @[lut_35.scala 1416:74 lut_35.scala 1429:39]
  wire  _GEN_10653 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10301; // @[lut_35.scala 1416:74 lut_35.scala 1430:39]
  wire  _GEN_10654 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10302; // @[lut_35.scala 1416:74 lut_35.scala 1431:39]
  wire  _GEN_10655 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10303; // @[lut_35.scala 1416:74 lut_35.scala 1432:39]
  wire  _GEN_10656 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10304; // @[lut_35.scala 1416:74 lut_35.scala 1433:39]
  wire  _GEN_10657 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10305; // @[lut_35.scala 1416:74 lut_35.scala 1434:39]
  wire  _GEN_10658 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10306; // @[lut_35.scala 1416:74 lut_35.scala 1435:39]
  wire  _GEN_10659 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10307; // @[lut_35.scala 1416:74 lut_35.scala 1436:39]
  wire  _GEN_10660 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10308; // @[lut_35.scala 1416:74 lut_35.scala 1437:39]
  wire  _GEN_10661 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid | _GEN_10309; // @[lut_35.scala 1416:74 lut_35.scala 1438:39]
  wire  _GEN_10662 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10310; // @[lut_35.scala 1416:74 lut_35.scala 1439:39]
  wire  _GEN_10663 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10311; // @[lut_35.scala 1416:74 lut_35.scala 1440:39]
  wire  _GEN_10664 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10312; // @[lut_35.scala 1416:74 lut_35.scala 1441:39]
  wire  _GEN_10665 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10313; // @[lut_35.scala 1416:74 lut_35.scala 1442:39]
  wire  _GEN_10666 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10314; // @[lut_35.scala 1416:74 lut_35.scala 1443:39]
  wire  _GEN_10667 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10315; // @[lut_35.scala 1416:74 lut_35.scala 1444:39]
  wire  _GEN_10668 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10316; // @[lut_35.scala 1416:74 lut_35.scala 1445:39]
  wire  _GEN_10669 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10317; // @[lut_35.scala 1416:74 lut_35.scala 1446:39]
  wire  _GEN_10670 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10318; // @[lut_35.scala 1416:74 lut_35.scala 1447:39]
  wire  _GEN_10671 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10319; // @[lut_35.scala 1416:74 lut_35.scala 1448:39]
  wire  _GEN_10672 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10320; // @[lut_35.scala 1416:74 lut_35.scala 1449:39]
  wire  _GEN_10673 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10321; // @[lut_35.scala 1416:74 lut_35.scala 1450:39]
  wire  _GEN_10674 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10322; // @[lut_35.scala 1416:74 lut_35.scala 1451:39]
  wire  _GEN_10675 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid | _GEN_10323; // @[lut_35.scala 1416:74 lut_35.scala 1452:34]
  wire  _GEN_10679 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1416:74 lut_35.scala 177:26 lut_35.scala 1454:28]
  wire  _GEN_10682 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10327; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10685 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10330; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10688 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10333; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10691 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10336; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10694 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10339; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10697 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10342; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10700 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10345; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10703 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10348; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10706 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10351; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10709 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10354; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10712 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10357; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10715 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10360; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10718 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10363; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10726 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10371; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10733 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10378; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10741 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10386; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10749 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10394; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10757 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10402; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10765 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10410; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10773 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10418; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10781 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10426; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10789 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10434; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10797 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10442; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10805 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10450; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10813 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10458; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10821 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10466; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10829 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10474; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10837 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10482; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10845 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10490; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10853 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10498; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10861 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10506; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10869 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10514; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10877 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10522; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10885 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10530; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10888 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10309; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10893 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10538; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10896 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10541; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10901 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10546; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10904 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10549; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10909 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10554; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10912 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10557; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10917 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10562; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10920 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10565; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10925 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10570; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10928 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10573; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10933 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10578; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10936 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10581; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10941 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10586; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10944 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10589; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10949 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10594; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10952 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10597; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10957 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10602; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10960 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10605; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10965 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10610; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10968 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10613; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10973 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10618; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10976 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10621; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10981 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10626; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10984 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10629; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10989 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10634; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10992 = LUT_mem_MPORT_196_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10637; // @[lut_35.scala 1416:74 lut_35.scala 177:26]
  wire  _GEN_10995 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10640; // @[lut_35.scala 1378:74 lut_35.scala 1379:38]
  wire  _GEN_10996 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10641; // @[lut_35.scala 1378:74 lut_35.scala 1380:38]
  wire  _GEN_10997 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10642; // @[lut_35.scala 1378:74 lut_35.scala 1381:38]
  wire  _GEN_10998 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10643; // @[lut_35.scala 1378:74 lut_35.scala 1382:38]
  wire  _GEN_10999 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10644; // @[lut_35.scala 1378:74 lut_35.scala 1383:38]
  wire  _GEN_11000 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10645; // @[lut_35.scala 1378:74 lut_35.scala 1384:38]
  wire  _GEN_11001 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10646; // @[lut_35.scala 1378:74 lut_35.scala 1385:38]
  wire  _GEN_11002 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10647; // @[lut_35.scala 1378:74 lut_35.scala 1386:38]
  wire  _GEN_11003 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10648; // @[lut_35.scala 1378:74 lut_35.scala 1387:38]
  wire  _GEN_11004 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10649; // @[lut_35.scala 1378:74 lut_35.scala 1388:38]
  wire  _GEN_11005 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10650; // @[lut_35.scala 1378:74 lut_35.scala 1389:39]
  wire  _GEN_11006 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10651; // @[lut_35.scala 1378:74 lut_35.scala 1390:39]
  wire  _GEN_11007 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10652; // @[lut_35.scala 1378:74 lut_35.scala 1391:39]
  wire  _GEN_11008 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10653; // @[lut_35.scala 1378:74 lut_35.scala 1392:39]
  wire  _GEN_11009 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10654; // @[lut_35.scala 1378:74 lut_35.scala 1393:39]
  wire  _GEN_11010 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10655; // @[lut_35.scala 1378:74 lut_35.scala 1394:39]
  wire  _GEN_11011 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10656; // @[lut_35.scala 1378:74 lut_35.scala 1395:39]
  wire  _GEN_11012 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10657; // @[lut_35.scala 1378:74 lut_35.scala 1396:39]
  wire  _GEN_11013 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10658; // @[lut_35.scala 1378:74 lut_35.scala 1397:39]
  wire  _GEN_11014 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10659; // @[lut_35.scala 1378:74 lut_35.scala 1398:39]
  wire  _GEN_11015 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid | _GEN_10660; // @[lut_35.scala 1378:74 lut_35.scala 1399:39]
  wire  _GEN_11016 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10661; // @[lut_35.scala 1378:74 lut_35.scala 1400:39]
  wire  _GEN_11017 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10662; // @[lut_35.scala 1378:74 lut_35.scala 1401:39]
  wire  _GEN_11018 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10663; // @[lut_35.scala 1378:74 lut_35.scala 1402:39]
  wire  _GEN_11019 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10664; // @[lut_35.scala 1378:74 lut_35.scala 1403:39]
  wire  _GEN_11020 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10665; // @[lut_35.scala 1378:74 lut_35.scala 1404:39]
  wire  _GEN_11021 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10666; // @[lut_35.scala 1378:74 lut_35.scala 1405:39]
  wire  _GEN_11022 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10667; // @[lut_35.scala 1378:74 lut_35.scala 1406:39]
  wire  _GEN_11023 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10668; // @[lut_35.scala 1378:74 lut_35.scala 1407:39]
  wire  _GEN_11024 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10669; // @[lut_35.scala 1378:74 lut_35.scala 1408:39]
  wire  _GEN_11025 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10670; // @[lut_35.scala 1378:74 lut_35.scala 1409:39]
  wire  _GEN_11026 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10671; // @[lut_35.scala 1378:74 lut_35.scala 1410:39]
  wire  _GEN_11027 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10672; // @[lut_35.scala 1378:74 lut_35.scala 1411:39]
  wire  _GEN_11028 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10673; // @[lut_35.scala 1378:74 lut_35.scala 1412:39]
  wire  _GEN_11029 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10674; // @[lut_35.scala 1378:74 lut_35.scala 1413:39]
  wire  _GEN_11030 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid | _GEN_10675; // @[lut_35.scala 1378:74 lut_35.scala 1414:34]
  wire  _GEN_11034 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1378:74 lut_35.scala 177:26 lut_35.scala 1416:27]
  wire  _GEN_11037 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10679; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11040 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10682; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11043 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10685; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11046 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10688; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11049 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10691; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11052 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10694; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11055 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10697; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11058 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10700; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11061 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10703; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11064 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10706; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11067 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10709; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11070 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10712; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11073 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10715; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11076 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10718; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11084 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10726; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11091 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10733; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11099 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10741; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11107 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10749; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11115 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10757; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11123 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10765; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11131 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10773; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11139 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10781; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11147 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10789; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11155 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10797; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11163 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10805; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11171 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10813; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11179 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10821; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11187 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10829; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11195 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10837; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11203 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10845; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11211 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10853; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11219 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10861; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11227 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10869; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11235 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10877; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11238 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10660; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11243 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10885; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11246 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10888; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11251 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10893; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11254 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10896; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11259 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10901; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11262 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10904; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11267 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10909; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11270 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10912; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11275 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10917; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11278 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10920; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11283 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10925; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11286 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10928; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11291 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10933; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11294 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10936; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11299 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10941; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11302 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10944; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11307 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10949; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11310 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10952; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11315 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10957; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11318 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10960; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11323 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10965; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11326 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10968; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11331 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10973; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11334 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10976; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11339 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10981; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11342 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10984; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11347 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10989; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11350 = LUT_mem_MPORT_195_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10992; // @[lut_35.scala 1378:74 lut_35.scala 177:26]
  wire  _GEN_11353 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10995; // @[lut_35.scala 1340:74 lut_35.scala 1341:38]
  wire  _GEN_11354 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10996; // @[lut_35.scala 1340:74 lut_35.scala 1342:38]
  wire  _GEN_11355 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10997; // @[lut_35.scala 1340:74 lut_35.scala 1343:38]
  wire  _GEN_11356 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10998; // @[lut_35.scala 1340:74 lut_35.scala 1344:38]
  wire  _GEN_11357 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_10999; // @[lut_35.scala 1340:74 lut_35.scala 1345:38]
  wire  _GEN_11358 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11000; // @[lut_35.scala 1340:74 lut_35.scala 1346:38]
  wire  _GEN_11359 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11001; // @[lut_35.scala 1340:74 lut_35.scala 1347:38]
  wire  _GEN_11360 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11002; // @[lut_35.scala 1340:74 lut_35.scala 1348:38]
  wire  _GEN_11361 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11003; // @[lut_35.scala 1340:74 lut_35.scala 1349:38]
  wire  _GEN_11362 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11004; // @[lut_35.scala 1340:74 lut_35.scala 1350:38]
  wire  _GEN_11363 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11005; // @[lut_35.scala 1340:74 lut_35.scala 1351:39]
  wire  _GEN_11364 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11006; // @[lut_35.scala 1340:74 lut_35.scala 1352:39]
  wire  _GEN_11365 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11007; // @[lut_35.scala 1340:74 lut_35.scala 1353:39]
  wire  _GEN_11366 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11008; // @[lut_35.scala 1340:74 lut_35.scala 1354:39]
  wire  _GEN_11367 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11009; // @[lut_35.scala 1340:74 lut_35.scala 1355:39]
  wire  _GEN_11368 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11010; // @[lut_35.scala 1340:74 lut_35.scala 1356:39]
  wire  _GEN_11369 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11011; // @[lut_35.scala 1340:74 lut_35.scala 1357:39]
  wire  _GEN_11370 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11012; // @[lut_35.scala 1340:74 lut_35.scala 1358:39]
  wire  _GEN_11371 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11013; // @[lut_35.scala 1340:74 lut_35.scala 1359:39]
  wire  _GEN_11372 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid | _GEN_11014; // @[lut_35.scala 1340:74 lut_35.scala 1360:39]
  wire  _GEN_11373 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11015; // @[lut_35.scala 1340:74 lut_35.scala 1361:39]
  wire  _GEN_11374 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11016; // @[lut_35.scala 1340:74 lut_35.scala 1362:39]
  wire  _GEN_11375 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11017; // @[lut_35.scala 1340:74 lut_35.scala 1363:39]
  wire  _GEN_11376 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11018; // @[lut_35.scala 1340:74 lut_35.scala 1364:39]
  wire  _GEN_11377 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11019; // @[lut_35.scala 1340:74 lut_35.scala 1365:39]
  wire  _GEN_11378 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11020; // @[lut_35.scala 1340:74 lut_35.scala 1366:39]
  wire  _GEN_11379 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11021; // @[lut_35.scala 1340:74 lut_35.scala 1367:39]
  wire  _GEN_11380 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11022; // @[lut_35.scala 1340:74 lut_35.scala 1368:39]
  wire  _GEN_11381 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11023; // @[lut_35.scala 1340:74 lut_35.scala 1369:39]
  wire  _GEN_11382 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11024; // @[lut_35.scala 1340:74 lut_35.scala 1370:39]
  wire  _GEN_11383 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11025; // @[lut_35.scala 1340:74 lut_35.scala 1371:39]
  wire  _GEN_11384 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11026; // @[lut_35.scala 1340:74 lut_35.scala 1372:39]
  wire  _GEN_11385 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11027; // @[lut_35.scala 1340:74 lut_35.scala 1373:39]
  wire  _GEN_11386 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11028; // @[lut_35.scala 1340:74 lut_35.scala 1374:39]
  wire  _GEN_11387 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11029; // @[lut_35.scala 1340:74 lut_35.scala 1375:39]
  wire  _GEN_11388 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid | _GEN_11030; // @[lut_35.scala 1340:74 lut_35.scala 1376:34]
  wire  _GEN_11392 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1340:74 lut_35.scala 177:26 lut_35.scala 1378:27]
  wire  _GEN_11395 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11034; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11398 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11037; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11401 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11040; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11404 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11043; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11407 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11046; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11410 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11049; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11413 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11052; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11416 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11055; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11419 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11058; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11422 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11061; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11425 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11064; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11428 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11067; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11431 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11070; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11434 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11073; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11437 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11076; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11445 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11084; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11452 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11091; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11460 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11099; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11468 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11107; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11476 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11115; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11484 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11123; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11492 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11131; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11500 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11139; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11508 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11147; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11516 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11155; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11524 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11163; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11532 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11171; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11540 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11179; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11548 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11187; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11556 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11195; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11564 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11203; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11572 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11211; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11580 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11219; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11588 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11227; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11591 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11014; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11596 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11235; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11599 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11238; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11604 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11243; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11607 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11246; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11612 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11251; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11615 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11254; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11620 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11259; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11623 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11262; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11628 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11267; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11631 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11270; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11636 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11275; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11639 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11278; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11644 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11283; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11647 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11286; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11652 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11291; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11655 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11294; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11660 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11299; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11663 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11302; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11668 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11307; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11671 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11310; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11676 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11315; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11679 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11318; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11684 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11323; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11687 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11326; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11692 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11331; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11695 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11334; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11700 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11339; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11703 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11342; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11708 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11347; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11711 = LUT_mem_MPORT_194_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11350; // @[lut_35.scala 1340:74 lut_35.scala 177:26]
  wire  _GEN_11714 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11353; // @[lut_35.scala 1302:74 lut_35.scala 1303:38]
  wire  _GEN_11715 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11354; // @[lut_35.scala 1302:74 lut_35.scala 1304:38]
  wire  _GEN_11716 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11355; // @[lut_35.scala 1302:74 lut_35.scala 1305:38]
  wire  _GEN_11717 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11356; // @[lut_35.scala 1302:74 lut_35.scala 1306:38]
  wire  _GEN_11718 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11357; // @[lut_35.scala 1302:74 lut_35.scala 1307:38]
  wire  _GEN_11719 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11358; // @[lut_35.scala 1302:74 lut_35.scala 1308:38]
  wire  _GEN_11720 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11359; // @[lut_35.scala 1302:74 lut_35.scala 1309:38]
  wire  _GEN_11721 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11360; // @[lut_35.scala 1302:74 lut_35.scala 1310:38]
  wire  _GEN_11722 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11361; // @[lut_35.scala 1302:74 lut_35.scala 1311:38]
  wire  _GEN_11723 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11362; // @[lut_35.scala 1302:74 lut_35.scala 1312:38]
  wire  _GEN_11724 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11363; // @[lut_35.scala 1302:74 lut_35.scala 1313:39]
  wire  _GEN_11725 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11364; // @[lut_35.scala 1302:74 lut_35.scala 1314:39]
  wire  _GEN_11726 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11365; // @[lut_35.scala 1302:74 lut_35.scala 1315:39]
  wire  _GEN_11727 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11366; // @[lut_35.scala 1302:74 lut_35.scala 1316:39]
  wire  _GEN_11728 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11367; // @[lut_35.scala 1302:74 lut_35.scala 1317:39]
  wire  _GEN_11729 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11368; // @[lut_35.scala 1302:74 lut_35.scala 1318:39]
  wire  _GEN_11730 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11369; // @[lut_35.scala 1302:74 lut_35.scala 1319:39]
  wire  _GEN_11731 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11370; // @[lut_35.scala 1302:74 lut_35.scala 1320:39]
  wire  _GEN_11732 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid | _GEN_11371; // @[lut_35.scala 1302:74 lut_35.scala 1321:39]
  wire  _GEN_11733 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11372; // @[lut_35.scala 1302:74 lut_35.scala 1322:39]
  wire  _GEN_11734 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11373; // @[lut_35.scala 1302:74 lut_35.scala 1323:39]
  wire  _GEN_11735 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11374; // @[lut_35.scala 1302:74 lut_35.scala 1324:39]
  wire  _GEN_11736 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11375; // @[lut_35.scala 1302:74 lut_35.scala 1325:39]
  wire  _GEN_11737 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11376; // @[lut_35.scala 1302:74 lut_35.scala 1326:39]
  wire  _GEN_11738 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11377; // @[lut_35.scala 1302:74 lut_35.scala 1327:39]
  wire  _GEN_11739 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11378; // @[lut_35.scala 1302:74 lut_35.scala 1328:39]
  wire  _GEN_11740 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11379; // @[lut_35.scala 1302:74 lut_35.scala 1329:39]
  wire  _GEN_11741 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11380; // @[lut_35.scala 1302:74 lut_35.scala 1330:39]
  wire  _GEN_11742 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11381; // @[lut_35.scala 1302:74 lut_35.scala 1331:39]
  wire  _GEN_11743 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11382; // @[lut_35.scala 1302:74 lut_35.scala 1332:39]
  wire  _GEN_11744 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11383; // @[lut_35.scala 1302:74 lut_35.scala 1333:39]
  wire  _GEN_11745 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11384; // @[lut_35.scala 1302:74 lut_35.scala 1334:39]
  wire  _GEN_11746 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11385; // @[lut_35.scala 1302:74 lut_35.scala 1335:39]
  wire  _GEN_11747 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11386; // @[lut_35.scala 1302:74 lut_35.scala 1336:39]
  wire  _GEN_11748 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11387; // @[lut_35.scala 1302:74 lut_35.scala 1337:39]
  wire  _GEN_11749 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid | _GEN_11388; // @[lut_35.scala 1302:74 lut_35.scala 1338:34]
  wire  _GEN_11753 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1302:74 lut_35.scala 177:26 lut_35.scala 1340:27]
  wire  _GEN_11756 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11392; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11759 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11395; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11762 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11398; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11765 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11401; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11768 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11404; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11771 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11407; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11774 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11410; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11777 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11413; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11780 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11416; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11783 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11419; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11786 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11422; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11789 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11425; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11792 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11428; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11795 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11431; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11798 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11434; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11801 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11437; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11809 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11445; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11816 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11452; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11824 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11460; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11832 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11468; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11840 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11476; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11848 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11484; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11856 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11492; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11864 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11500; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11872 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11508; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11880 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11516; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11888 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11524; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11896 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11532; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11904 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11540; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11912 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11548; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11920 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11556; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11928 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11564; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11936 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11572; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11944 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11580; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11947 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11371; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11952 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11588; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11955 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11591; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11960 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11596; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11963 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11599; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11968 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11604; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11971 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11607; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11976 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11612; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11979 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11615; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11984 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11620; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11987 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11623; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11992 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11628; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_11995 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11631; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_12000 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11636; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_12003 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11639; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_12008 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11644; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_12011 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11647; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_12016 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11652; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_12019 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11655; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_12024 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11660; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_12027 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11663; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_12032 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11668; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_12035 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11671; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_12040 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11676; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_12043 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11679; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_12048 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11684; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_12051 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11687; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_12056 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11692; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_12059 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11695; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_12064 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11700; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_12067 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11703; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_12072 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11708; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_12075 = LUT_mem_MPORT_193_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11711; // @[lut_35.scala 1302:74 lut_35.scala 177:26]
  wire  _GEN_12078 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11714; // @[lut_35.scala 1264:74 lut_35.scala 1265:38]
  wire  _GEN_12079 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11715; // @[lut_35.scala 1264:74 lut_35.scala 1266:38]
  wire  _GEN_12080 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11716; // @[lut_35.scala 1264:74 lut_35.scala 1267:38]
  wire  _GEN_12081 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11717; // @[lut_35.scala 1264:74 lut_35.scala 1268:38]
  wire  _GEN_12082 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11718; // @[lut_35.scala 1264:74 lut_35.scala 1269:38]
  wire  _GEN_12083 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11719; // @[lut_35.scala 1264:74 lut_35.scala 1270:38]
  wire  _GEN_12084 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11720; // @[lut_35.scala 1264:74 lut_35.scala 1271:38]
  wire  _GEN_12085 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11721; // @[lut_35.scala 1264:74 lut_35.scala 1272:38]
  wire  _GEN_12086 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11722; // @[lut_35.scala 1264:74 lut_35.scala 1273:38]
  wire  _GEN_12087 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11723; // @[lut_35.scala 1264:74 lut_35.scala 1274:38]
  wire  _GEN_12088 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11724; // @[lut_35.scala 1264:74 lut_35.scala 1275:39]
  wire  _GEN_12089 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11725; // @[lut_35.scala 1264:74 lut_35.scala 1276:39]
  wire  _GEN_12090 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11726; // @[lut_35.scala 1264:74 lut_35.scala 1277:39]
  wire  _GEN_12091 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11727; // @[lut_35.scala 1264:74 lut_35.scala 1278:39]
  wire  _GEN_12092 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11728; // @[lut_35.scala 1264:74 lut_35.scala 1279:39]
  wire  _GEN_12093 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11729; // @[lut_35.scala 1264:74 lut_35.scala 1280:39]
  wire  _GEN_12094 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11730; // @[lut_35.scala 1264:74 lut_35.scala 1281:39]
  wire  _GEN_12095 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid | _GEN_11731; // @[lut_35.scala 1264:74 lut_35.scala 1282:39]
  wire  _GEN_12096 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11732; // @[lut_35.scala 1264:74 lut_35.scala 1283:39]
  wire  _GEN_12097 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11733; // @[lut_35.scala 1264:74 lut_35.scala 1284:39]
  wire  _GEN_12098 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11734; // @[lut_35.scala 1264:74 lut_35.scala 1285:39]
  wire  _GEN_12099 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11735; // @[lut_35.scala 1264:74 lut_35.scala 1286:39]
  wire  _GEN_12100 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11736; // @[lut_35.scala 1264:74 lut_35.scala 1287:39]
  wire  _GEN_12101 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11737; // @[lut_35.scala 1264:74 lut_35.scala 1288:39]
  wire  _GEN_12102 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11738; // @[lut_35.scala 1264:74 lut_35.scala 1289:39]
  wire  _GEN_12103 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11739; // @[lut_35.scala 1264:74 lut_35.scala 1290:39]
  wire  _GEN_12104 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11740; // @[lut_35.scala 1264:74 lut_35.scala 1291:39]
  wire  _GEN_12105 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11741; // @[lut_35.scala 1264:74 lut_35.scala 1292:39]
  wire  _GEN_12106 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11742; // @[lut_35.scala 1264:74 lut_35.scala 1293:39]
  wire  _GEN_12107 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11743; // @[lut_35.scala 1264:74 lut_35.scala 1294:39]
  wire  _GEN_12108 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11744; // @[lut_35.scala 1264:74 lut_35.scala 1295:39]
  wire  _GEN_12109 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11745; // @[lut_35.scala 1264:74 lut_35.scala 1296:39]
  wire  _GEN_12110 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11746; // @[lut_35.scala 1264:74 lut_35.scala 1297:39]
  wire  _GEN_12111 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11747; // @[lut_35.scala 1264:74 lut_35.scala 1298:39]
  wire  _GEN_12112 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11748; // @[lut_35.scala 1264:74 lut_35.scala 1299:39]
  wire  _GEN_12113 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid | _GEN_11749; // @[lut_35.scala 1264:74 lut_35.scala 1300:34]
  wire  _GEN_12117 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1264:74 lut_35.scala 177:26 lut_35.scala 1302:27]
  wire  _GEN_12120 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11753; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12123 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11756; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12126 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11759; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12129 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11762; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12132 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11765; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12135 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11768; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12138 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11771; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12141 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11774; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12144 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11777; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12147 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11780; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12150 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11783; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12153 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11786; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12156 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11789; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12159 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11792; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12162 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11795; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12165 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11798; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12168 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11801; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12176 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11809; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12183 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11816; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12191 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11824; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12199 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11832; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12207 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11840; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12215 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11848; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12223 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11856; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12231 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11864; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12239 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11872; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12247 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11880; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12255 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11888; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12263 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11896; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12271 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11904; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12279 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11912; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12287 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11920; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12295 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11928; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12303 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11936; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12306 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11731; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12311 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11944; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12314 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11947; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12319 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11952; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12322 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11955; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12327 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11960; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12330 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11963; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12335 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11968; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12338 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11971; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12343 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11976; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12346 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11979; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12351 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11984; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12354 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11987; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12359 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11992; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12362 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_11995; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12367 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12000; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12370 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12003; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12375 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12008; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12378 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12011; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12383 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12016; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12386 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12019; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12391 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12024; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12394 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12027; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12399 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12032; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12402 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12035; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12407 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12040; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12410 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12043; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12415 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12048; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12418 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12051; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12423 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12056; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12426 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12059; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12431 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12064; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12434 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12067; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12439 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12072; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12442 = LUT_mem_MPORT_192_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12075; // @[lut_35.scala 1264:74 lut_35.scala 177:26]
  wire  _GEN_12445 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12078; // @[lut_35.scala 1226:74 lut_35.scala 1227:38]
  wire  _GEN_12446 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12079; // @[lut_35.scala 1226:74 lut_35.scala 1228:38]
  wire  _GEN_12447 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12080; // @[lut_35.scala 1226:74 lut_35.scala 1229:38]
  wire  _GEN_12448 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12081; // @[lut_35.scala 1226:74 lut_35.scala 1230:38]
  wire  _GEN_12449 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12082; // @[lut_35.scala 1226:74 lut_35.scala 1231:38]
  wire  _GEN_12450 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12083; // @[lut_35.scala 1226:74 lut_35.scala 1232:38]
  wire  _GEN_12451 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12084; // @[lut_35.scala 1226:74 lut_35.scala 1233:38]
  wire  _GEN_12452 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12085; // @[lut_35.scala 1226:74 lut_35.scala 1234:38]
  wire  _GEN_12453 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12086; // @[lut_35.scala 1226:74 lut_35.scala 1235:38]
  wire  _GEN_12454 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12087; // @[lut_35.scala 1226:74 lut_35.scala 1236:38]
  wire  _GEN_12455 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12088; // @[lut_35.scala 1226:74 lut_35.scala 1237:39]
  wire  _GEN_12456 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12089; // @[lut_35.scala 1226:74 lut_35.scala 1238:39]
  wire  _GEN_12457 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12090; // @[lut_35.scala 1226:74 lut_35.scala 1239:39]
  wire  _GEN_12458 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12091; // @[lut_35.scala 1226:74 lut_35.scala 1240:39]
  wire  _GEN_12459 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12092; // @[lut_35.scala 1226:74 lut_35.scala 1241:39]
  wire  _GEN_12460 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12093; // @[lut_35.scala 1226:74 lut_35.scala 1242:39]
  wire  _GEN_12461 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid | _GEN_12094; // @[lut_35.scala 1226:74 lut_35.scala 1243:39]
  wire  _GEN_12462 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12095; // @[lut_35.scala 1226:74 lut_35.scala 1244:39]
  wire  _GEN_12463 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12096; // @[lut_35.scala 1226:74 lut_35.scala 1245:39]
  wire  _GEN_12464 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12097; // @[lut_35.scala 1226:74 lut_35.scala 1246:39]
  wire  _GEN_12465 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12098; // @[lut_35.scala 1226:74 lut_35.scala 1247:39]
  wire  _GEN_12466 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12099; // @[lut_35.scala 1226:74 lut_35.scala 1248:39]
  wire  _GEN_12467 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12100; // @[lut_35.scala 1226:74 lut_35.scala 1249:39]
  wire  _GEN_12468 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12101; // @[lut_35.scala 1226:74 lut_35.scala 1250:39]
  wire  _GEN_12469 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12102; // @[lut_35.scala 1226:74 lut_35.scala 1251:39]
  wire  _GEN_12470 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12103; // @[lut_35.scala 1226:74 lut_35.scala 1252:39]
  wire  _GEN_12471 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12104; // @[lut_35.scala 1226:74 lut_35.scala 1253:39]
  wire  _GEN_12472 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12105; // @[lut_35.scala 1226:74 lut_35.scala 1254:39]
  wire  _GEN_12473 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12106; // @[lut_35.scala 1226:74 lut_35.scala 1255:39]
  wire  _GEN_12474 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12107; // @[lut_35.scala 1226:74 lut_35.scala 1256:39]
  wire  _GEN_12475 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12108; // @[lut_35.scala 1226:74 lut_35.scala 1257:39]
  wire  _GEN_12476 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12109; // @[lut_35.scala 1226:74 lut_35.scala 1258:39]
  wire  _GEN_12477 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12110; // @[lut_35.scala 1226:74 lut_35.scala 1259:39]
  wire  _GEN_12478 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12111; // @[lut_35.scala 1226:74 lut_35.scala 1260:39]
  wire  _GEN_12479 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12112; // @[lut_35.scala 1226:74 lut_35.scala 1261:39]
  wire  _GEN_12480 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid | _GEN_12113; // @[lut_35.scala 1226:74 lut_35.scala 1262:34]
  wire  _GEN_12484 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1226:74 lut_35.scala 177:26 lut_35.scala 1264:27]
  wire  _GEN_12487 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12117; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12490 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12120; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12493 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12123; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12496 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12126; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12499 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12129; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12502 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12132; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12505 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12135; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12508 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12138; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12511 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12141; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12514 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12144; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12517 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12147; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12520 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12150; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12523 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12153; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12526 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12156; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12529 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12159; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12532 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12162; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12535 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12165; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12538 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12168; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12546 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12176; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12553 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12183; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12561 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12191; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12569 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12199; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12577 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12207; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12585 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12215; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12593 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12223; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12601 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12231; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12609 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12239; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12617 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12247; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12625 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12255; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12633 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12263; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12641 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12271; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12649 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12279; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12657 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12287; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12665 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12295; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12668 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12094; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12673 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12303; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12676 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12306; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12681 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12311; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12684 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12314; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12689 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12319; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12692 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12322; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12697 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12327; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12700 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12330; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12705 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12335; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12708 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12338; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12713 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12343; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12716 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12346; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12721 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12351; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12724 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12354; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12729 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12359; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12732 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12362; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12737 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12367; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12740 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12370; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12745 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12375; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12748 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12378; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12753 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12383; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12756 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12386; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12761 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12391; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12764 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12394; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12769 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12399; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12772 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12402; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12777 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12407; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12780 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12410; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12785 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12415; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12788 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12418; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12793 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12423; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12796 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12426; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12801 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12431; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12804 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12434; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12809 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12439; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12812 = LUT_mem_MPORT_191_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12442; // @[lut_35.scala 1226:74 lut_35.scala 177:26]
  wire  _GEN_12815 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12445; // @[lut_35.scala 1188:74 lut_35.scala 1189:38]
  wire  _GEN_12816 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12446; // @[lut_35.scala 1188:74 lut_35.scala 1190:38]
  wire  _GEN_12817 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12447; // @[lut_35.scala 1188:74 lut_35.scala 1191:38]
  wire  _GEN_12818 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12448; // @[lut_35.scala 1188:74 lut_35.scala 1192:38]
  wire  _GEN_12819 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12449; // @[lut_35.scala 1188:74 lut_35.scala 1193:38]
  wire  _GEN_12820 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12450; // @[lut_35.scala 1188:74 lut_35.scala 1194:38]
  wire  _GEN_12821 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12451; // @[lut_35.scala 1188:74 lut_35.scala 1195:38]
  wire  _GEN_12822 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12452; // @[lut_35.scala 1188:74 lut_35.scala 1196:38]
  wire  _GEN_12823 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12453; // @[lut_35.scala 1188:74 lut_35.scala 1197:38]
  wire  _GEN_12824 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12454; // @[lut_35.scala 1188:74 lut_35.scala 1198:38]
  wire  _GEN_12825 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12455; // @[lut_35.scala 1188:74 lut_35.scala 1199:39]
  wire  _GEN_12826 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12456; // @[lut_35.scala 1188:74 lut_35.scala 1200:39]
  wire  _GEN_12827 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12457; // @[lut_35.scala 1188:74 lut_35.scala 1201:39]
  wire  _GEN_12828 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12458; // @[lut_35.scala 1188:74 lut_35.scala 1202:39]
  wire  _GEN_12829 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12459; // @[lut_35.scala 1188:74 lut_35.scala 1203:39]
  wire  _GEN_12830 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid | _GEN_12460; // @[lut_35.scala 1188:74 lut_35.scala 1204:39]
  wire  _GEN_12831 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12461; // @[lut_35.scala 1188:74 lut_35.scala 1205:39]
  wire  _GEN_12832 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12462; // @[lut_35.scala 1188:74 lut_35.scala 1206:39]
  wire  _GEN_12833 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12463; // @[lut_35.scala 1188:74 lut_35.scala 1207:39]
  wire  _GEN_12834 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12464; // @[lut_35.scala 1188:74 lut_35.scala 1208:39]
  wire  _GEN_12835 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12465; // @[lut_35.scala 1188:74 lut_35.scala 1209:39]
  wire  _GEN_12836 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12466; // @[lut_35.scala 1188:74 lut_35.scala 1210:39]
  wire  _GEN_12837 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12467; // @[lut_35.scala 1188:74 lut_35.scala 1211:39]
  wire  _GEN_12838 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12468; // @[lut_35.scala 1188:74 lut_35.scala 1212:39]
  wire  _GEN_12839 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12469; // @[lut_35.scala 1188:74 lut_35.scala 1213:39]
  wire  _GEN_12840 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12470; // @[lut_35.scala 1188:74 lut_35.scala 1214:39]
  wire  _GEN_12841 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12471; // @[lut_35.scala 1188:74 lut_35.scala 1215:39]
  wire  _GEN_12842 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12472; // @[lut_35.scala 1188:74 lut_35.scala 1216:39]
  wire  _GEN_12843 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12473; // @[lut_35.scala 1188:74 lut_35.scala 1217:39]
  wire  _GEN_12844 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12474; // @[lut_35.scala 1188:74 lut_35.scala 1218:39]
  wire  _GEN_12845 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12475; // @[lut_35.scala 1188:74 lut_35.scala 1219:39]
  wire  _GEN_12846 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12476; // @[lut_35.scala 1188:74 lut_35.scala 1220:39]
  wire  _GEN_12847 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12477; // @[lut_35.scala 1188:74 lut_35.scala 1221:39]
  wire  _GEN_12848 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12478; // @[lut_35.scala 1188:74 lut_35.scala 1222:39]
  wire  _GEN_12849 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12479; // @[lut_35.scala 1188:74 lut_35.scala 1223:39]
  wire  _GEN_12850 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid | _GEN_12480; // @[lut_35.scala 1188:74 lut_35.scala 1224:34]
  wire  _GEN_12854 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1188:74 lut_35.scala 177:26 lut_35.scala 1226:27]
  wire  _GEN_12857 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12484; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_12860 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12487; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_12863 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12490; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_12866 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12493; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_12869 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12496; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_12872 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12499; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_12875 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12502; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_12878 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12505; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_12881 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12508; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_12884 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12511; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_12887 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12514; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_12890 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12517; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_12893 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12520; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_12896 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12523; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_12899 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12526; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_12902 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12529; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_12905 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12532; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_12908 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12535; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_12911 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12538; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_12919 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12546; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_12926 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12553; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_12934 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12561; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_12942 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12569; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_12950 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12577; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_12958 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12585; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_12966 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12593; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_12974 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12601; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_12982 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12609; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_12990 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12617; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_12998 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12625; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13006 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12633; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13014 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12641; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13022 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12649; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13030 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12657; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13033 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12460; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13038 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12665; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13041 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12668; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13046 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12673; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13049 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12676; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13054 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12681; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13057 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12684; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13062 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12689; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13065 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12692; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13070 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12697; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13073 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12700; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13078 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12705; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13081 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12708; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13086 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12713; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13089 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12716; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13094 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12721; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13097 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12724; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13102 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12729; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13105 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12732; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13110 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12737; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13113 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12740; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13118 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12745; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13121 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12748; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13126 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12753; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13129 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12756; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13134 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12761; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13137 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12764; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13142 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12769; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13145 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12772; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13150 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12777; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13153 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12780; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13158 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12785; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13161 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12788; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13166 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12793; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13169 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12796; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13174 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12801; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13177 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12804; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13182 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12809; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13185 = LUT_mem_MPORT_190_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12812; // @[lut_35.scala 1188:74 lut_35.scala 177:26]
  wire  _GEN_13188 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12815; // @[lut_35.scala 1150:74 lut_35.scala 1151:38]
  wire  _GEN_13189 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12816; // @[lut_35.scala 1150:74 lut_35.scala 1152:38]
  wire  _GEN_13190 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12817; // @[lut_35.scala 1150:74 lut_35.scala 1153:38]
  wire  _GEN_13191 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12818; // @[lut_35.scala 1150:74 lut_35.scala 1154:38]
  wire  _GEN_13192 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12819; // @[lut_35.scala 1150:74 lut_35.scala 1155:38]
  wire  _GEN_13193 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12820; // @[lut_35.scala 1150:74 lut_35.scala 1156:38]
  wire  _GEN_13194 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12821; // @[lut_35.scala 1150:74 lut_35.scala 1157:38]
  wire  _GEN_13195 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12822; // @[lut_35.scala 1150:74 lut_35.scala 1158:38]
  wire  _GEN_13196 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12823; // @[lut_35.scala 1150:74 lut_35.scala 1159:38]
  wire  _GEN_13197 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12824; // @[lut_35.scala 1150:74 lut_35.scala 1160:38]
  wire  _GEN_13198 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12825; // @[lut_35.scala 1150:74 lut_35.scala 1161:39]
  wire  _GEN_13199 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12826; // @[lut_35.scala 1150:74 lut_35.scala 1162:39]
  wire  _GEN_13200 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12827; // @[lut_35.scala 1150:74 lut_35.scala 1163:39]
  wire  _GEN_13201 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12828; // @[lut_35.scala 1150:74 lut_35.scala 1164:39]
  wire  _GEN_13202 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid | _GEN_12829; // @[lut_35.scala 1150:74 lut_35.scala 1165:39]
  wire  _GEN_13203 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12830; // @[lut_35.scala 1150:74 lut_35.scala 1166:39]
  wire  _GEN_13204 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12831; // @[lut_35.scala 1150:74 lut_35.scala 1167:39]
  wire  _GEN_13205 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12832; // @[lut_35.scala 1150:74 lut_35.scala 1168:39]
  wire  _GEN_13206 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12833; // @[lut_35.scala 1150:74 lut_35.scala 1169:39]
  wire  _GEN_13207 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12834; // @[lut_35.scala 1150:74 lut_35.scala 1170:39]
  wire  _GEN_13208 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12835; // @[lut_35.scala 1150:74 lut_35.scala 1171:39]
  wire  _GEN_13209 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12836; // @[lut_35.scala 1150:74 lut_35.scala 1172:39]
  wire  _GEN_13210 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12837; // @[lut_35.scala 1150:74 lut_35.scala 1173:39]
  wire  _GEN_13211 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12838; // @[lut_35.scala 1150:74 lut_35.scala 1174:39]
  wire  _GEN_13212 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12839; // @[lut_35.scala 1150:74 lut_35.scala 1175:39]
  wire  _GEN_13213 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12840; // @[lut_35.scala 1150:74 lut_35.scala 1176:39]
  wire  _GEN_13214 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12841; // @[lut_35.scala 1150:74 lut_35.scala 1177:39]
  wire  _GEN_13215 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12842; // @[lut_35.scala 1150:74 lut_35.scala 1178:39]
  wire  _GEN_13216 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12843; // @[lut_35.scala 1150:74 lut_35.scala 1179:39]
  wire  _GEN_13217 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12844; // @[lut_35.scala 1150:74 lut_35.scala 1180:39]
  wire  _GEN_13218 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12845; // @[lut_35.scala 1150:74 lut_35.scala 1181:39]
  wire  _GEN_13219 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12846; // @[lut_35.scala 1150:74 lut_35.scala 1182:39]
  wire  _GEN_13220 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12847; // @[lut_35.scala 1150:74 lut_35.scala 1183:39]
  wire  _GEN_13221 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12848; // @[lut_35.scala 1150:74 lut_35.scala 1184:39]
  wire  _GEN_13222 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12849; // @[lut_35.scala 1150:74 lut_35.scala 1185:39]
  wire  _GEN_13223 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid | _GEN_12850; // @[lut_35.scala 1150:74 lut_35.scala 1186:34]
  wire  _GEN_13227 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1150:74 lut_35.scala 177:26 lut_35.scala 1188:27]
  wire  _GEN_13230 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12854; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13233 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12857; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13236 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12860; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13239 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12863; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13242 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12866; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13245 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12869; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13248 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12872; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13251 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12875; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13254 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12878; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13257 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12881; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13260 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12884; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13263 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12887; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13266 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12890; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13269 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12893; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13272 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12896; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13275 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12899; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13278 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12902; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13281 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12905; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13284 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12908; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13287 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12911; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13295 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12919; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13302 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12926; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13310 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12934; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13318 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12942; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13326 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12950; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13334 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12958; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13342 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12966; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13350 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12974; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13358 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12982; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13366 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12990; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13374 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12998; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13382 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13006; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13390 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13014; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13398 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13022; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13401 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_12829; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13406 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13030; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13409 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13033; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13414 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13038; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13417 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13041; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13422 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13046; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13425 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13049; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13430 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13054; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13433 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13057; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13438 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13062; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13441 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13065; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13446 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13070; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13449 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13073; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13454 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13078; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13457 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13081; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13462 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13086; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13465 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13089; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13470 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13094; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13473 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13097; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13478 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13102; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13481 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13105; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13486 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13110; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13489 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13113; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13494 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13118; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13497 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13121; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13502 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13126; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13505 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13129; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13510 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13134; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13513 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13137; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13518 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13142; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13521 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13145; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13526 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13150; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13529 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13153; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13534 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13158; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13537 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13161; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13542 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13166; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13545 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13169; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13550 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13174; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13553 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13177; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13558 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13182; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13561 = LUT_mem_MPORT_189_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13185; // @[lut_35.scala 1150:74 lut_35.scala 177:26]
  wire  _GEN_13564 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13188; // @[lut_35.scala 1112:74 lut_35.scala 1113:38]
  wire  _GEN_13565 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13189; // @[lut_35.scala 1112:74 lut_35.scala 1114:38]
  wire  _GEN_13566 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13190; // @[lut_35.scala 1112:74 lut_35.scala 1115:38]
  wire  _GEN_13567 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13191; // @[lut_35.scala 1112:74 lut_35.scala 1116:38]
  wire  _GEN_13568 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13192; // @[lut_35.scala 1112:74 lut_35.scala 1117:38]
  wire  _GEN_13569 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13193; // @[lut_35.scala 1112:74 lut_35.scala 1118:38]
  wire  _GEN_13570 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13194; // @[lut_35.scala 1112:74 lut_35.scala 1119:38]
  wire  _GEN_13571 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13195; // @[lut_35.scala 1112:74 lut_35.scala 1120:38]
  wire  _GEN_13572 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13196; // @[lut_35.scala 1112:74 lut_35.scala 1121:38]
  wire  _GEN_13573 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13197; // @[lut_35.scala 1112:74 lut_35.scala 1122:38]
  wire  _GEN_13574 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13198; // @[lut_35.scala 1112:74 lut_35.scala 1123:39]
  wire  _GEN_13575 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13199; // @[lut_35.scala 1112:74 lut_35.scala 1124:39]
  wire  _GEN_13576 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13200; // @[lut_35.scala 1112:74 lut_35.scala 1125:39]
  wire  _GEN_13577 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid | _GEN_13201; // @[lut_35.scala 1112:74 lut_35.scala 1126:39]
  wire  _GEN_13578 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13202; // @[lut_35.scala 1112:74 lut_35.scala 1127:39]
  wire  _GEN_13579 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13203; // @[lut_35.scala 1112:74 lut_35.scala 1128:39]
  wire  _GEN_13580 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13204; // @[lut_35.scala 1112:74 lut_35.scala 1129:39]
  wire  _GEN_13581 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13205; // @[lut_35.scala 1112:74 lut_35.scala 1130:39]
  wire  _GEN_13582 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13206; // @[lut_35.scala 1112:74 lut_35.scala 1131:39]
  wire  _GEN_13583 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13207; // @[lut_35.scala 1112:74 lut_35.scala 1132:39]
  wire  _GEN_13584 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13208; // @[lut_35.scala 1112:74 lut_35.scala 1133:39]
  wire  _GEN_13585 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13209; // @[lut_35.scala 1112:74 lut_35.scala 1134:39]
  wire  _GEN_13586 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13210; // @[lut_35.scala 1112:74 lut_35.scala 1135:39]
  wire  _GEN_13587 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13211; // @[lut_35.scala 1112:74 lut_35.scala 1136:39]
  wire  _GEN_13588 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13212; // @[lut_35.scala 1112:74 lut_35.scala 1137:39]
  wire  _GEN_13589 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13213; // @[lut_35.scala 1112:74 lut_35.scala 1138:39]
  wire  _GEN_13590 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13214; // @[lut_35.scala 1112:74 lut_35.scala 1139:39]
  wire  _GEN_13591 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13215; // @[lut_35.scala 1112:74 lut_35.scala 1140:39]
  wire  _GEN_13592 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13216; // @[lut_35.scala 1112:74 lut_35.scala 1141:39]
  wire  _GEN_13593 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13217; // @[lut_35.scala 1112:74 lut_35.scala 1142:39]
  wire  _GEN_13594 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13218; // @[lut_35.scala 1112:74 lut_35.scala 1143:39]
  wire  _GEN_13595 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13219; // @[lut_35.scala 1112:74 lut_35.scala 1144:39]
  wire  _GEN_13596 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13220; // @[lut_35.scala 1112:74 lut_35.scala 1145:39]
  wire  _GEN_13597 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13221; // @[lut_35.scala 1112:74 lut_35.scala 1146:39]
  wire  _GEN_13598 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13222; // @[lut_35.scala 1112:74 lut_35.scala 1147:39]
  wire  _GEN_13599 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid | _GEN_13223; // @[lut_35.scala 1112:74 lut_35.scala 1148:34]
  wire  _GEN_13603 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1112:74 lut_35.scala 177:26 lut_35.scala 1150:27]
  wire  _GEN_13606 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13227; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13609 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13230; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13612 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13233; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13615 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13236; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13618 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13239; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13621 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13242; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13624 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13245; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13627 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13248; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13630 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13251; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13633 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13254; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13636 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13257; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13639 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13260; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13642 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13263; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13645 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13266; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13648 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13269; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13651 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13272; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13654 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13275; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13657 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13278; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13660 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13281; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13663 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13284; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13666 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13287; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13674 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13295; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13681 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13302; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13689 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13310; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13697 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13318; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13705 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13326; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13713 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13334; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13721 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13342; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13729 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13350; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13737 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13358; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13745 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13366; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13753 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13374; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13761 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13382; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13769 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13390; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13772 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13201; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13777 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13398; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13780 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13401; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13785 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13406; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13788 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13409; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13793 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13414; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13796 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13417; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13801 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13422; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13804 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13425; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13809 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13430; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13812 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13433; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13817 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13438; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13820 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13441; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13825 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13446; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13828 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13449; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13833 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13454; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13836 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13457; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13841 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13462; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13844 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13465; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13849 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13470; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13852 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13473; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13857 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13478; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13860 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13481; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13865 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13486; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13868 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13489; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13873 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13494; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13876 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13497; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13881 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13502; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13884 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13505; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13889 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13510; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13892 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13513; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13897 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13518; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13900 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13521; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13905 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13526; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13908 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13529; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13913 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13534; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13916 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13537; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13921 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13542; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13924 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13545; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13929 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13550; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13932 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13553; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13937 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13558; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13940 = LUT_mem_MPORT_188_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13561; // @[lut_35.scala 1112:74 lut_35.scala 177:26]
  wire  _GEN_13943 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13564; // @[lut_35.scala 1074:74 lut_35.scala 1075:38]
  wire  _GEN_13944 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13565; // @[lut_35.scala 1074:74 lut_35.scala 1076:38]
  wire  _GEN_13945 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13566; // @[lut_35.scala 1074:74 lut_35.scala 1077:38]
  wire  _GEN_13946 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13567; // @[lut_35.scala 1074:74 lut_35.scala 1078:38]
  wire  _GEN_13947 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13568; // @[lut_35.scala 1074:74 lut_35.scala 1079:38]
  wire  _GEN_13948 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13569; // @[lut_35.scala 1074:74 lut_35.scala 1080:38]
  wire  _GEN_13949 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13570; // @[lut_35.scala 1074:74 lut_35.scala 1081:38]
  wire  _GEN_13950 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13571; // @[lut_35.scala 1074:74 lut_35.scala 1082:38]
  wire  _GEN_13951 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13572; // @[lut_35.scala 1074:74 lut_35.scala 1083:38]
  wire  _GEN_13952 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13573; // @[lut_35.scala 1074:74 lut_35.scala 1084:38]
  wire  _GEN_13953 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13574; // @[lut_35.scala 1074:74 lut_35.scala 1085:39]
  wire  _GEN_13954 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13575; // @[lut_35.scala 1074:74 lut_35.scala 1086:39]
  wire  _GEN_13955 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid | _GEN_13576; // @[lut_35.scala 1074:74 lut_35.scala 1087:39]
  wire  _GEN_13956 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13577; // @[lut_35.scala 1074:74 lut_35.scala 1088:39]
  wire  _GEN_13957 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13578; // @[lut_35.scala 1074:74 lut_35.scala 1089:39]
  wire  _GEN_13958 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13579; // @[lut_35.scala 1074:74 lut_35.scala 1090:39]
  wire  _GEN_13959 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13580; // @[lut_35.scala 1074:74 lut_35.scala 1091:39]
  wire  _GEN_13960 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13581; // @[lut_35.scala 1074:74 lut_35.scala 1092:39]
  wire  _GEN_13961 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13582; // @[lut_35.scala 1074:74 lut_35.scala 1093:39]
  wire  _GEN_13962 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13583; // @[lut_35.scala 1074:74 lut_35.scala 1094:39]
  wire  _GEN_13963 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13584; // @[lut_35.scala 1074:74 lut_35.scala 1095:39]
  wire  _GEN_13964 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13585; // @[lut_35.scala 1074:74 lut_35.scala 1096:39]
  wire  _GEN_13965 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13586; // @[lut_35.scala 1074:74 lut_35.scala 1097:39]
  wire  _GEN_13966 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13587; // @[lut_35.scala 1074:74 lut_35.scala 1098:39]
  wire  _GEN_13967 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13588; // @[lut_35.scala 1074:74 lut_35.scala 1099:39]
  wire  _GEN_13968 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13589; // @[lut_35.scala 1074:74 lut_35.scala 1100:39]
  wire  _GEN_13969 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13590; // @[lut_35.scala 1074:74 lut_35.scala 1101:39]
  wire  _GEN_13970 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13591; // @[lut_35.scala 1074:74 lut_35.scala 1102:39]
  wire  _GEN_13971 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13592; // @[lut_35.scala 1074:74 lut_35.scala 1103:39]
  wire  _GEN_13972 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13593; // @[lut_35.scala 1074:74 lut_35.scala 1104:39]
  wire  _GEN_13973 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13594; // @[lut_35.scala 1074:74 lut_35.scala 1105:39]
  wire  _GEN_13974 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13595; // @[lut_35.scala 1074:74 lut_35.scala 1106:39]
  wire  _GEN_13975 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13596; // @[lut_35.scala 1074:74 lut_35.scala 1107:39]
  wire  _GEN_13976 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13597; // @[lut_35.scala 1074:74 lut_35.scala 1108:39]
  wire  _GEN_13977 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13598; // @[lut_35.scala 1074:74 lut_35.scala 1109:39]
  wire  _GEN_13978 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid | _GEN_13599; // @[lut_35.scala 1074:74 lut_35.scala 1110:34]
  wire  _GEN_13982 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1074:74 lut_35.scala 177:26 lut_35.scala 1112:27]
  wire  _GEN_13985 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13603; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_13988 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13606; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_13991 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13609; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_13994 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13612; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_13997 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13615; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14000 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13618; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14003 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13621; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14006 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13624; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14009 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13627; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14012 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13630; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14015 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13633; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14018 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13636; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14021 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13639; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14024 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13642; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14027 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13645; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14030 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13648; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14033 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13651; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14036 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13654; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14039 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13657; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14042 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13660; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14045 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13663; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14048 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13666; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14056 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13674; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14063 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13681; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14071 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13689; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14079 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13697; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14087 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13705; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14095 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13713; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14103 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13721; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14111 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13729; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14119 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13737; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14127 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13745; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14135 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13753; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14143 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13761; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14146 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13576; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14151 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13769; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14154 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13772; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14159 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13777; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14162 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13780; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14167 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13785; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14170 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13788; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14175 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13793; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14178 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13796; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14183 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13801; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14186 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13804; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14191 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13809; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14194 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13812; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14199 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13817; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14202 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13820; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14207 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13825; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14210 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13828; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14215 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13833; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14218 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13836; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14223 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13841; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14226 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13844; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14231 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13849; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14234 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13852; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14239 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13857; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14242 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13860; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14247 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13865; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14250 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13868; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14255 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13873; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14258 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13876; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14263 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13881; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14266 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13884; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14271 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13889; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14274 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13892; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14279 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13897; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14282 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13900; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14287 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13905; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14290 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13908; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14295 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13913; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14298 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13916; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14303 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13921; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14306 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13924; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14311 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13929; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14314 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13932; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14319 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13937; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14322 = LUT_mem_MPORT_187_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13940; // @[lut_35.scala 1074:74 lut_35.scala 177:26]
  wire  _GEN_14325 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13943; // @[lut_35.scala 1036:74 lut_35.scala 1037:38]
  wire  _GEN_14326 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13944; // @[lut_35.scala 1036:74 lut_35.scala 1038:38]
  wire  _GEN_14327 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13945; // @[lut_35.scala 1036:74 lut_35.scala 1039:38]
  wire  _GEN_14328 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13946; // @[lut_35.scala 1036:74 lut_35.scala 1040:38]
  wire  _GEN_14329 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13947; // @[lut_35.scala 1036:74 lut_35.scala 1041:38]
  wire  _GEN_14330 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13948; // @[lut_35.scala 1036:74 lut_35.scala 1042:38]
  wire  _GEN_14331 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13949; // @[lut_35.scala 1036:74 lut_35.scala 1043:38]
  wire  _GEN_14332 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13950; // @[lut_35.scala 1036:74 lut_35.scala 1044:38]
  wire  _GEN_14333 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13951; // @[lut_35.scala 1036:74 lut_35.scala 1045:38]
  wire  _GEN_14334 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13952; // @[lut_35.scala 1036:74 lut_35.scala 1046:38]
  wire  _GEN_14335 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13953; // @[lut_35.scala 1036:74 lut_35.scala 1047:39]
  wire  _GEN_14336 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid | _GEN_13954; // @[lut_35.scala 1036:74 lut_35.scala 1048:39]
  wire  _GEN_14337 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13955; // @[lut_35.scala 1036:74 lut_35.scala 1049:39]
  wire  _GEN_14338 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13956; // @[lut_35.scala 1036:74 lut_35.scala 1050:39]
  wire  _GEN_14339 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13957; // @[lut_35.scala 1036:74 lut_35.scala 1051:39]
  wire  _GEN_14340 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13958; // @[lut_35.scala 1036:74 lut_35.scala 1052:39]
  wire  _GEN_14341 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13959; // @[lut_35.scala 1036:74 lut_35.scala 1053:39]
  wire  _GEN_14342 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13960; // @[lut_35.scala 1036:74 lut_35.scala 1054:39]
  wire  _GEN_14343 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13961; // @[lut_35.scala 1036:74 lut_35.scala 1055:39]
  wire  _GEN_14344 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13962; // @[lut_35.scala 1036:74 lut_35.scala 1056:39]
  wire  _GEN_14345 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13963; // @[lut_35.scala 1036:74 lut_35.scala 1057:39]
  wire  _GEN_14346 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13964; // @[lut_35.scala 1036:74 lut_35.scala 1058:39]
  wire  _GEN_14347 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13965; // @[lut_35.scala 1036:74 lut_35.scala 1059:39]
  wire  _GEN_14348 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13966; // @[lut_35.scala 1036:74 lut_35.scala 1060:39]
  wire  _GEN_14349 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13967; // @[lut_35.scala 1036:74 lut_35.scala 1061:39]
  wire  _GEN_14350 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13968; // @[lut_35.scala 1036:74 lut_35.scala 1062:39]
  wire  _GEN_14351 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13969; // @[lut_35.scala 1036:74 lut_35.scala 1063:39]
  wire  _GEN_14352 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13970; // @[lut_35.scala 1036:74 lut_35.scala 1064:39]
  wire  _GEN_14353 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13971; // @[lut_35.scala 1036:74 lut_35.scala 1065:39]
  wire  _GEN_14354 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13972; // @[lut_35.scala 1036:74 lut_35.scala 1066:39]
  wire  _GEN_14355 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13973; // @[lut_35.scala 1036:74 lut_35.scala 1067:39]
  wire  _GEN_14356 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13974; // @[lut_35.scala 1036:74 lut_35.scala 1068:39]
  wire  _GEN_14357 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13975; // @[lut_35.scala 1036:74 lut_35.scala 1069:39]
  wire  _GEN_14358 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13976; // @[lut_35.scala 1036:74 lut_35.scala 1070:39]
  wire  _GEN_14359 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13977; // @[lut_35.scala 1036:74 lut_35.scala 1071:39]
  wire  _GEN_14360 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid | _GEN_13978; // @[lut_35.scala 1036:74 lut_35.scala 1072:34]
  wire  _GEN_14364 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 1036:74 lut_35.scala 177:26 lut_35.scala 1074:27]
  wire  _GEN_14367 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13982; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14370 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13985; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14373 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13988; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14376 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13991; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14379 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13994; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14382 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13997; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14385 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14000; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14388 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14003; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14391 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14006; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14394 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14009; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14397 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14012; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14400 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14015; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14403 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14018; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14406 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14021; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14409 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14024; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14412 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14027; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14415 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14030; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14418 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14033; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14421 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14036; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14424 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14039; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14427 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14042; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14430 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14045; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14433 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14048; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14441 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14056; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14448 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14063; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14456 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14071; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14464 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14079; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14472 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14087; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14480 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14095; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14488 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14103; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14496 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14111; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14504 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14119; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14512 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14127; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14520 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14135; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14523 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_13954; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14528 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14143; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14531 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14146; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14536 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14151; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14539 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14154; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14544 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14159; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14547 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14162; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14552 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14167; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14555 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14170; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14560 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14175; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14563 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14178; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14568 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14183; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14571 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14186; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14576 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14191; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14579 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14194; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14584 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14199; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14587 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14202; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14592 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14207; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14595 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14210; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14600 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14215; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14603 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14218; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14608 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14223; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14611 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14226; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14616 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14231; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14619 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14234; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14624 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14239; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14627 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14242; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14632 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14247; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14635 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14250; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14640 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14255; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14643 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14258; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14648 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14263; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14651 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14266; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14656 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14271; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14659 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14274; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14664 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14279; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14667 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14282; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14672 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14287; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14675 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14290; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14680 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14295; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14683 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14298; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14688 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14303; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14691 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14306; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14696 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14311; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14699 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14314; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14704 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14319; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14707 = LUT_mem_MPORT_186_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14322; // @[lut_35.scala 1036:74 lut_35.scala 177:26]
  wire  _GEN_14710 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14325; // @[lut_35.scala 998:74 lut_35.scala 999:38]
  wire  _GEN_14711 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14326; // @[lut_35.scala 998:74 lut_35.scala 1000:38]
  wire  _GEN_14712 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14327; // @[lut_35.scala 998:74 lut_35.scala 1001:38]
  wire  _GEN_14713 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14328; // @[lut_35.scala 998:74 lut_35.scala 1002:38]
  wire  _GEN_14714 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14329; // @[lut_35.scala 998:74 lut_35.scala 1003:38]
  wire  _GEN_14715 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14330; // @[lut_35.scala 998:74 lut_35.scala 1004:38]
  wire  _GEN_14716 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14331; // @[lut_35.scala 998:74 lut_35.scala 1005:38]
  wire  _GEN_14717 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14332; // @[lut_35.scala 998:74 lut_35.scala 1006:38]
  wire  _GEN_14718 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14333; // @[lut_35.scala 998:74 lut_35.scala 1007:38]
  wire  _GEN_14719 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14334; // @[lut_35.scala 998:74 lut_35.scala 1008:38]
  wire  _GEN_14720 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid | _GEN_14335; // @[lut_35.scala 998:74 lut_35.scala 1009:39]
  wire  _GEN_14721 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14336; // @[lut_35.scala 998:74 lut_35.scala 1010:39]
  wire  _GEN_14722 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14337; // @[lut_35.scala 998:74 lut_35.scala 1011:39]
  wire  _GEN_14723 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14338; // @[lut_35.scala 998:74 lut_35.scala 1012:39]
  wire  _GEN_14724 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14339; // @[lut_35.scala 998:74 lut_35.scala 1013:39]
  wire  _GEN_14725 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14340; // @[lut_35.scala 998:74 lut_35.scala 1014:39]
  wire  _GEN_14726 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14341; // @[lut_35.scala 998:74 lut_35.scala 1015:39]
  wire  _GEN_14727 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14342; // @[lut_35.scala 998:74 lut_35.scala 1016:39]
  wire  _GEN_14728 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14343; // @[lut_35.scala 998:74 lut_35.scala 1017:39]
  wire  _GEN_14729 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14344; // @[lut_35.scala 998:74 lut_35.scala 1018:39]
  wire  _GEN_14730 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14345; // @[lut_35.scala 998:74 lut_35.scala 1019:39]
  wire  _GEN_14731 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14346; // @[lut_35.scala 998:74 lut_35.scala 1020:39]
  wire  _GEN_14732 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14347; // @[lut_35.scala 998:74 lut_35.scala 1021:39]
  wire  _GEN_14733 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14348; // @[lut_35.scala 998:74 lut_35.scala 1022:39]
  wire  _GEN_14734 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14349; // @[lut_35.scala 998:74 lut_35.scala 1023:39]
  wire  _GEN_14735 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14350; // @[lut_35.scala 998:74 lut_35.scala 1024:39]
  wire  _GEN_14736 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14351; // @[lut_35.scala 998:74 lut_35.scala 1025:39]
  wire  _GEN_14737 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14352; // @[lut_35.scala 998:74 lut_35.scala 1026:39]
  wire  _GEN_14738 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14353; // @[lut_35.scala 998:74 lut_35.scala 1027:39]
  wire  _GEN_14739 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14354; // @[lut_35.scala 998:74 lut_35.scala 1028:39]
  wire  _GEN_14740 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14355; // @[lut_35.scala 998:74 lut_35.scala 1029:39]
  wire  _GEN_14741 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14356; // @[lut_35.scala 998:74 lut_35.scala 1030:39]
  wire  _GEN_14742 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14357; // @[lut_35.scala 998:74 lut_35.scala 1031:39]
  wire  _GEN_14743 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14358; // @[lut_35.scala 998:74 lut_35.scala 1032:39]
  wire  _GEN_14744 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14359; // @[lut_35.scala 998:74 lut_35.scala 1033:39]
  wire  _GEN_14745 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid | _GEN_14360; // @[lut_35.scala 998:74 lut_35.scala 1034:34]
  wire  _GEN_14749 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 998:74 lut_35.scala 177:26 lut_35.scala 1036:27]
  wire  _GEN_14752 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14364; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14755 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14367; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14758 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14370; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14761 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14373; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14764 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14376; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14767 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14379; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14770 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14382; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14773 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14385; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14776 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14388; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14779 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14391; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14782 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14394; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14785 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14397; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14788 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14400; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14791 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14403; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14794 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14406; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14797 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14409; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14800 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14412; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14803 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14415; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14806 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14418; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14809 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14421; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14812 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14424; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14815 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14427; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14818 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14430; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14821 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14433; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14829 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14441; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14836 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14448; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14844 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14456; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14852 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14464; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14860 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14472; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14868 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14480; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14876 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14488; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14884 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14496; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14892 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14504; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14900 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14512; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14903 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14335; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14908 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14520; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14911 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14523; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14916 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14528; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14919 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14531; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14924 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14536; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14927 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14539; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14932 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14544; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14935 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14547; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14940 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14552; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14943 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14555; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14948 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14560; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14951 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14563; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14956 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14568; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14959 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14571; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14964 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14576; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14967 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14579; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14972 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14584; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14975 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14587; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14980 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14592; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14983 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14595; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14988 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14600; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14991 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14603; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14996 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14608; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_14999 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14611; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_15004 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14616; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_15007 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14619; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_15012 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14624; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_15015 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14627; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_15020 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14632; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_15023 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14635; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_15028 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14640; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_15031 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14643; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_15036 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14648; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_15039 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14651; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_15044 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14656; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_15047 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14659; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_15052 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14664; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_15055 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14667; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_15060 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14672; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_15063 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14675; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_15068 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14680; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_15071 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14683; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_15076 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14688; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_15079 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14691; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_15084 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14696; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_15087 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14699; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_15092 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14704; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_15095 = LUT_mem_MPORT_185_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14707; // @[lut_35.scala 998:74 lut_35.scala 177:26]
  wire  _GEN_15098 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14710; // @[lut_35.scala 960:73 lut_35.scala 961:38]
  wire  _GEN_15099 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14711; // @[lut_35.scala 960:73 lut_35.scala 962:38]
  wire  _GEN_15100 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14712; // @[lut_35.scala 960:73 lut_35.scala 963:38]
  wire  _GEN_15101 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14713; // @[lut_35.scala 960:73 lut_35.scala 964:38]
  wire  _GEN_15102 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14714; // @[lut_35.scala 960:73 lut_35.scala 965:38]
  wire  _GEN_15103 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14715; // @[lut_35.scala 960:73 lut_35.scala 966:38]
  wire  _GEN_15104 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14716; // @[lut_35.scala 960:73 lut_35.scala 967:38]
  wire  _GEN_15105 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14717; // @[lut_35.scala 960:73 lut_35.scala 968:38]
  wire  _GEN_15106 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14718; // @[lut_35.scala 960:73 lut_35.scala 969:38]
  wire  _GEN_15107 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid | _GEN_14719; // @[lut_35.scala 960:73 lut_35.scala 970:38]
  wire  _GEN_15108 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14720; // @[lut_35.scala 960:73 lut_35.scala 971:39]
  wire  _GEN_15109 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14721; // @[lut_35.scala 960:73 lut_35.scala 972:39]
  wire  _GEN_15110 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14722; // @[lut_35.scala 960:73 lut_35.scala 973:39]
  wire  _GEN_15111 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14723; // @[lut_35.scala 960:73 lut_35.scala 974:39]
  wire  _GEN_15112 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14724; // @[lut_35.scala 960:73 lut_35.scala 975:39]
  wire  _GEN_15113 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14725; // @[lut_35.scala 960:73 lut_35.scala 976:39]
  wire  _GEN_15114 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14726; // @[lut_35.scala 960:73 lut_35.scala 977:39]
  wire  _GEN_15115 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14727; // @[lut_35.scala 960:73 lut_35.scala 978:39]
  wire  _GEN_15116 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14728; // @[lut_35.scala 960:73 lut_35.scala 979:39]
  wire  _GEN_15117 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14729; // @[lut_35.scala 960:73 lut_35.scala 980:39]
  wire  _GEN_15118 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14730; // @[lut_35.scala 960:73 lut_35.scala 981:39]
  wire  _GEN_15119 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14731; // @[lut_35.scala 960:73 lut_35.scala 982:39]
  wire  _GEN_15120 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14732; // @[lut_35.scala 960:73 lut_35.scala 983:39]
  wire  _GEN_15121 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14733; // @[lut_35.scala 960:73 lut_35.scala 984:39]
  wire  _GEN_15122 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14734; // @[lut_35.scala 960:73 lut_35.scala 985:39]
  wire  _GEN_15123 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14735; // @[lut_35.scala 960:73 lut_35.scala 986:39]
  wire  _GEN_15124 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14736; // @[lut_35.scala 960:73 lut_35.scala 987:39]
  wire  _GEN_15125 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14737; // @[lut_35.scala 960:73 lut_35.scala 988:39]
  wire  _GEN_15126 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14738; // @[lut_35.scala 960:73 lut_35.scala 989:39]
  wire  _GEN_15127 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14739; // @[lut_35.scala 960:73 lut_35.scala 990:39]
  wire  _GEN_15128 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14740; // @[lut_35.scala 960:73 lut_35.scala 991:39]
  wire  _GEN_15129 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14741; // @[lut_35.scala 960:73 lut_35.scala 992:39]
  wire  _GEN_15130 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14742; // @[lut_35.scala 960:73 lut_35.scala 993:39]
  wire  _GEN_15131 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14743; // @[lut_35.scala 960:73 lut_35.scala 994:39]
  wire  _GEN_15132 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14744; // @[lut_35.scala 960:73 lut_35.scala 995:39]
  wire  _GEN_15133 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid | _GEN_14745; // @[lut_35.scala 960:73 lut_35.scala 996:34]
  wire  _GEN_15137 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 960:73 lut_35.scala 177:26 lut_35.scala 998:27]
  wire  _GEN_15140 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14749; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15143 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14752; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15146 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14755; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15149 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14758; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15152 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14761; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15155 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14764; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15158 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14767; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15161 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14770; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15164 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14773; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15167 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14776; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15170 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14779; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15173 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14782; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15176 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14785; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15179 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14788; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15182 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14791; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15185 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14794; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15188 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14797; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15191 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14800; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15194 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14803; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15197 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14806; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15200 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14809; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15203 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14812; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15206 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14815; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15209 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14818; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15212 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14821; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15220 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14829; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15227 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14836; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15235 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14844; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15243 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14852; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15251 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14860; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15259 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14868; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15267 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14876; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15275 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14884; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15283 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14892; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15286 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14719; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15291 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14900; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15294 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14903; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15299 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14908; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15302 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14911; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15307 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14916; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15310 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14919; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15315 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14924; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15318 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14927; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15323 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14932; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15326 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14935; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15331 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14940; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15334 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14943; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15339 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14948; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15342 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14951; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15347 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14956; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15350 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14959; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15355 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14964; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15358 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14967; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15363 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14972; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15366 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14975; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15371 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14980; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15374 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14983; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15379 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14988; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15382 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14991; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15387 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14996; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15390 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_14999; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15395 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15004; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15398 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15007; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15403 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15012; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15406 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15015; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15411 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15020; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15414 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15023; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15419 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15028; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15422 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15031; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15427 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15036; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15430 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15039; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15435 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15044; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15438 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15047; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15443 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15052; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15446 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15055; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15451 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15060; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15454 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15063; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15459 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15068; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15462 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15071; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15467 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15076; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15470 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15079; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15475 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15084; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15478 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15087; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15483 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15092; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15486 = LUT_mem_MPORT_184_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15095; // @[lut_35.scala 960:73 lut_35.scala 177:26]
  wire  _GEN_15489 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15098; // @[lut_35.scala 922:73 lut_35.scala 923:38]
  wire  _GEN_15490 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15099; // @[lut_35.scala 922:73 lut_35.scala 924:38]
  wire  _GEN_15491 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15100; // @[lut_35.scala 922:73 lut_35.scala 925:38]
  wire  _GEN_15492 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15101; // @[lut_35.scala 922:73 lut_35.scala 926:38]
  wire  _GEN_15493 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15102; // @[lut_35.scala 922:73 lut_35.scala 927:38]
  wire  _GEN_15494 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15103; // @[lut_35.scala 922:73 lut_35.scala 928:38]
  wire  _GEN_15495 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15104; // @[lut_35.scala 922:73 lut_35.scala 929:38]
  wire  _GEN_15496 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15105; // @[lut_35.scala 922:73 lut_35.scala 930:38]
  wire  _GEN_15497 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid | _GEN_15106; // @[lut_35.scala 922:73 lut_35.scala 931:38]
  wire  _GEN_15498 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15107; // @[lut_35.scala 922:73 lut_35.scala 932:38]
  wire  _GEN_15499 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15108; // @[lut_35.scala 922:73 lut_35.scala 933:39]
  wire  _GEN_15500 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15109; // @[lut_35.scala 922:73 lut_35.scala 934:39]
  wire  _GEN_15501 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15110; // @[lut_35.scala 922:73 lut_35.scala 935:39]
  wire  _GEN_15502 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15111; // @[lut_35.scala 922:73 lut_35.scala 936:39]
  wire  _GEN_15503 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15112; // @[lut_35.scala 922:73 lut_35.scala 937:39]
  wire  _GEN_15504 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15113; // @[lut_35.scala 922:73 lut_35.scala 938:39]
  wire  _GEN_15505 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15114; // @[lut_35.scala 922:73 lut_35.scala 939:39]
  wire  _GEN_15506 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15115; // @[lut_35.scala 922:73 lut_35.scala 940:39]
  wire  _GEN_15507 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15116; // @[lut_35.scala 922:73 lut_35.scala 941:39]
  wire  _GEN_15508 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15117; // @[lut_35.scala 922:73 lut_35.scala 942:39]
  wire  _GEN_15509 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15118; // @[lut_35.scala 922:73 lut_35.scala 943:39]
  wire  _GEN_15510 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15119; // @[lut_35.scala 922:73 lut_35.scala 944:39]
  wire  _GEN_15511 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15120; // @[lut_35.scala 922:73 lut_35.scala 945:39]
  wire  _GEN_15512 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15121; // @[lut_35.scala 922:73 lut_35.scala 946:39]
  wire  _GEN_15513 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15122; // @[lut_35.scala 922:73 lut_35.scala 947:39]
  wire  _GEN_15514 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15123; // @[lut_35.scala 922:73 lut_35.scala 948:39]
  wire  _GEN_15515 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15124; // @[lut_35.scala 922:73 lut_35.scala 949:39]
  wire  _GEN_15516 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15125; // @[lut_35.scala 922:73 lut_35.scala 950:39]
  wire  _GEN_15517 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15126; // @[lut_35.scala 922:73 lut_35.scala 951:39]
  wire  _GEN_15518 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15127; // @[lut_35.scala 922:73 lut_35.scala 952:39]
  wire  _GEN_15519 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15128; // @[lut_35.scala 922:73 lut_35.scala 953:39]
  wire  _GEN_15520 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15129; // @[lut_35.scala 922:73 lut_35.scala 954:39]
  wire  _GEN_15521 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15130; // @[lut_35.scala 922:73 lut_35.scala 955:39]
  wire  _GEN_15522 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15131; // @[lut_35.scala 922:73 lut_35.scala 956:39]
  wire  _GEN_15523 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15132; // @[lut_35.scala 922:73 lut_35.scala 957:39]
  wire  _GEN_15524 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid | _GEN_15133; // @[lut_35.scala 922:73 lut_35.scala 958:34]
  wire  _GEN_15528 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 922:73 lut_35.scala 177:26 lut_35.scala 960:27]
  wire  _GEN_15531 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15137; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15534 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15140; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15537 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15143; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15540 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15146; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15543 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15149; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15546 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15152; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15549 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15155; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15552 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15158; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15555 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15161; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15558 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15164; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15561 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15167; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15564 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15170; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15567 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15173; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15570 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15176; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15573 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15179; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15576 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15182; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15579 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15185; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15582 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15188; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15585 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15191; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15588 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15194; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15591 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15197; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15594 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15200; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15597 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15203; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15600 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15206; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15603 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15209; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15606 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15212; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15614 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15220; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15621 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15227; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15629 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15235; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15637 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15243; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15645 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15251; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15653 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15259; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15661 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15267; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15669 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15275; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15672 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15106; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15677 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15283; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15680 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15286; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15685 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15291; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15688 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15294; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15693 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15299; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15696 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15302; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15701 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15307; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15704 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15310; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15709 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15315; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15712 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15318; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15717 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15323; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15720 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15326; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15725 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15331; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15728 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15334; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15733 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15339; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15736 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15342; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15741 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15347; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15744 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15350; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15749 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15355; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15752 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15358; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15757 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15363; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15760 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15366; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15765 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15371; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15768 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15374; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15773 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15379; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15776 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15382; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15781 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15387; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15784 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15390; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15789 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15395; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15792 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15398; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15797 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15403; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15800 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15406; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15805 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15411; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15808 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15414; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15813 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15419; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15816 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15422; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15821 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15427; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15824 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15430; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15829 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15435; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15832 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15438; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15837 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15443; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15840 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15446; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15845 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15451; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15848 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15454; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15853 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15459; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15856 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15462; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15861 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15467; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15864 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15470; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15869 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15475; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15872 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15478; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15877 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15483; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15880 = LUT_mem_MPORT_183_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15486; // @[lut_35.scala 922:73 lut_35.scala 177:26]
  wire  _GEN_15883 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15489; // @[lut_35.scala 884:73 lut_35.scala 885:38]
  wire  _GEN_15884 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15490; // @[lut_35.scala 884:73 lut_35.scala 886:38]
  wire  _GEN_15885 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15491; // @[lut_35.scala 884:73 lut_35.scala 887:38]
  wire  _GEN_15886 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15492; // @[lut_35.scala 884:73 lut_35.scala 888:38]
  wire  _GEN_15887 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15493; // @[lut_35.scala 884:73 lut_35.scala 889:38]
  wire  _GEN_15888 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15494; // @[lut_35.scala 884:73 lut_35.scala 890:38]
  wire  _GEN_15889 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15495; // @[lut_35.scala 884:73 lut_35.scala 891:38]
  wire  _GEN_15890 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid | _GEN_15496; // @[lut_35.scala 884:73 lut_35.scala 892:38]
  wire  _GEN_15891 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15497; // @[lut_35.scala 884:73 lut_35.scala 893:38]
  wire  _GEN_15892 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15498; // @[lut_35.scala 884:73 lut_35.scala 894:38]
  wire  _GEN_15893 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15499; // @[lut_35.scala 884:73 lut_35.scala 895:39]
  wire  _GEN_15894 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15500; // @[lut_35.scala 884:73 lut_35.scala 896:39]
  wire  _GEN_15895 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15501; // @[lut_35.scala 884:73 lut_35.scala 897:39]
  wire  _GEN_15896 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15502; // @[lut_35.scala 884:73 lut_35.scala 898:39]
  wire  _GEN_15897 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15503; // @[lut_35.scala 884:73 lut_35.scala 899:39]
  wire  _GEN_15898 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15504; // @[lut_35.scala 884:73 lut_35.scala 900:39]
  wire  _GEN_15899 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15505; // @[lut_35.scala 884:73 lut_35.scala 901:39]
  wire  _GEN_15900 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15506; // @[lut_35.scala 884:73 lut_35.scala 902:39]
  wire  _GEN_15901 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15507; // @[lut_35.scala 884:73 lut_35.scala 903:39]
  wire  _GEN_15902 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15508; // @[lut_35.scala 884:73 lut_35.scala 904:39]
  wire  _GEN_15903 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15509; // @[lut_35.scala 884:73 lut_35.scala 905:39]
  wire  _GEN_15904 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15510; // @[lut_35.scala 884:73 lut_35.scala 906:39]
  wire  _GEN_15905 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15511; // @[lut_35.scala 884:73 lut_35.scala 907:39]
  wire  _GEN_15906 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15512; // @[lut_35.scala 884:73 lut_35.scala 908:39]
  wire  _GEN_15907 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15513; // @[lut_35.scala 884:73 lut_35.scala 909:39]
  wire  _GEN_15908 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15514; // @[lut_35.scala 884:73 lut_35.scala 910:39]
  wire  _GEN_15909 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15515; // @[lut_35.scala 884:73 lut_35.scala 911:39]
  wire  _GEN_15910 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15516; // @[lut_35.scala 884:73 lut_35.scala 912:39]
  wire  _GEN_15911 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15517; // @[lut_35.scala 884:73 lut_35.scala 913:39]
  wire  _GEN_15912 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15518; // @[lut_35.scala 884:73 lut_35.scala 914:39]
  wire  _GEN_15913 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15519; // @[lut_35.scala 884:73 lut_35.scala 915:39]
  wire  _GEN_15914 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15520; // @[lut_35.scala 884:73 lut_35.scala 916:39]
  wire  _GEN_15915 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15521; // @[lut_35.scala 884:73 lut_35.scala 917:39]
  wire  _GEN_15916 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15522; // @[lut_35.scala 884:73 lut_35.scala 918:39]
  wire  _GEN_15917 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15523; // @[lut_35.scala 884:73 lut_35.scala 919:39]
  wire  _GEN_15918 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid | _GEN_15524; // @[lut_35.scala 884:73 lut_35.scala 920:34]
  wire  _GEN_15922 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 884:73 lut_35.scala 177:26 lut_35.scala 922:27]
  wire  _GEN_15925 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15528; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_15928 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15531; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_15931 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15534; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_15934 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15537; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_15937 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15540; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_15940 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15543; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_15943 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15546; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_15946 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15549; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_15949 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15552; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_15952 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15555; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_15955 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15558; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_15958 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15561; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_15961 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15564; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_15964 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15567; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_15967 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15570; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_15970 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15573; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_15973 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15576; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_15976 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15579; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_15979 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15582; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_15982 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15585; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_15985 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15588; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_15988 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15591; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_15991 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15594; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_15994 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15597; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_15997 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15600; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16000 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15603; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16003 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15606; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16011 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15614; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16018 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15621; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16026 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15629; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16034 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15637; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16042 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15645; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16050 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15653; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16058 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15661; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16061 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15496; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16066 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15669; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16069 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15672; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16074 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15677; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16077 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15680; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16082 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15685; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16085 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15688; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16090 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15693; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16093 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15696; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16098 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15701; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16101 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15704; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16106 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15709; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16109 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15712; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16114 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15717; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16117 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15720; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16122 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15725; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16125 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15728; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16130 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15733; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16133 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15736; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16138 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15741; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16141 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15744; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16146 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15749; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16149 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15752; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16154 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15757; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16157 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15760; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16162 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15765; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16165 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15768; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16170 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15773; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16173 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15776; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16178 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15781; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16181 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15784; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16186 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15789; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16189 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15792; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16194 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15797; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16197 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15800; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16202 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15805; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16205 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15808; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16210 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15813; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16213 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15816; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16218 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15821; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16221 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15824; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16226 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15829; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16229 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15832; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16234 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15837; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16237 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15840; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16242 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15845; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16245 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15848; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16250 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15853; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16253 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15856; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16258 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15861; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16261 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15864; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16266 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15869; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16269 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15872; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16274 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15877; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16277 = LUT_mem_MPORT_182_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15880; // @[lut_35.scala 884:73 lut_35.scala 177:26]
  wire  _GEN_16280 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15883; // @[lut_35.scala 846:73 lut_35.scala 847:38]
  wire  _GEN_16281 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15884; // @[lut_35.scala 846:73 lut_35.scala 848:38]
  wire  _GEN_16282 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15885; // @[lut_35.scala 846:73 lut_35.scala 849:38]
  wire  _GEN_16283 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15886; // @[lut_35.scala 846:73 lut_35.scala 850:38]
  wire  _GEN_16284 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15887; // @[lut_35.scala 846:73 lut_35.scala 851:38]
  wire  _GEN_16285 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15888; // @[lut_35.scala 846:73 lut_35.scala 852:38]
  wire  _GEN_16286 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid | _GEN_15889; // @[lut_35.scala 846:73 lut_35.scala 853:38]
  wire  _GEN_16287 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15890; // @[lut_35.scala 846:73 lut_35.scala 854:38]
  wire  _GEN_16288 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15891; // @[lut_35.scala 846:73 lut_35.scala 855:38]
  wire  _GEN_16289 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15892; // @[lut_35.scala 846:73 lut_35.scala 856:38]
  wire  _GEN_16290 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15893; // @[lut_35.scala 846:73 lut_35.scala 857:39]
  wire  _GEN_16291 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15894; // @[lut_35.scala 846:73 lut_35.scala 858:39]
  wire  _GEN_16292 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15895; // @[lut_35.scala 846:73 lut_35.scala 859:39]
  wire  _GEN_16293 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15896; // @[lut_35.scala 846:73 lut_35.scala 860:39]
  wire  _GEN_16294 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15897; // @[lut_35.scala 846:73 lut_35.scala 861:39]
  wire  _GEN_16295 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15898; // @[lut_35.scala 846:73 lut_35.scala 862:39]
  wire  _GEN_16296 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15899; // @[lut_35.scala 846:73 lut_35.scala 863:39]
  wire  _GEN_16297 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15900; // @[lut_35.scala 846:73 lut_35.scala 864:39]
  wire  _GEN_16298 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15901; // @[lut_35.scala 846:73 lut_35.scala 865:39]
  wire  _GEN_16299 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15902; // @[lut_35.scala 846:73 lut_35.scala 866:39]
  wire  _GEN_16300 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15903; // @[lut_35.scala 846:73 lut_35.scala 867:39]
  wire  _GEN_16301 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15904; // @[lut_35.scala 846:73 lut_35.scala 868:39]
  wire  _GEN_16302 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15905; // @[lut_35.scala 846:73 lut_35.scala 869:39]
  wire  _GEN_16303 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15906; // @[lut_35.scala 846:73 lut_35.scala 870:39]
  wire  _GEN_16304 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15907; // @[lut_35.scala 846:73 lut_35.scala 871:39]
  wire  _GEN_16305 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15908; // @[lut_35.scala 846:73 lut_35.scala 872:39]
  wire  _GEN_16306 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15909; // @[lut_35.scala 846:73 lut_35.scala 873:39]
  wire  _GEN_16307 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15910; // @[lut_35.scala 846:73 lut_35.scala 874:39]
  wire  _GEN_16308 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15911; // @[lut_35.scala 846:73 lut_35.scala 875:39]
  wire  _GEN_16309 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15912; // @[lut_35.scala 846:73 lut_35.scala 876:39]
  wire  _GEN_16310 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15913; // @[lut_35.scala 846:73 lut_35.scala 877:39]
  wire  _GEN_16311 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15914; // @[lut_35.scala 846:73 lut_35.scala 878:39]
  wire  _GEN_16312 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15915; // @[lut_35.scala 846:73 lut_35.scala 879:39]
  wire  _GEN_16313 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15916; // @[lut_35.scala 846:73 lut_35.scala 880:39]
  wire  _GEN_16314 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15917; // @[lut_35.scala 846:73 lut_35.scala 881:39]
  wire  _GEN_16315 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid | _GEN_15918; // @[lut_35.scala 846:73 lut_35.scala 882:34]
  wire  _GEN_16319 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 846:73 lut_35.scala 177:26 lut_35.scala 884:27]
  wire  _GEN_16322 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15922; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16325 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15925; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16328 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15928; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16331 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15931; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16334 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15934; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16337 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15937; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16340 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15940; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16343 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15943; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16346 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15946; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16349 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15949; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16352 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15952; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16355 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15955; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16358 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15958; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16361 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15961; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16364 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15964; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16367 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15967; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16370 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15970; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16373 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15973; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16376 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15976; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16379 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15979; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16382 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15982; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16385 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15985; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16388 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15988; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16391 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15991; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16394 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15994; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16397 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15997; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16400 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16000; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16403 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16003; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16411 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16011; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16418 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16018; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16426 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16026; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16434 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16034; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16442 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16042; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16450 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16050; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16453 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_15889; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16458 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16058; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16461 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16061; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16466 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16066; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16469 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16069; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16474 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16074; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16477 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16077; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16482 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16082; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16485 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16085; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16490 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16090; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16493 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16093; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16498 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16098; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16501 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16101; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16506 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16106; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16509 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16109; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16514 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16114; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16517 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16117; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16522 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16122; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16525 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16125; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16530 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16130; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16533 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16133; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16538 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16138; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16541 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16141; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16546 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16146; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16549 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16149; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16554 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16154; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16557 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16157; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16562 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16162; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16565 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16165; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16570 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16170; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16573 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16173; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16578 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16178; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16581 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16181; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16586 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16186; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16589 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16189; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16594 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16194; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16597 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16197; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16602 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16202; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16605 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16205; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16610 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16210; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16613 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16213; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16618 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16218; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16621 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16221; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16626 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16226; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16629 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16229; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16634 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16234; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16637 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16237; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16642 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16242; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16645 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16245; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16650 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16250; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16653 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16253; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16658 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16258; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16661 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16261; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16666 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16266; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16669 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16269; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16674 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16274; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16677 = LUT_mem_MPORT_181_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16277; // @[lut_35.scala 846:73 lut_35.scala 177:26]
  wire  _GEN_16680 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16280; // @[lut_35.scala 808:73 lut_35.scala 809:38]
  wire  _GEN_16681 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16281; // @[lut_35.scala 808:73 lut_35.scala 810:38]
  wire  _GEN_16682 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16282; // @[lut_35.scala 808:73 lut_35.scala 811:38]
  wire  _GEN_16683 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16283; // @[lut_35.scala 808:73 lut_35.scala 812:38]
  wire  _GEN_16684 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16284; // @[lut_35.scala 808:73 lut_35.scala 813:38]
  wire  _GEN_16685 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid | _GEN_16285; // @[lut_35.scala 808:73 lut_35.scala 814:38]
  wire  _GEN_16686 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16286; // @[lut_35.scala 808:73 lut_35.scala 815:38]
  wire  _GEN_16687 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16287; // @[lut_35.scala 808:73 lut_35.scala 816:38]
  wire  _GEN_16688 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16288; // @[lut_35.scala 808:73 lut_35.scala 817:38]
  wire  _GEN_16689 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16289; // @[lut_35.scala 808:73 lut_35.scala 818:38]
  wire  _GEN_16690 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16290; // @[lut_35.scala 808:73 lut_35.scala 819:39]
  wire  _GEN_16691 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16291; // @[lut_35.scala 808:73 lut_35.scala 820:39]
  wire  _GEN_16692 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16292; // @[lut_35.scala 808:73 lut_35.scala 821:39]
  wire  _GEN_16693 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16293; // @[lut_35.scala 808:73 lut_35.scala 822:39]
  wire  _GEN_16694 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16294; // @[lut_35.scala 808:73 lut_35.scala 823:39]
  wire  _GEN_16695 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16295; // @[lut_35.scala 808:73 lut_35.scala 824:39]
  wire  _GEN_16696 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16296; // @[lut_35.scala 808:73 lut_35.scala 825:39]
  wire  _GEN_16697 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16297; // @[lut_35.scala 808:73 lut_35.scala 826:39]
  wire  _GEN_16698 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16298; // @[lut_35.scala 808:73 lut_35.scala 827:39]
  wire  _GEN_16699 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16299; // @[lut_35.scala 808:73 lut_35.scala 828:39]
  wire  _GEN_16700 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16300; // @[lut_35.scala 808:73 lut_35.scala 829:39]
  wire  _GEN_16701 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16301; // @[lut_35.scala 808:73 lut_35.scala 830:39]
  wire  _GEN_16702 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16302; // @[lut_35.scala 808:73 lut_35.scala 831:39]
  wire  _GEN_16703 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16303; // @[lut_35.scala 808:73 lut_35.scala 832:39]
  wire  _GEN_16704 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16304; // @[lut_35.scala 808:73 lut_35.scala 833:39]
  wire  _GEN_16705 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16305; // @[lut_35.scala 808:73 lut_35.scala 834:39]
  wire  _GEN_16706 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16306; // @[lut_35.scala 808:73 lut_35.scala 835:39]
  wire  _GEN_16707 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16307; // @[lut_35.scala 808:73 lut_35.scala 836:39]
  wire  _GEN_16708 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16308; // @[lut_35.scala 808:73 lut_35.scala 837:39]
  wire  _GEN_16709 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16309; // @[lut_35.scala 808:73 lut_35.scala 838:39]
  wire  _GEN_16710 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16310; // @[lut_35.scala 808:73 lut_35.scala 839:39]
  wire  _GEN_16711 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16311; // @[lut_35.scala 808:73 lut_35.scala 840:39]
  wire  _GEN_16712 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16312; // @[lut_35.scala 808:73 lut_35.scala 841:39]
  wire  _GEN_16713 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16313; // @[lut_35.scala 808:73 lut_35.scala 842:39]
  wire  _GEN_16714 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16314; // @[lut_35.scala 808:73 lut_35.scala 843:39]
  wire  _GEN_16715 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid | _GEN_16315; // @[lut_35.scala 808:73 lut_35.scala 844:34]
  wire  _GEN_16719 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 808:73 lut_35.scala 177:26 lut_35.scala 846:27]
  wire  _GEN_16722 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16319; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16725 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16322; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16728 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16325; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16731 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16328; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16734 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16331; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16737 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16334; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16740 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16337; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16743 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16340; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16746 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16343; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16749 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16346; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16752 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16349; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16755 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16352; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16758 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16355; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16761 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16358; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16764 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16361; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16767 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16364; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16770 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16367; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16773 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16370; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16776 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16373; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16779 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16376; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16782 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16379; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16785 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16382; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16788 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16385; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16791 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16388; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16794 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16391; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16797 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16394; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16800 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16397; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16803 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16400; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16806 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16403; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16814 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16411; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16821 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16418; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16829 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16426; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16837 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16434; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16845 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16442; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16848 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16285; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16853 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16450; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16856 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16453; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16861 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16458; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16864 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16461; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16869 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16466; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16872 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16469; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16877 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16474; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16880 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16477; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16885 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16482; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16888 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16485; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16893 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16490; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16896 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16493; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16901 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16498; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16904 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16501; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16909 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16506; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16912 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16509; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16917 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16514; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16920 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16517; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16925 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16522; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16928 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16525; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16933 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16530; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16936 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16533; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16941 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16538; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16944 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16541; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16949 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16546; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16952 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16549; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16957 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16554; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16960 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16557; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16965 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16562; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16968 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16565; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16973 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16570; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16976 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16573; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16981 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16578; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16984 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16581; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16989 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16586; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16992 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16589; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_16997 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16594; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_17000 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16597; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_17005 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16602; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_17008 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16605; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_17013 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16610; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_17016 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16613; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_17021 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16618; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_17024 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16621; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_17029 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16626; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_17032 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16629; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_17037 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16634; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_17040 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16637; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_17045 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16642; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_17048 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16645; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_17053 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16650; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_17056 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16653; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_17061 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16658; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_17064 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16661; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_17069 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16666; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_17072 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16669; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_17077 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16674; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_17080 = LUT_mem_MPORT_180_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16677; // @[lut_35.scala 808:73 lut_35.scala 177:26]
  wire  _GEN_17083 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16680; // @[lut_35.scala 770:73 lut_35.scala 771:38]
  wire  _GEN_17084 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16681; // @[lut_35.scala 770:73 lut_35.scala 772:38]
  wire  _GEN_17085 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16682; // @[lut_35.scala 770:73 lut_35.scala 773:38]
  wire  _GEN_17086 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16683; // @[lut_35.scala 770:73 lut_35.scala 774:38]
  wire  _GEN_17087 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid | _GEN_16684; // @[lut_35.scala 770:73 lut_35.scala 775:38]
  wire  _GEN_17088 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16685; // @[lut_35.scala 770:73 lut_35.scala 776:38]
  wire  _GEN_17089 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16686; // @[lut_35.scala 770:73 lut_35.scala 777:38]
  wire  _GEN_17090 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16687; // @[lut_35.scala 770:73 lut_35.scala 778:38]
  wire  _GEN_17091 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16688; // @[lut_35.scala 770:73 lut_35.scala 779:38]
  wire  _GEN_17092 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16689; // @[lut_35.scala 770:73 lut_35.scala 780:38]
  wire  _GEN_17093 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16690; // @[lut_35.scala 770:73 lut_35.scala 781:39]
  wire  _GEN_17094 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16691; // @[lut_35.scala 770:73 lut_35.scala 782:39]
  wire  _GEN_17095 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16692; // @[lut_35.scala 770:73 lut_35.scala 783:39]
  wire  _GEN_17096 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16693; // @[lut_35.scala 770:73 lut_35.scala 784:39]
  wire  _GEN_17097 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16694; // @[lut_35.scala 770:73 lut_35.scala 785:39]
  wire  _GEN_17098 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16695; // @[lut_35.scala 770:73 lut_35.scala 786:39]
  wire  _GEN_17099 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16696; // @[lut_35.scala 770:73 lut_35.scala 787:39]
  wire  _GEN_17100 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16697; // @[lut_35.scala 770:73 lut_35.scala 788:39]
  wire  _GEN_17101 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16698; // @[lut_35.scala 770:73 lut_35.scala 789:39]
  wire  _GEN_17102 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16699; // @[lut_35.scala 770:73 lut_35.scala 790:39]
  wire  _GEN_17103 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16700; // @[lut_35.scala 770:73 lut_35.scala 791:39]
  wire  _GEN_17104 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16701; // @[lut_35.scala 770:73 lut_35.scala 792:39]
  wire  _GEN_17105 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16702; // @[lut_35.scala 770:73 lut_35.scala 793:39]
  wire  _GEN_17106 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16703; // @[lut_35.scala 770:73 lut_35.scala 794:39]
  wire  _GEN_17107 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16704; // @[lut_35.scala 770:73 lut_35.scala 795:39]
  wire  _GEN_17108 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16705; // @[lut_35.scala 770:73 lut_35.scala 796:39]
  wire  _GEN_17109 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16706; // @[lut_35.scala 770:73 lut_35.scala 797:39]
  wire  _GEN_17110 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16707; // @[lut_35.scala 770:73 lut_35.scala 798:39]
  wire  _GEN_17111 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16708; // @[lut_35.scala 770:73 lut_35.scala 799:39]
  wire  _GEN_17112 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16709; // @[lut_35.scala 770:73 lut_35.scala 800:39]
  wire  _GEN_17113 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16710; // @[lut_35.scala 770:73 lut_35.scala 801:39]
  wire  _GEN_17114 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16711; // @[lut_35.scala 770:73 lut_35.scala 802:39]
  wire  _GEN_17115 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16712; // @[lut_35.scala 770:73 lut_35.scala 803:39]
  wire  _GEN_17116 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16713; // @[lut_35.scala 770:73 lut_35.scala 804:39]
  wire  _GEN_17117 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16714; // @[lut_35.scala 770:73 lut_35.scala 805:39]
  wire  _GEN_17118 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid | _GEN_16715; // @[lut_35.scala 770:73 lut_35.scala 806:34]
  wire  _GEN_17122 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 770:73 lut_35.scala 177:26 lut_35.scala 808:27]
  wire  _GEN_17125 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16719; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17128 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16722; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17131 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16725; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17134 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16728; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17137 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16731; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17140 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16734; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17143 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16737; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17146 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16740; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17149 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16743; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17152 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16746; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17155 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16749; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17158 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16752; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17161 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16755; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17164 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16758; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17167 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16761; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17170 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16764; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17173 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16767; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17176 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16770; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17179 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16773; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17182 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16776; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17185 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16779; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17188 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16782; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17191 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16785; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17194 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16788; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17197 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16791; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17200 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16794; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17203 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16797; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17206 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16800; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17209 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16803; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17212 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16806; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17220 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16814; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17227 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16821; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17235 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16829; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17243 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16837; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17246 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16684; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17251 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16845; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17254 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16848; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17259 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16853; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17262 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16856; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17267 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16861; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17270 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16864; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17275 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16869; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17278 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16872; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17283 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16877; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17286 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16880; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17291 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16885; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17294 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16888; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17299 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16893; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17302 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16896; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17307 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16901; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17310 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16904; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17315 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16909; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17318 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16912; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17323 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16917; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17326 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16920; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17331 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16925; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17334 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16928; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17339 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16933; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17342 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16936; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17347 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16941; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17350 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16944; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17355 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16949; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17358 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16952; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17363 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16957; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17366 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16960; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17371 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16965; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17374 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16968; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17379 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16973; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17382 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16976; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17387 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16981; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17390 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16984; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17395 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16989; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17398 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16992; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17403 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_16997; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17406 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17000; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17411 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17005; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17414 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17008; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17419 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17013; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17422 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17016; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17427 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17021; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17430 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17024; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17435 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17029; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17438 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17032; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17443 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17037; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17446 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17040; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17451 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17045; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17454 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17048; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17459 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17053; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17462 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17056; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17467 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17061; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17470 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17064; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17475 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17069; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17478 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17072; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17483 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17077; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17486 = LUT_mem_MPORT_179_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17080; // @[lut_35.scala 770:73 lut_35.scala 177:26]
  wire  _GEN_17489 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17083; // @[lut_35.scala 732:73 lut_35.scala 733:38]
  wire  _GEN_17490 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17084; // @[lut_35.scala 732:73 lut_35.scala 734:38]
  wire  _GEN_17491 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17085; // @[lut_35.scala 732:73 lut_35.scala 735:38]
  wire  _GEN_17492 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid | _GEN_17086; // @[lut_35.scala 732:73 lut_35.scala 736:38]
  wire  _GEN_17493 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17087; // @[lut_35.scala 732:73 lut_35.scala 737:38]
  wire  _GEN_17494 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17088; // @[lut_35.scala 732:73 lut_35.scala 738:38]
  wire  _GEN_17495 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17089; // @[lut_35.scala 732:73 lut_35.scala 739:38]
  wire  _GEN_17496 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17090; // @[lut_35.scala 732:73 lut_35.scala 740:38]
  wire  _GEN_17497 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17091; // @[lut_35.scala 732:73 lut_35.scala 741:38]
  wire  _GEN_17498 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17092; // @[lut_35.scala 732:73 lut_35.scala 742:38]
  wire  _GEN_17499 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17093; // @[lut_35.scala 732:73 lut_35.scala 743:39]
  wire  _GEN_17500 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17094; // @[lut_35.scala 732:73 lut_35.scala 744:39]
  wire  _GEN_17501 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17095; // @[lut_35.scala 732:73 lut_35.scala 745:39]
  wire  _GEN_17502 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17096; // @[lut_35.scala 732:73 lut_35.scala 746:39]
  wire  _GEN_17503 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17097; // @[lut_35.scala 732:73 lut_35.scala 747:39]
  wire  _GEN_17504 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17098; // @[lut_35.scala 732:73 lut_35.scala 748:39]
  wire  _GEN_17505 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17099; // @[lut_35.scala 732:73 lut_35.scala 749:39]
  wire  _GEN_17506 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17100; // @[lut_35.scala 732:73 lut_35.scala 750:39]
  wire  _GEN_17507 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17101; // @[lut_35.scala 732:73 lut_35.scala 751:39]
  wire  _GEN_17508 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17102; // @[lut_35.scala 732:73 lut_35.scala 752:39]
  wire  _GEN_17509 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17103; // @[lut_35.scala 732:73 lut_35.scala 753:39]
  wire  _GEN_17510 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17104; // @[lut_35.scala 732:73 lut_35.scala 754:39]
  wire  _GEN_17511 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17105; // @[lut_35.scala 732:73 lut_35.scala 755:39]
  wire  _GEN_17512 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17106; // @[lut_35.scala 732:73 lut_35.scala 756:39]
  wire  _GEN_17513 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17107; // @[lut_35.scala 732:73 lut_35.scala 757:39]
  wire  _GEN_17514 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17108; // @[lut_35.scala 732:73 lut_35.scala 758:39]
  wire  _GEN_17515 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17109; // @[lut_35.scala 732:73 lut_35.scala 759:39]
  wire  _GEN_17516 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17110; // @[lut_35.scala 732:73 lut_35.scala 760:39]
  wire  _GEN_17517 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17111; // @[lut_35.scala 732:73 lut_35.scala 761:39]
  wire  _GEN_17518 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17112; // @[lut_35.scala 732:73 lut_35.scala 762:39]
  wire  _GEN_17519 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17113; // @[lut_35.scala 732:73 lut_35.scala 763:39]
  wire  _GEN_17520 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17114; // @[lut_35.scala 732:73 lut_35.scala 764:39]
  wire  _GEN_17521 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17115; // @[lut_35.scala 732:73 lut_35.scala 765:39]
  wire  _GEN_17522 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17116; // @[lut_35.scala 732:73 lut_35.scala 766:39]
  wire  _GEN_17523 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17117; // @[lut_35.scala 732:73 lut_35.scala 767:39]
  wire  _GEN_17524 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid | _GEN_17118; // @[lut_35.scala 732:73 lut_35.scala 768:34]
  wire  _GEN_17528 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 732:73 lut_35.scala 177:26 lut_35.scala 770:27]
  wire  _GEN_17531 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17122; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17534 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17125; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17537 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17128; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17540 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17131; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17543 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17134; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17546 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17137; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17549 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17140; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17552 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17143; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17555 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17146; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17558 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17149; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17561 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17152; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17564 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17155; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17567 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17158; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17570 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17161; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17573 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17164; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17576 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17167; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17579 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17170; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17582 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17173; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17585 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17176; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17588 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17179; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17591 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17182; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17594 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17185; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17597 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17188; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17600 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17191; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17603 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17194; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17606 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17197; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17609 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17200; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17612 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17203; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17615 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17206; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17618 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17209; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17621 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17212; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17629 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17220; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17636 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17227; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17644 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17235; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17647 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17086; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17652 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17243; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17655 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17246; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17660 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17251; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17663 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17254; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17668 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17259; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17671 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17262; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17676 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17267; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17679 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17270; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17684 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17275; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17687 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17278; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17692 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17283; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17695 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17286; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17700 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17291; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17703 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17294; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17708 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17299; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17711 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17302; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17716 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17307; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17719 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17310; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17724 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17315; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17727 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17318; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17732 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17323; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17735 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17326; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17740 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17331; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17743 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17334; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17748 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17339; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17751 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17342; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17756 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17347; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17759 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17350; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17764 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17355; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17767 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17358; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17772 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17363; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17775 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17366; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17780 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17371; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17783 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17374; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17788 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17379; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17791 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17382; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17796 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17387; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17799 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17390; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17804 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17395; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17807 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17398; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17812 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17403; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17815 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17406; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17820 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17411; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17823 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17414; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17828 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17419; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17831 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17422; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17836 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17427; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17839 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17430; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17844 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17435; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17847 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17438; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17852 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17443; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17855 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17446; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17860 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17451; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17863 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17454; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17868 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17459; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17871 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17462; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17876 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17467; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17879 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17470; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17884 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17475; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17887 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17478; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17892 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17483; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17895 = LUT_mem_MPORT_178_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17486; // @[lut_35.scala 732:73 lut_35.scala 177:26]
  wire  _GEN_17898 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17489; // @[lut_35.scala 694:73 lut_35.scala 695:38]
  wire  _GEN_17899 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17490; // @[lut_35.scala 694:73 lut_35.scala 696:38]
  wire  _GEN_17900 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid | _GEN_17491; // @[lut_35.scala 694:73 lut_35.scala 697:38]
  wire  _GEN_17901 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17492; // @[lut_35.scala 694:73 lut_35.scala 698:38]
  wire  _GEN_17902 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17493; // @[lut_35.scala 694:73 lut_35.scala 699:38]
  wire  _GEN_17903 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17494; // @[lut_35.scala 694:73 lut_35.scala 700:38]
  wire  _GEN_17904 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17495; // @[lut_35.scala 694:73 lut_35.scala 701:38]
  wire  _GEN_17905 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17496; // @[lut_35.scala 694:73 lut_35.scala 702:38]
  wire  _GEN_17906 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17497; // @[lut_35.scala 694:73 lut_35.scala 703:38]
  wire  _GEN_17907 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17498; // @[lut_35.scala 694:73 lut_35.scala 704:38]
  wire  _GEN_17908 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17499; // @[lut_35.scala 694:73 lut_35.scala 705:39]
  wire  _GEN_17909 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17500; // @[lut_35.scala 694:73 lut_35.scala 706:39]
  wire  _GEN_17910 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17501; // @[lut_35.scala 694:73 lut_35.scala 707:39]
  wire  _GEN_17911 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17502; // @[lut_35.scala 694:73 lut_35.scala 708:39]
  wire  _GEN_17912 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17503; // @[lut_35.scala 694:73 lut_35.scala 709:39]
  wire  _GEN_17913 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17504; // @[lut_35.scala 694:73 lut_35.scala 710:39]
  wire  _GEN_17914 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17505; // @[lut_35.scala 694:73 lut_35.scala 711:39]
  wire  _GEN_17915 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17506; // @[lut_35.scala 694:73 lut_35.scala 712:39]
  wire  _GEN_17916 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17507; // @[lut_35.scala 694:73 lut_35.scala 713:39]
  wire  _GEN_17917 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17508; // @[lut_35.scala 694:73 lut_35.scala 714:39]
  wire  _GEN_17918 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17509; // @[lut_35.scala 694:73 lut_35.scala 715:39]
  wire  _GEN_17919 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17510; // @[lut_35.scala 694:73 lut_35.scala 716:39]
  wire  _GEN_17920 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17511; // @[lut_35.scala 694:73 lut_35.scala 717:39]
  wire  _GEN_17921 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17512; // @[lut_35.scala 694:73 lut_35.scala 718:39]
  wire  _GEN_17922 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17513; // @[lut_35.scala 694:73 lut_35.scala 719:39]
  wire  _GEN_17923 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17514; // @[lut_35.scala 694:73 lut_35.scala 720:39]
  wire  _GEN_17924 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17515; // @[lut_35.scala 694:73 lut_35.scala 721:39]
  wire  _GEN_17925 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17516; // @[lut_35.scala 694:73 lut_35.scala 722:39]
  wire  _GEN_17926 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17517; // @[lut_35.scala 694:73 lut_35.scala 723:39]
  wire  _GEN_17927 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17518; // @[lut_35.scala 694:73 lut_35.scala 724:39]
  wire  _GEN_17928 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17519; // @[lut_35.scala 694:73 lut_35.scala 725:39]
  wire  _GEN_17929 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17520; // @[lut_35.scala 694:73 lut_35.scala 726:39]
  wire  _GEN_17930 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17521; // @[lut_35.scala 694:73 lut_35.scala 727:39]
  wire  _GEN_17931 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17522; // @[lut_35.scala 694:73 lut_35.scala 728:39]
  wire  _GEN_17932 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17523; // @[lut_35.scala 694:73 lut_35.scala 729:39]
  wire  _GEN_17933 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid | _GEN_17524; // @[lut_35.scala 694:73 lut_35.scala 730:34]
  wire  _GEN_17937 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 694:73 lut_35.scala 177:26 lut_35.scala 732:27]
  wire  _GEN_17940 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17528; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_17943 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17531; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_17946 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17534; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_17949 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17537; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_17952 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17540; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_17955 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17543; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_17958 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17546; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_17961 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17549; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_17964 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17552; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_17967 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17555; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_17970 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17558; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_17973 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17561; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_17976 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17564; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_17979 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17567; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_17982 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17570; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_17985 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17573; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_17988 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17576; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_17991 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17579; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_17994 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17582; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_17997 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17585; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18000 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17588; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18003 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17591; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18006 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17594; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18009 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17597; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18012 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17600; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18015 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17603; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18018 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17606; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18021 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17609; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18024 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17612; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18027 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17615; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18030 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17618; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18033 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17621; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18041 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17629; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18048 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17636; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18051 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17491; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18056 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17644; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18059 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17647; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18064 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17652; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18067 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17655; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18072 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17660; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18075 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17663; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18080 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17668; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18083 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17671; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18088 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17676; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18091 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17679; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18096 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17684; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18099 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17687; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18104 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17692; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18107 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17695; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18112 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17700; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18115 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17703; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18120 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17708; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18123 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17711; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18128 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17716; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18131 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17719; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18136 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17724; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18139 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17727; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18144 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17732; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18147 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17735; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18152 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17740; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18155 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17743; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18160 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17748; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18163 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17751; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18168 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17756; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18171 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17759; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18176 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17764; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18179 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17767; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18184 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17772; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18187 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17775; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18192 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17780; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18195 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17783; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18200 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17788; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18203 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17791; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18208 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17796; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18211 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17799; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18216 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17804; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18219 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17807; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18224 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17812; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18227 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17815; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18232 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17820; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18235 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17823; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18240 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17828; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18243 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17831; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18248 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17836; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18251 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17839; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18256 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17844; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18259 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17847; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18264 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17852; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18267 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17855; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18272 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17860; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18275 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17863; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18280 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17868; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18283 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17871; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18288 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17876; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18291 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17879; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18296 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17884; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18299 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17887; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18304 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17892; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18307 = LUT_mem_MPORT_177_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17895; // @[lut_35.scala 694:73 lut_35.scala 177:26]
  wire  _GEN_18310 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17898; // @[lut_35.scala 656:74 lut_35.scala 657:38]
  wire  _GEN_18311 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid | _GEN_17899; // @[lut_35.scala 656:74 lut_35.scala 658:38]
  wire  _GEN_18312 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17900; // @[lut_35.scala 656:74 lut_35.scala 659:38]
  wire  _GEN_18313 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17901; // @[lut_35.scala 656:74 lut_35.scala 660:38]
  wire  _GEN_18314 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17902; // @[lut_35.scala 656:74 lut_35.scala 661:38]
  wire  _GEN_18315 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17903; // @[lut_35.scala 656:74 lut_35.scala 662:38]
  wire  _GEN_18316 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17904; // @[lut_35.scala 656:74 lut_35.scala 663:38]
  wire  _GEN_18317 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17905; // @[lut_35.scala 656:74 lut_35.scala 664:38]
  wire  _GEN_18318 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17906; // @[lut_35.scala 656:74 lut_35.scala 665:38]
  wire  _GEN_18319 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17907; // @[lut_35.scala 656:74 lut_35.scala 666:38]
  wire  _GEN_18320 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17908; // @[lut_35.scala 656:74 lut_35.scala 667:39]
  wire  _GEN_18321 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17909; // @[lut_35.scala 656:74 lut_35.scala 668:39]
  wire  _GEN_18322 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17910; // @[lut_35.scala 656:74 lut_35.scala 669:39]
  wire  _GEN_18323 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17911; // @[lut_35.scala 656:74 lut_35.scala 670:39]
  wire  _GEN_18324 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17912; // @[lut_35.scala 656:74 lut_35.scala 671:39]
  wire  _GEN_18325 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17913; // @[lut_35.scala 656:74 lut_35.scala 672:39]
  wire  _GEN_18326 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17914; // @[lut_35.scala 656:74 lut_35.scala 673:39]
  wire  _GEN_18327 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17915; // @[lut_35.scala 656:74 lut_35.scala 674:39]
  wire  _GEN_18328 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17916; // @[lut_35.scala 656:74 lut_35.scala 675:39]
  wire  _GEN_18329 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17917; // @[lut_35.scala 656:74 lut_35.scala 676:39]
  wire  _GEN_18330 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17918; // @[lut_35.scala 656:74 lut_35.scala 677:39]
  wire  _GEN_18331 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17919; // @[lut_35.scala 656:74 lut_35.scala 678:39]
  wire  _GEN_18332 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17920; // @[lut_35.scala 656:74 lut_35.scala 679:39]
  wire  _GEN_18333 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17921; // @[lut_35.scala 656:74 lut_35.scala 680:39]
  wire  _GEN_18334 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17922; // @[lut_35.scala 656:74 lut_35.scala 681:39]
  wire  _GEN_18335 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17923; // @[lut_35.scala 656:74 lut_35.scala 682:39]
  wire  _GEN_18336 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17924; // @[lut_35.scala 656:74 lut_35.scala 683:39]
  wire  _GEN_18337 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17925; // @[lut_35.scala 656:74 lut_35.scala 684:39]
  wire  _GEN_18338 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17926; // @[lut_35.scala 656:74 lut_35.scala 685:39]
  wire  _GEN_18339 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17927; // @[lut_35.scala 656:74 lut_35.scala 686:39]
  wire  _GEN_18340 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17928; // @[lut_35.scala 656:74 lut_35.scala 687:39]
  wire  _GEN_18341 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17929; // @[lut_35.scala 656:74 lut_35.scala 688:39]
  wire  _GEN_18342 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17930; // @[lut_35.scala 656:74 lut_35.scala 689:39]
  wire  _GEN_18343 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17931; // @[lut_35.scala 656:74 lut_35.scala 690:39]
  wire  _GEN_18344 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17932; // @[lut_35.scala 656:74 lut_35.scala 691:39]
  wire  _GEN_18345 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid | _GEN_17933; // @[lut_35.scala 656:74 lut_35.scala 692:34]
  wire  _GEN_18349 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 656:74 lut_35.scala 177:26 lut_35.scala 694:27]
  wire  _GEN_18352 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17937; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18355 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17940; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18358 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17943; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18361 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17946; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18364 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17949; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18367 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17952; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18370 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17955; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18373 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17958; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18376 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17961; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18379 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17964; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18382 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17967; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18385 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17970; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18388 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17973; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18391 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17976; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18394 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17979; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18397 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17982; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18400 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17985; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18403 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17988; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18406 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17991; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18409 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17994; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18412 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17997; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18415 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18000; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18418 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18003; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18421 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18006; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18424 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18009; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18427 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18012; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18430 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18015; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18433 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18018; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18436 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18021; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18439 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18024; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18442 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18027; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18445 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18030; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18448 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18033; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18456 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18041; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18459 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_17899; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18463 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18048; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18466 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18051; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18471 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18056; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18474 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18059; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18479 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18064; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18482 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18067; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18487 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18072; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18490 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18075; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18495 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18080; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18498 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18083; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18503 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18088; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18506 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18091; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18511 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18096; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18514 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18099; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18519 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18104; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18522 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18107; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18527 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18112; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18530 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18115; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18535 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18120; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18538 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18123; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18543 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18128; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18546 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18131; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18551 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18136; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18554 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18139; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18559 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18144; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18562 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18147; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18567 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18152; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18570 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18155; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18575 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18160; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18578 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18163; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18583 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18168; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18586 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18171; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18591 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18176; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18594 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18179; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18599 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18184; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18602 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18187; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18607 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18192; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18610 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18195; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18615 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18200; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18618 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18203; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18623 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18208; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18626 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18211; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18631 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18216; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18634 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18219; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18639 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18224; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18642 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18227; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18647 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18232; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18650 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18235; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18655 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18240; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18658 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18243; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18663 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18248; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18666 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18251; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18671 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18256; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18674 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18259; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18679 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18264; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18682 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18267; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18687 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18272; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18690 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18275; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18695 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18280; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18698 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18283; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18703 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18288; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18706 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18291; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18711 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18296; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18714 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18299; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18719 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18304; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18722 = LUT_mem_MPORT_176_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18307; // @[lut_35.scala 656:74 lut_35.scala 177:26]
  wire  _GEN_18725 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid | _GEN_18310; // @[lut_35.scala 618:68 lut_35.scala 619:38]
  wire  _GEN_18726 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18311; // @[lut_35.scala 618:68 lut_35.scala 620:38]
  wire  _GEN_18727 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18312; // @[lut_35.scala 618:68 lut_35.scala 621:38]
  wire  _GEN_18728 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18313; // @[lut_35.scala 618:68 lut_35.scala 622:38]
  wire  _GEN_18729 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18314; // @[lut_35.scala 618:68 lut_35.scala 623:38]
  wire  _GEN_18730 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18315; // @[lut_35.scala 618:68 lut_35.scala 624:38]
  wire  _GEN_18731 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18316; // @[lut_35.scala 618:68 lut_35.scala 625:38]
  wire  _GEN_18732 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18317; // @[lut_35.scala 618:68 lut_35.scala 626:38]
  wire  _GEN_18733 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18318; // @[lut_35.scala 618:68 lut_35.scala 627:38]
  wire  _GEN_18734 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18319; // @[lut_35.scala 618:68 lut_35.scala 628:38]
  wire  _GEN_18735 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18320; // @[lut_35.scala 618:68 lut_35.scala 629:39]
  wire  _GEN_18736 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18321; // @[lut_35.scala 618:68 lut_35.scala 630:39]
  wire  _GEN_18737 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18322; // @[lut_35.scala 618:68 lut_35.scala 631:39]
  wire  _GEN_18738 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18323; // @[lut_35.scala 618:68 lut_35.scala 632:39]
  wire  _GEN_18739 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18324; // @[lut_35.scala 618:68 lut_35.scala 633:39]
  wire  _GEN_18740 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18325; // @[lut_35.scala 618:68 lut_35.scala 634:39]
  wire  _GEN_18741 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18326; // @[lut_35.scala 618:68 lut_35.scala 635:39]
  wire  _GEN_18742 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18327; // @[lut_35.scala 618:68 lut_35.scala 636:39]
  wire  _GEN_18743 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18328; // @[lut_35.scala 618:68 lut_35.scala 637:39]
  wire  _GEN_18744 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18329; // @[lut_35.scala 618:68 lut_35.scala 638:39]
  wire  _GEN_18745 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18330; // @[lut_35.scala 618:68 lut_35.scala 639:39]
  wire  _GEN_18746 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18331; // @[lut_35.scala 618:68 lut_35.scala 640:39]
  wire  _GEN_18747 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18332; // @[lut_35.scala 618:68 lut_35.scala 641:39]
  wire  _GEN_18748 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18333; // @[lut_35.scala 618:68 lut_35.scala 642:39]
  wire  _GEN_18749 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18334; // @[lut_35.scala 618:68 lut_35.scala 643:39]
  wire  _GEN_18750 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18335; // @[lut_35.scala 618:68 lut_35.scala 644:39]
  wire  _GEN_18751 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18336; // @[lut_35.scala 618:68 lut_35.scala 645:39]
  wire  _GEN_18752 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18337; // @[lut_35.scala 618:68 lut_35.scala 646:39]
  wire  _GEN_18753 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18338; // @[lut_35.scala 618:68 lut_35.scala 647:39]
  wire  _GEN_18754 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18339; // @[lut_35.scala 618:68 lut_35.scala 648:39]
  wire  _GEN_18755 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18340; // @[lut_35.scala 618:68 lut_35.scala 649:39]
  wire  _GEN_18756 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18341; // @[lut_35.scala 618:68 lut_35.scala 650:39]
  wire  _GEN_18757 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18342; // @[lut_35.scala 618:68 lut_35.scala 651:39]
  wire  _GEN_18758 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18343; // @[lut_35.scala 618:68 lut_35.scala 652:39]
  wire  _GEN_18759 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18344; // @[lut_35.scala 618:68 lut_35.scala 653:39]
  wire  _GEN_18760 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid | _GEN_18345; // @[lut_35.scala 618:68 lut_35.scala 654:34]
  wire  _GEN_18764 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : 1'h1; // @[lut_35.scala 618:68 lut_35.scala 177:26 lut_35.scala 656:27]
  wire  _GEN_18767 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18349; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18770 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18352; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18773 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18355; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18776 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18358; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18779 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18361; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18782 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18364; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18785 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18367; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18788 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18370; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18791 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18373; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18794 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18376; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18797 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18379; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18800 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18382; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18803 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18385; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18806 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18388; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18809 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18391; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18812 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18394; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18815 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18397; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18818 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18400; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18821 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18403; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18824 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18406; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18827 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18409; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18830 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18412; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18833 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18415; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18836 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18418; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18839 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18421; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18842 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18424; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18845 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18427; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18848 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18430; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18851 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18433; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18854 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18436; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18857 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18439; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18860 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18442; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18863 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18445; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18866 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18448; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18869 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18310; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18874 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18456; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18877 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18459; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18881 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18463; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18884 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18466; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18889 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18471; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18892 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18474; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18897 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18479; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18900 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18482; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18905 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18487; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18908 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18490; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18913 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18495; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18916 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18498; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18921 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18503; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18924 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18506; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18929 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18511; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18932 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18514; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18937 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18519; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18940 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18522; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18945 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18527; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18948 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18530; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18953 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18535; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18956 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18538; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18961 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18543; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18964 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18546; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18969 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18551; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18972 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18554; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18977 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18559; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18980 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18562; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18985 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18567; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18988 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18570; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18993 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18575; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_18996 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18578; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_19001 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18583; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_19004 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18586; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_19009 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18591; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_19012 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18594; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_19017 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18599; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_19020 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18602; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_19025 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18607; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_19028 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18610; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_19033 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18615; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_19036 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18618; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_19041 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18623; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_19044 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18626; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_19049 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18631; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_19052 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18634; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_19057 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18639; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_19060 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18642; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_19065 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18647; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_19068 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18650; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_19073 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18655; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_19076 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18658; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_19081 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18663; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_19084 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18666; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_19089 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18671; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_19092 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18674; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_19097 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18679; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_19100 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18682; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_19105 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18687; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_19108 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18690; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_19113 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18695; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_19116 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18698; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_19121 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18703; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_19124 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18706; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_19129 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18711; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_19132 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18714; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_19137 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18719; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_19140 = LUT_mem_MPORT_175_data[31:0] == push_ray_id & push_valid ? 1'h0 : _GEN_18722; // @[lut_35.scala 618:68 lut_35.scala 177:26]
  wire  _GEN_19146 = push_1 & push_valid & _GEN_18725; // @[lut_35.scala 617:46 lut_35.scala 3432:32]
  wire  _GEN_19147 = push_1 & push_valid & _GEN_18726; // @[lut_35.scala 617:46 lut_35.scala 3433:32]
  wire  _GEN_19148 = push_1 & push_valid & _GEN_18727; // @[lut_35.scala 617:46 lut_35.scala 3434:32]
  wire  _GEN_19149 = push_1 & push_valid & _GEN_18728; // @[lut_35.scala 617:46 lut_35.scala 3435:32]
  wire  _GEN_19150 = push_1 & push_valid & _GEN_18729; // @[lut_35.scala 617:46 lut_35.scala 3436:32]
  wire  _GEN_19151 = push_1 & push_valid & _GEN_18730; // @[lut_35.scala 617:46 lut_35.scala 3437:32]
  wire  _GEN_19152 = push_1 & push_valid & _GEN_18731; // @[lut_35.scala 617:46 lut_35.scala 3438:32]
  wire  _GEN_19153 = push_1 & push_valid & _GEN_18732; // @[lut_35.scala 617:46 lut_35.scala 3439:32]
  wire  _GEN_19154 = push_1 & push_valid & _GEN_18733; // @[lut_35.scala 617:46 lut_35.scala 3440:42]
  wire  _GEN_19155 = push_1 & push_valid & _GEN_18734; // @[lut_35.scala 617:46 lut_35.scala 3441:42]
  wire  _GEN_19156 = push_1 & push_valid & _GEN_18735; // @[lut_35.scala 617:46 lut_35.scala 3442:43]
  wire  _GEN_19157 = push_1 & push_valid & _GEN_18736; // @[lut_35.scala 617:46 lut_35.scala 3443:43]
  wire  _GEN_19158 = push_1 & push_valid & _GEN_18737; // @[lut_35.scala 617:46 lut_35.scala 3444:43]
  wire  _GEN_19159 = push_1 & push_valid & _GEN_18738; // @[lut_35.scala 617:46 lut_35.scala 3445:43]
  wire  _GEN_19160 = push_1 & push_valid & _GEN_18739; // @[lut_35.scala 617:46 lut_35.scala 3446:43]
  wire  _GEN_19161 = push_1 & push_valid & _GEN_18740; // @[lut_35.scala 617:46 lut_35.scala 3447:43]
  wire  _GEN_19162 = push_1 & push_valid & _GEN_18741; // @[lut_35.scala 617:46 lut_35.scala 3448:43]
  wire  _GEN_19163 = push_1 & push_valid & _GEN_18742; // @[lut_35.scala 617:46 lut_35.scala 3449:43]
  wire  _GEN_19164 = push_1 & push_valid & _GEN_18743; // @[lut_35.scala 617:46 lut_35.scala 3450:43]
  wire  _GEN_19165 = push_1 & push_valid & _GEN_18744; // @[lut_35.scala 617:46 lut_35.scala 3451:43]
  wire  _GEN_19166 = push_1 & push_valid & _GEN_18745; // @[lut_35.scala 617:46 lut_35.scala 3452:43]
  wire  _GEN_19167 = push_1 & push_valid & _GEN_18746; // @[lut_35.scala 617:46 lut_35.scala 3453:43]
  wire  _GEN_19168 = push_1 & push_valid & _GEN_18747; // @[lut_35.scala 617:46 lut_35.scala 3454:43]
  wire  _GEN_19169 = push_1 & push_valid & _GEN_18748; // @[lut_35.scala 617:46 lut_35.scala 3455:43]
  wire  _GEN_19170 = push_1 & push_valid & _GEN_18749; // @[lut_35.scala 617:46 lut_35.scala 3456:43]
  wire  _GEN_19171 = push_1 & push_valid & _GEN_18750; // @[lut_35.scala 617:46 lut_35.scala 3457:43]
  wire  _GEN_19172 = push_1 & push_valid & _GEN_18751; // @[lut_35.scala 617:46 lut_35.scala 3458:43]
  wire  _GEN_19173 = push_1 & push_valid & _GEN_18752; // @[lut_35.scala 617:46 lut_35.scala 3459:43]
  wire  _GEN_19174 = push_1 & push_valid & _GEN_18753; // @[lut_35.scala 617:46 lut_35.scala 3460:43]
  wire  _GEN_19175 = push_1 & push_valid & _GEN_18754; // @[lut_35.scala 617:46 lut_35.scala 3461:43]
  wire  _GEN_19176 = push_1 & push_valid & _GEN_18755; // @[lut_35.scala 617:46 lut_35.scala 3462:43]
  wire  _GEN_19177 = push_1 & push_valid & _GEN_18756; // @[lut_35.scala 617:46 lut_35.scala 3463:43]
  wire  _GEN_19178 = push_1 & push_valid & _GEN_18757; // @[lut_35.scala 617:46 lut_35.scala 3464:43]
  wire  _GEN_19179 = push_1 & push_valid & _GEN_18758; // @[lut_35.scala 617:46 lut_35.scala 3465:43]
  wire  _GEN_19180 = push_1 & push_valid & _GEN_18759; // @[lut_35.scala 617:46 lut_35.scala 3466:43]
  wire  _GEN_19181 = push_1 & push_valid & _GEN_18760; // @[lut_35.scala 617:46 lut_35.scala 3467:30]
  reg  pop_1; // @[lut_35.scala 3532:50]
  reg [31:0] read_stack0_pop; // @[lut_35.scala 3533:38]
  reg [31:0] read_stack1_pop; // @[lut_35.scala 3534:38]
  reg [31:0] read_stack2_pop; // @[lut_35.scala 3535:38]
  reg [31:0] read_stack3_pop; // @[lut_35.scala 3536:38]
  reg [31:0] read_stack4_pop; // @[lut_35.scala 3537:38]
  reg [31:0] read_stack5_pop; // @[lut_35.scala 3538:38]
  reg [31:0] read_stack6_pop; // @[lut_35.scala 3539:38]
  reg [31:0] read_stack7_pop; // @[lut_35.scala 3540:38]
  reg [31:0] read_stack8_pop; // @[lut_35.scala 3541:38]
  reg [31:0] read_stack9_pop; // @[lut_35.scala 3542:38]
  reg [31:0] read_stack10_pop; // @[lut_35.scala 3543:39]
  reg [31:0] read_stack11_pop; // @[lut_35.scala 3544:39]
  reg [31:0] read_stack12_pop; // @[lut_35.scala 3545:39]
  reg [31:0] read_stack13_pop; // @[lut_35.scala 3546:39]
  reg [31:0] read_stack14_pop; // @[lut_35.scala 3547:39]
  reg [31:0] read_stack15_pop; // @[lut_35.scala 3548:39]
  reg [31:0] read_stack16_pop; // @[lut_35.scala 3549:39]
  reg [31:0] read_stack17_pop; // @[lut_35.scala 3550:39]
  reg [31:0] read_stack18_pop; // @[lut_35.scala 3551:39]
  reg [31:0] read_stack19_pop; // @[lut_35.scala 3552:39]
  reg [31:0] read_stack20_pop; // @[lut_35.scala 3553:39]
  reg [31:0] read_stack21_pop; // @[lut_35.scala 3554:39]
  reg [31:0] read_stack22_pop; // @[lut_35.scala 3555:39]
  reg [31:0] read_stack23_pop; // @[lut_35.scala 3556:39]
  reg [31:0] read_stack24_pop; // @[lut_35.scala 3557:39]
  reg [31:0] read_stack25_pop; // @[lut_35.scala 3558:39]
  reg [31:0] read_stack26_pop; // @[lut_35.scala 3559:39]
  reg [31:0] read_stack27_pop; // @[lut_35.scala 3560:39]
  reg [31:0] read_stack28_pop; // @[lut_35.scala 3561:39]
  reg [31:0] read_stack29_pop; // @[lut_35.scala 3562:39]
  reg [31:0] read_stack30_pop; // @[lut_35.scala 3563:39]
  reg [31:0] read_stack31_pop; // @[lut_35.scala 3564:39]
  reg [31:0] read_stack32_pop; // @[lut_35.scala 3565:39]
  reg [31:0] read_stack33_pop; // @[lut_35.scala 3566:39]
  reg [31:0] read_stack34_pop; // @[lut_35.scala 3567:39]
  reg [31:0] pop_ray_id; // @[lut_35.scala 3570:37]
  reg [31:0] pop_hitT_1; // @[lut_35.scala 3571:37]
  reg  pop_valid; // @[lut_35.scala 3572:36]
  reg  pop_0_1; // @[lut_35.scala 3575:46]
  reg  pop_1_1; // @[lut_35.scala 3576:46]
  reg  pop_2_1; // @[lut_35.scala 3577:46]
  reg  pop_3_1; // @[lut_35.scala 3578:46]
  reg  pop_4_1; // @[lut_35.scala 3579:46]
  reg  pop_5_1; // @[lut_35.scala 3580:46]
  reg  pop_6_1; // @[lut_35.scala 3581:46]
  reg  pop_7_1; // @[lut_35.scala 3582:46]
  reg  pop_8_1; // @[lut_35.scala 3583:46]
  reg  pop_9_1; // @[lut_35.scala 3584:46]
  reg  pop_10_1; // @[lut_35.scala 3585:47]
  reg  pop_11_1; // @[lut_35.scala 3586:47]
  reg  pop_12_1; // @[lut_35.scala 3587:47]
  reg  pop_13_1; // @[lut_35.scala 3588:47]
  reg  pop_14_1; // @[lut_35.scala 3589:47]
  reg  pop_15_1; // @[lut_35.scala 3590:47]
  reg  pop_16_1; // @[lut_35.scala 3591:47]
  reg  pop_17_1; // @[lut_35.scala 3592:47]
  reg  pop_18_1; // @[lut_35.scala 3593:47]
  reg  pop_19_1; // @[lut_35.scala 3594:47]
  reg  pop_20_1; // @[lut_35.scala 3595:47]
  reg  pop_21_1; // @[lut_35.scala 3596:47]
  reg  pop_22_1; // @[lut_35.scala 3597:47]
  reg  pop_23_1; // @[lut_35.scala 3598:47]
  reg  pop_24_1; // @[lut_35.scala 3599:47]
  reg  pop_25_1; // @[lut_35.scala 3600:47]
  reg  pop_26_1; // @[lut_35.scala 3601:47]
  reg  pop_27_1; // @[lut_35.scala 3602:47]
  reg  pop_28_1; // @[lut_35.scala 3603:47]
  reg  pop_29_1; // @[lut_35.scala 3604:47]
  reg  pop_30_1; // @[lut_35.scala 3605:47]
  reg  pop_31_1; // @[lut_35.scala 3606:47]
  reg  pop_32_1; // @[lut_35.scala 3607:47]
  reg  pop_33_1; // @[lut_35.scala 3608:47]
  reg  pop_34_1; // @[lut_35.scala 3609:47]
  reg  pop_valid_2; // @[lut_35.scala 3611:47]
  reg [31:0] pop_ray_id_2; // @[lut_35.scala 3613:47]
  reg [31:0] pop_hitT_2; // @[lut_35.scala 3614:47]
  reg  no_match; // @[lut_35.scala 3616:47]
  wire  _T_672 = io_pop & io_pop_valid; // @[lut_35.scala 3657:28]
  wire  _T_681 = pop_1 & pop_ray_id != read_stack0_pop & pop_ray_id != read_stack1_pop & pop_ray_id != read_stack2_pop
     & pop_ray_id != read_stack3_pop; // @[lut_35.scala 3669:124]
  wire  _T_689 = _T_681 & pop_ray_id != read_stack4_pop & pop_ray_id != read_stack5_pop & pop_ray_id != read_stack6_pop
     & pop_ray_id != read_stack7_pop; // @[lut_35.scala 3670:108]
  wire  _T_697 = _T_689 & pop_ray_id != read_stack8_pop & pop_ray_id != read_stack9_pop & pop_ray_id != read_stack10_pop
     & pop_ray_id != read_stack11_pop; // @[lut_35.scala 3671:109]
  wire  _T_705 = _T_697 & pop_ray_id != read_stack12_pop & pop_ray_id != read_stack13_pop & pop_ray_id !=
    read_stack14_pop & pop_ray_id != read_stack15_pop; // @[lut_35.scala 3672:111]
  wire  _T_713 = _T_705 & pop_ray_id != read_stack16_pop & pop_ray_id != read_stack17_pop & pop_ray_id !=
    read_stack18_pop & pop_ray_id != read_stack19_pop; // @[lut_35.scala 3673:111]
  wire  _T_721 = _T_713 & pop_ray_id != read_stack20_pop & pop_ray_id != read_stack21_pop & pop_ray_id !=
    read_stack22_pop & pop_ray_id != read_stack23_pop; // @[lut_35.scala 3674:111]
  wire  _T_729 = _T_721 & pop_ray_id != read_stack24_pop & pop_ray_id != read_stack25_pop & pop_ray_id !=
    read_stack26_pop & pop_ray_id != read_stack27_pop; // @[lut_35.scala 3675:111]
  wire  _T_736 = pop_ray_id != read_stack31_pop; // @[lut_35.scala 3676:125]
  wire  _T_737 = _T_729 & pop_ray_id != read_stack28_pop & pop_ray_id != read_stack29_pop & pop_ray_id !=
    read_stack30_pop & pop_ray_id != read_stack31_pop; // @[lut_35.scala 3676:111]
  wire  _T_745 = _T_737 & _T_736 & pop_ray_id != read_stack32_pop & pop_ray_id != read_stack33_pop & pop_ray_id !=
    read_stack34_pop; // @[lut_35.scala 3677:111]
  reg  no_match_1; // @[lut_35.scala 3682:51]
  reg  no_match_2; // @[lut_35.scala 3683:51]
  wire  _T_751 = read_stack0_pop == pop_ray_id & pop_valid; // @[lut_35.scala 3688:45]
  wire  _T_754 = read_stack1_pop == pop_ray_id & pop_valid; // @[lut_35.scala 3728:55]
  wire  _T_757 = read_stack2_pop == pop_ray_id & pop_valid; // @[lut_35.scala 3768:55]
  wire  _T_760 = read_stack3_pop == pop_ray_id & pop_valid; // @[lut_35.scala 3808:55]
  wire  _T_763 = read_stack4_pop == pop_ray_id & pop_valid; // @[lut_35.scala 3848:55]
  wire  _T_766 = read_stack5_pop == pop_ray_id & pop_valid; // @[lut_35.scala 3888:55]
  wire  _T_769 = read_stack6_pop == pop_ray_id & pop_valid; // @[lut_35.scala 3928:55]
  wire  _T_772 = read_stack7_pop == pop_ray_id & pop_valid; // @[lut_35.scala 3968:55]
  wire  _T_775 = read_stack8_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4008:55]
  wire  _T_778 = read_stack9_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4049:55]
  wire  _T_781 = read_stack10_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4089:56]
  wire  _T_784 = read_stack11_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4129:56]
  wire  _T_787 = read_stack12_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4169:56]
  wire  _T_790 = read_stack13_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4209:56]
  wire  _T_793 = read_stack14_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4249:56]
  wire  _T_796 = read_stack15_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4289:56]
  wire  _T_799 = read_stack16_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4329:56]
  wire  _T_802 = read_stack17_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4369:56]
  wire  _T_805 = read_stack18_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4409:56]
  wire  _T_808 = read_stack19_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4449:56]
  wire  _T_811 = read_stack20_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4489:56]
  wire  _T_814 = read_stack21_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4529:56]
  wire  _T_817 = read_stack22_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4569:56]
  wire  _T_820 = read_stack23_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4609:56]
  wire  _T_823 = read_stack24_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4649:56]
  wire  _T_826 = read_stack25_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4689:56]
  wire  _T_829 = read_stack26_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4729:56]
  wire  _T_832 = read_stack27_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4769:56]
  wire  _T_835 = read_stack28_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4809:56]
  wire  _T_838 = read_stack29_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4849:56]
  wire  _T_841 = read_stack30_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4889:56]
  wire  _T_844 = read_stack31_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4929:56]
  wire  _T_847 = read_stack32_pop == pop_ray_id & pop_valid; // @[lut_35.scala 4969:56]
  wire  _T_850 = read_stack33_pop == pop_ray_id & pop_valid; // @[lut_35.scala 5009:56]
  wire  _T_853 = read_stack34_pop == pop_ray_id & pop_valid; // @[lut_35.scala 5049:56]
  wire [31:0] _GEN_19572 = read_stack34_pop == pop_ray_id & pop_valid ? pop_ray_id : pop_ray_id_2; // @[lut_35.scala 5049:78 lut_35.scala 5087:38 lut_35.scala 3613:47]
  wire [31:0] _GEN_19573 = read_stack34_pop == pop_ray_id & pop_valid ? pop_hitT_1 : pop_hitT_2; // @[lut_35.scala 5049:78 lut_35.scala 5088:41 lut_35.scala 3614:47]
  wire  _GEN_19576 = read_stack33_pop == pop_ray_id & pop_valid ? 1'h0 : _T_853; // @[lut_35.scala 5009:78 lut_35.scala 5044:45]
  wire  _GEN_19577 = read_stack33_pop == pop_ray_id & pop_valid | _T_853; // @[lut_35.scala 5009:78 lut_35.scala 5045:40]
  wire [31:0] _GEN_19579 = read_stack33_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_19572; // @[lut_35.scala 5009:78 lut_35.scala 5047:38]
  wire [31:0] _GEN_19580 = read_stack33_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_19573; // @[lut_35.scala 5009:78 lut_35.scala 5048:41]
  wire  _GEN_19583 = read_stack32_pop == pop_ray_id & pop_valid ? 1'h0 : _T_850; // @[lut_35.scala 4969:78 lut_35.scala 5003:45]
  wire  _GEN_19584 = read_stack32_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19576; // @[lut_35.scala 4969:78 lut_35.scala 5004:45]
  wire  _GEN_19585 = read_stack32_pop == pop_ray_id & pop_valid | _GEN_19577; // @[lut_35.scala 4969:78 lut_35.scala 5005:40]
  wire [31:0] _GEN_19587 = read_stack32_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_19579; // @[lut_35.scala 4969:78 lut_35.scala 5007:38]
  wire [31:0] _GEN_19588 = read_stack32_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_19580; // @[lut_35.scala 4969:78 lut_35.scala 5008:41]
  wire  _GEN_19591 = read_stack31_pop == pop_ray_id & pop_valid ? 1'h0 : _T_847; // @[lut_35.scala 4929:78 lut_35.scala 4962:45]
  wire  _GEN_19592 = read_stack31_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19583; // @[lut_35.scala 4929:78 lut_35.scala 4963:45]
  wire  _GEN_19593 = read_stack31_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19584; // @[lut_35.scala 4929:78 lut_35.scala 4964:45]
  wire  _GEN_19594 = read_stack31_pop == pop_ray_id & pop_valid | _GEN_19585; // @[lut_35.scala 4929:78 lut_35.scala 4965:40]
  wire [31:0] _GEN_19596 = read_stack31_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_19587; // @[lut_35.scala 4929:78 lut_35.scala 4967:38]
  wire [31:0] _GEN_19597 = read_stack31_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_19588; // @[lut_35.scala 4929:78 lut_35.scala 4968:41]
  wire  _GEN_19600 = read_stack30_pop == pop_ray_id & pop_valid ? 1'h0 : _T_844; // @[lut_35.scala 4889:78 lut_35.scala 4921:45]
  wire  _GEN_19601 = read_stack30_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19591; // @[lut_35.scala 4889:78 lut_35.scala 4922:45]
  wire  _GEN_19602 = read_stack30_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19592; // @[lut_35.scala 4889:78 lut_35.scala 4923:45]
  wire  _GEN_19603 = read_stack30_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19593; // @[lut_35.scala 4889:78 lut_35.scala 4924:45]
  wire  _GEN_19604 = read_stack30_pop == pop_ray_id & pop_valid | _GEN_19594; // @[lut_35.scala 4889:78 lut_35.scala 4925:40]
  wire [31:0] _GEN_19606 = read_stack30_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_19596; // @[lut_35.scala 4889:78 lut_35.scala 4927:38]
  wire [31:0] _GEN_19607 = read_stack30_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_19597; // @[lut_35.scala 4889:78 lut_35.scala 4928:41]
  wire  _GEN_19610 = read_stack29_pop == pop_ray_id & pop_valid ? 1'h0 : _T_841; // @[lut_35.scala 4849:78 lut_35.scala 4880:45]
  wire  _GEN_19611 = read_stack29_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19600; // @[lut_35.scala 4849:78 lut_35.scala 4881:45]
  wire  _GEN_19612 = read_stack29_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19601; // @[lut_35.scala 4849:78 lut_35.scala 4882:45]
  wire  _GEN_19613 = read_stack29_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19602; // @[lut_35.scala 4849:78 lut_35.scala 4883:45]
  wire  _GEN_19614 = read_stack29_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19603; // @[lut_35.scala 4849:78 lut_35.scala 4884:45]
  wire  _GEN_19615 = read_stack29_pop == pop_ray_id & pop_valid | _GEN_19604; // @[lut_35.scala 4849:78 lut_35.scala 4885:40]
  wire [31:0] _GEN_19617 = read_stack29_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_19606; // @[lut_35.scala 4849:78 lut_35.scala 4887:38]
  wire [31:0] _GEN_19618 = read_stack29_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_19607; // @[lut_35.scala 4849:78 lut_35.scala 4888:41]
  wire  _GEN_19621 = read_stack28_pop == pop_ray_id & pop_valid ? 1'h0 : _T_838; // @[lut_35.scala 4809:78 lut_35.scala 4839:45]
  wire  _GEN_19622 = read_stack28_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19610; // @[lut_35.scala 4809:78 lut_35.scala 4840:45]
  wire  _GEN_19623 = read_stack28_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19611; // @[lut_35.scala 4809:78 lut_35.scala 4841:45]
  wire  _GEN_19624 = read_stack28_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19612; // @[lut_35.scala 4809:78 lut_35.scala 4842:45]
  wire  _GEN_19625 = read_stack28_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19613; // @[lut_35.scala 4809:78 lut_35.scala 4843:45]
  wire  _GEN_19626 = read_stack28_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19614; // @[lut_35.scala 4809:78 lut_35.scala 4844:45]
  wire  _GEN_19627 = read_stack28_pop == pop_ray_id & pop_valid | _GEN_19615; // @[lut_35.scala 4809:78 lut_35.scala 4845:40]
  wire [31:0] _GEN_19629 = read_stack28_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_19617; // @[lut_35.scala 4809:78 lut_35.scala 4847:38]
  wire [31:0] _GEN_19630 = read_stack28_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_19618; // @[lut_35.scala 4809:78 lut_35.scala 4848:41]
  wire  _GEN_19633 = read_stack27_pop == pop_ray_id & pop_valid ? 1'h0 : _T_835; // @[lut_35.scala 4769:78 lut_35.scala 4798:45]
  wire  _GEN_19634 = read_stack27_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19621; // @[lut_35.scala 4769:78 lut_35.scala 4799:45]
  wire  _GEN_19635 = read_stack27_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19622; // @[lut_35.scala 4769:78 lut_35.scala 4800:45]
  wire  _GEN_19636 = read_stack27_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19623; // @[lut_35.scala 4769:78 lut_35.scala 4801:45]
  wire  _GEN_19637 = read_stack27_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19624; // @[lut_35.scala 4769:78 lut_35.scala 4802:45]
  wire  _GEN_19638 = read_stack27_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19625; // @[lut_35.scala 4769:78 lut_35.scala 4803:45]
  wire  _GEN_19639 = read_stack27_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19626; // @[lut_35.scala 4769:78 lut_35.scala 4804:45]
  wire  _GEN_19640 = read_stack27_pop == pop_ray_id & pop_valid | _GEN_19627; // @[lut_35.scala 4769:78 lut_35.scala 4805:40]
  wire [31:0] _GEN_19642 = read_stack27_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_19629; // @[lut_35.scala 4769:78 lut_35.scala 4807:38]
  wire [31:0] _GEN_19643 = read_stack27_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_19630; // @[lut_35.scala 4769:78 lut_35.scala 4808:41]
  wire  _GEN_19646 = read_stack26_pop == pop_ray_id & pop_valid ? 1'h0 : _T_832; // @[lut_35.scala 4729:78 lut_35.scala 4757:45]
  wire  _GEN_19647 = read_stack26_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19633; // @[lut_35.scala 4729:78 lut_35.scala 4758:45]
  wire  _GEN_19648 = read_stack26_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19634; // @[lut_35.scala 4729:78 lut_35.scala 4759:45]
  wire  _GEN_19649 = read_stack26_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19635; // @[lut_35.scala 4729:78 lut_35.scala 4760:45]
  wire  _GEN_19650 = read_stack26_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19636; // @[lut_35.scala 4729:78 lut_35.scala 4761:45]
  wire  _GEN_19651 = read_stack26_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19637; // @[lut_35.scala 4729:78 lut_35.scala 4762:45]
  wire  _GEN_19652 = read_stack26_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19638; // @[lut_35.scala 4729:78 lut_35.scala 4763:45]
  wire  _GEN_19653 = read_stack26_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19639; // @[lut_35.scala 4729:78 lut_35.scala 4764:45]
  wire  _GEN_19654 = read_stack26_pop == pop_ray_id & pop_valid | _GEN_19640; // @[lut_35.scala 4729:78 lut_35.scala 4765:40]
  wire [31:0] _GEN_19656 = read_stack26_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_19642; // @[lut_35.scala 4729:78 lut_35.scala 4767:38]
  wire [31:0] _GEN_19657 = read_stack26_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_19643; // @[lut_35.scala 4729:78 lut_35.scala 4768:41]
  wire  _GEN_19660 = read_stack25_pop == pop_ray_id & pop_valid ? 1'h0 : _T_829; // @[lut_35.scala 4689:78 lut_35.scala 4716:45]
  wire  _GEN_19661 = read_stack25_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19646; // @[lut_35.scala 4689:78 lut_35.scala 4717:45]
  wire  _GEN_19662 = read_stack25_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19647; // @[lut_35.scala 4689:78 lut_35.scala 4718:45]
  wire  _GEN_19663 = read_stack25_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19648; // @[lut_35.scala 4689:78 lut_35.scala 4719:45]
  wire  _GEN_19664 = read_stack25_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19649; // @[lut_35.scala 4689:78 lut_35.scala 4720:45]
  wire  _GEN_19665 = read_stack25_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19650; // @[lut_35.scala 4689:78 lut_35.scala 4721:45]
  wire  _GEN_19666 = read_stack25_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19651; // @[lut_35.scala 4689:78 lut_35.scala 4722:45]
  wire  _GEN_19667 = read_stack25_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19652; // @[lut_35.scala 4689:78 lut_35.scala 4723:45]
  wire  _GEN_19668 = read_stack25_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19653; // @[lut_35.scala 4689:78 lut_35.scala 4724:45]
  wire  _GEN_19669 = read_stack25_pop == pop_ray_id & pop_valid | _GEN_19654; // @[lut_35.scala 4689:78 lut_35.scala 4725:40]
  wire [31:0] _GEN_19671 = read_stack25_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_19656; // @[lut_35.scala 4689:78 lut_35.scala 4727:38]
  wire [31:0] _GEN_19672 = read_stack25_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_19657; // @[lut_35.scala 4689:78 lut_35.scala 4728:41]
  wire  _GEN_19675 = read_stack24_pop == pop_ray_id & pop_valid ? 1'h0 : _T_826; // @[lut_35.scala 4649:78 lut_35.scala 4675:45]
  wire  _GEN_19676 = read_stack24_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19660; // @[lut_35.scala 4649:78 lut_35.scala 4676:45]
  wire  _GEN_19677 = read_stack24_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19661; // @[lut_35.scala 4649:78 lut_35.scala 4677:45]
  wire  _GEN_19678 = read_stack24_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19662; // @[lut_35.scala 4649:78 lut_35.scala 4678:45]
  wire  _GEN_19679 = read_stack24_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19663; // @[lut_35.scala 4649:78 lut_35.scala 4679:45]
  wire  _GEN_19680 = read_stack24_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19664; // @[lut_35.scala 4649:78 lut_35.scala 4680:45]
  wire  _GEN_19681 = read_stack24_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19665; // @[lut_35.scala 4649:78 lut_35.scala 4681:45]
  wire  _GEN_19682 = read_stack24_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19666; // @[lut_35.scala 4649:78 lut_35.scala 4682:45]
  wire  _GEN_19683 = read_stack24_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19667; // @[lut_35.scala 4649:78 lut_35.scala 4683:45]
  wire  _GEN_19684 = read_stack24_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19668; // @[lut_35.scala 4649:78 lut_35.scala 4684:45]
  wire  _GEN_19685 = read_stack24_pop == pop_ray_id & pop_valid | _GEN_19669; // @[lut_35.scala 4649:78 lut_35.scala 4685:40]
  wire [31:0] _GEN_19687 = read_stack24_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_19671; // @[lut_35.scala 4649:78 lut_35.scala 4687:38]
  wire [31:0] _GEN_19688 = read_stack24_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_19672; // @[lut_35.scala 4649:78 lut_35.scala 4688:41]
  wire  _GEN_19691 = read_stack23_pop == pop_ray_id & pop_valid ? 1'h0 : _T_823; // @[lut_35.scala 4609:78 lut_35.scala 4634:45]
  wire  _GEN_19692 = read_stack23_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19675; // @[lut_35.scala 4609:78 lut_35.scala 4635:45]
  wire  _GEN_19693 = read_stack23_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19676; // @[lut_35.scala 4609:78 lut_35.scala 4636:45]
  wire  _GEN_19694 = read_stack23_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19677; // @[lut_35.scala 4609:78 lut_35.scala 4637:45]
  wire  _GEN_19695 = read_stack23_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19678; // @[lut_35.scala 4609:78 lut_35.scala 4638:45]
  wire  _GEN_19696 = read_stack23_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19679; // @[lut_35.scala 4609:78 lut_35.scala 4639:45]
  wire  _GEN_19697 = read_stack23_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19680; // @[lut_35.scala 4609:78 lut_35.scala 4640:45]
  wire  _GEN_19698 = read_stack23_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19681; // @[lut_35.scala 4609:78 lut_35.scala 4641:45]
  wire  _GEN_19699 = read_stack23_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19682; // @[lut_35.scala 4609:78 lut_35.scala 4642:45]
  wire  _GEN_19700 = read_stack23_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19683; // @[lut_35.scala 4609:78 lut_35.scala 4643:45]
  wire  _GEN_19701 = read_stack23_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19684; // @[lut_35.scala 4609:78 lut_35.scala 4644:45]
  wire  _GEN_19702 = read_stack23_pop == pop_ray_id & pop_valid | _GEN_19685; // @[lut_35.scala 4609:78 lut_35.scala 4645:40]
  wire [31:0] _GEN_19704 = read_stack23_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_19687; // @[lut_35.scala 4609:78 lut_35.scala 4647:38]
  wire [31:0] _GEN_19705 = read_stack23_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_19688; // @[lut_35.scala 4609:78 lut_35.scala 4648:41]
  wire  _GEN_19708 = read_stack22_pop == pop_ray_id & pop_valid ? 1'h0 : _T_820; // @[lut_35.scala 4569:78 lut_35.scala 4593:45]
  wire  _GEN_19709 = read_stack22_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19691; // @[lut_35.scala 4569:78 lut_35.scala 4594:45]
  wire  _GEN_19710 = read_stack22_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19692; // @[lut_35.scala 4569:78 lut_35.scala 4595:45]
  wire  _GEN_19711 = read_stack22_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19693; // @[lut_35.scala 4569:78 lut_35.scala 4596:45]
  wire  _GEN_19712 = read_stack22_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19694; // @[lut_35.scala 4569:78 lut_35.scala 4597:45]
  wire  _GEN_19713 = read_stack22_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19695; // @[lut_35.scala 4569:78 lut_35.scala 4598:45]
  wire  _GEN_19714 = read_stack22_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19696; // @[lut_35.scala 4569:78 lut_35.scala 4599:45]
  wire  _GEN_19715 = read_stack22_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19697; // @[lut_35.scala 4569:78 lut_35.scala 4600:45]
  wire  _GEN_19716 = read_stack22_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19698; // @[lut_35.scala 4569:78 lut_35.scala 4601:45]
  wire  _GEN_19717 = read_stack22_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19699; // @[lut_35.scala 4569:78 lut_35.scala 4602:45]
  wire  _GEN_19718 = read_stack22_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19700; // @[lut_35.scala 4569:78 lut_35.scala 4603:45]
  wire  _GEN_19719 = read_stack22_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19701; // @[lut_35.scala 4569:78 lut_35.scala 4604:45]
  wire  _GEN_19720 = read_stack22_pop == pop_ray_id & pop_valid | _GEN_19702; // @[lut_35.scala 4569:78 lut_35.scala 4605:40]
  wire [31:0] _GEN_19722 = read_stack22_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_19704; // @[lut_35.scala 4569:78 lut_35.scala 4607:38]
  wire [31:0] _GEN_19723 = read_stack22_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_19705; // @[lut_35.scala 4569:78 lut_35.scala 4608:41]
  wire  _GEN_19726 = read_stack21_pop == pop_ray_id & pop_valid ? 1'h0 : _T_817; // @[lut_35.scala 4529:78 lut_35.scala 4552:45]
  wire  _GEN_19727 = read_stack21_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19708; // @[lut_35.scala 4529:78 lut_35.scala 4553:45]
  wire  _GEN_19728 = read_stack21_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19709; // @[lut_35.scala 4529:78 lut_35.scala 4554:45]
  wire  _GEN_19729 = read_stack21_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19710; // @[lut_35.scala 4529:78 lut_35.scala 4555:45]
  wire  _GEN_19730 = read_stack21_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19711; // @[lut_35.scala 4529:78 lut_35.scala 4556:45]
  wire  _GEN_19731 = read_stack21_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19712; // @[lut_35.scala 4529:78 lut_35.scala 4557:45]
  wire  _GEN_19732 = read_stack21_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19713; // @[lut_35.scala 4529:78 lut_35.scala 4558:45]
  wire  _GEN_19733 = read_stack21_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19714; // @[lut_35.scala 4529:78 lut_35.scala 4559:45]
  wire  _GEN_19734 = read_stack21_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19715; // @[lut_35.scala 4529:78 lut_35.scala 4560:45]
  wire  _GEN_19735 = read_stack21_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19716; // @[lut_35.scala 4529:78 lut_35.scala 4561:45]
  wire  _GEN_19736 = read_stack21_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19717; // @[lut_35.scala 4529:78 lut_35.scala 4562:45]
  wire  _GEN_19737 = read_stack21_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19718; // @[lut_35.scala 4529:78 lut_35.scala 4563:45]
  wire  _GEN_19738 = read_stack21_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19719; // @[lut_35.scala 4529:78 lut_35.scala 4564:45]
  wire  _GEN_19739 = read_stack21_pop == pop_ray_id & pop_valid | _GEN_19720; // @[lut_35.scala 4529:78 lut_35.scala 4565:40]
  wire [31:0] _GEN_19741 = read_stack21_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_19722; // @[lut_35.scala 4529:78 lut_35.scala 4567:38]
  wire [31:0] _GEN_19742 = read_stack21_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_19723; // @[lut_35.scala 4529:78 lut_35.scala 4568:41]
  wire  _GEN_19745 = read_stack20_pop == pop_ray_id & pop_valid ? 1'h0 : _T_814; // @[lut_35.scala 4489:78 lut_35.scala 4511:45]
  wire  _GEN_19746 = read_stack20_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19726; // @[lut_35.scala 4489:78 lut_35.scala 4512:45]
  wire  _GEN_19747 = read_stack20_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19727; // @[lut_35.scala 4489:78 lut_35.scala 4513:45]
  wire  _GEN_19748 = read_stack20_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19728; // @[lut_35.scala 4489:78 lut_35.scala 4514:45]
  wire  _GEN_19749 = read_stack20_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19729; // @[lut_35.scala 4489:78 lut_35.scala 4515:45]
  wire  _GEN_19750 = read_stack20_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19730; // @[lut_35.scala 4489:78 lut_35.scala 4516:45]
  wire  _GEN_19751 = read_stack20_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19731; // @[lut_35.scala 4489:78 lut_35.scala 4517:45]
  wire  _GEN_19752 = read_stack20_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19732; // @[lut_35.scala 4489:78 lut_35.scala 4518:45]
  wire  _GEN_19753 = read_stack20_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19733; // @[lut_35.scala 4489:78 lut_35.scala 4519:45]
  wire  _GEN_19754 = read_stack20_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19734; // @[lut_35.scala 4489:78 lut_35.scala 4520:45]
  wire  _GEN_19755 = read_stack20_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19735; // @[lut_35.scala 4489:78 lut_35.scala 4521:45]
  wire  _GEN_19756 = read_stack20_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19736; // @[lut_35.scala 4489:78 lut_35.scala 4522:45]
  wire  _GEN_19757 = read_stack20_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19737; // @[lut_35.scala 4489:78 lut_35.scala 4523:45]
  wire  _GEN_19758 = read_stack20_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19738; // @[lut_35.scala 4489:78 lut_35.scala 4524:45]
  wire  _GEN_19759 = read_stack20_pop == pop_ray_id & pop_valid | _GEN_19739; // @[lut_35.scala 4489:78 lut_35.scala 4525:40]
  wire [31:0] _GEN_19761 = read_stack20_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_19741; // @[lut_35.scala 4489:78 lut_35.scala 4527:38]
  wire [31:0] _GEN_19762 = read_stack20_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_19742; // @[lut_35.scala 4489:78 lut_35.scala 4528:41]
  wire  _GEN_19765 = read_stack19_pop == pop_ray_id & pop_valid ? 1'h0 : _T_811; // @[lut_35.scala 4449:78 lut_35.scala 4470:45]
  wire  _GEN_19766 = read_stack19_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19745; // @[lut_35.scala 4449:78 lut_35.scala 4471:45]
  wire  _GEN_19767 = read_stack19_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19746; // @[lut_35.scala 4449:78 lut_35.scala 4472:45]
  wire  _GEN_19768 = read_stack19_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19747; // @[lut_35.scala 4449:78 lut_35.scala 4473:45]
  wire  _GEN_19769 = read_stack19_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19748; // @[lut_35.scala 4449:78 lut_35.scala 4474:45]
  wire  _GEN_19770 = read_stack19_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19749; // @[lut_35.scala 4449:78 lut_35.scala 4475:45]
  wire  _GEN_19771 = read_stack19_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19750; // @[lut_35.scala 4449:78 lut_35.scala 4476:45]
  wire  _GEN_19772 = read_stack19_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19751; // @[lut_35.scala 4449:78 lut_35.scala 4477:45]
  wire  _GEN_19773 = read_stack19_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19752; // @[lut_35.scala 4449:78 lut_35.scala 4478:45]
  wire  _GEN_19774 = read_stack19_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19753; // @[lut_35.scala 4449:78 lut_35.scala 4479:45]
  wire  _GEN_19775 = read_stack19_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19754; // @[lut_35.scala 4449:78 lut_35.scala 4480:45]
  wire  _GEN_19776 = read_stack19_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19755; // @[lut_35.scala 4449:78 lut_35.scala 4481:45]
  wire  _GEN_19777 = read_stack19_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19756; // @[lut_35.scala 4449:78 lut_35.scala 4482:45]
  wire  _GEN_19778 = read_stack19_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19757; // @[lut_35.scala 4449:78 lut_35.scala 4483:45]
  wire  _GEN_19779 = read_stack19_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19758; // @[lut_35.scala 4449:78 lut_35.scala 4484:45]
  wire  _GEN_19780 = read_stack19_pop == pop_ray_id & pop_valid | _GEN_19759; // @[lut_35.scala 4449:78 lut_35.scala 4485:40]
  wire [31:0] _GEN_19782 = read_stack19_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_19761; // @[lut_35.scala 4449:78 lut_35.scala 4487:38]
  wire [31:0] _GEN_19783 = read_stack19_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_19762; // @[lut_35.scala 4449:78 lut_35.scala 4488:41]
  wire  _GEN_19786 = read_stack18_pop == pop_ray_id & pop_valid ? 1'h0 : _T_808; // @[lut_35.scala 4409:78 lut_35.scala 4429:45]
  wire  _GEN_19787 = read_stack18_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19765; // @[lut_35.scala 4409:78 lut_35.scala 4430:45]
  wire  _GEN_19788 = read_stack18_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19766; // @[lut_35.scala 4409:78 lut_35.scala 4431:45]
  wire  _GEN_19789 = read_stack18_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19767; // @[lut_35.scala 4409:78 lut_35.scala 4432:45]
  wire  _GEN_19790 = read_stack18_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19768; // @[lut_35.scala 4409:78 lut_35.scala 4433:45]
  wire  _GEN_19791 = read_stack18_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19769; // @[lut_35.scala 4409:78 lut_35.scala 4434:45]
  wire  _GEN_19792 = read_stack18_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19770; // @[lut_35.scala 4409:78 lut_35.scala 4435:45]
  wire  _GEN_19793 = read_stack18_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19771; // @[lut_35.scala 4409:78 lut_35.scala 4436:45]
  wire  _GEN_19794 = read_stack18_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19772; // @[lut_35.scala 4409:78 lut_35.scala 4437:45]
  wire  _GEN_19795 = read_stack18_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19773; // @[lut_35.scala 4409:78 lut_35.scala 4438:45]
  wire  _GEN_19796 = read_stack18_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19774; // @[lut_35.scala 4409:78 lut_35.scala 4439:45]
  wire  _GEN_19797 = read_stack18_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19775; // @[lut_35.scala 4409:78 lut_35.scala 4440:45]
  wire  _GEN_19798 = read_stack18_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19776; // @[lut_35.scala 4409:78 lut_35.scala 4441:45]
  wire  _GEN_19799 = read_stack18_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19777; // @[lut_35.scala 4409:78 lut_35.scala 4442:45]
  wire  _GEN_19800 = read_stack18_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19778; // @[lut_35.scala 4409:78 lut_35.scala 4443:45]
  wire  _GEN_19801 = read_stack18_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19779; // @[lut_35.scala 4409:78 lut_35.scala 4444:45]
  wire  _GEN_19802 = read_stack18_pop == pop_ray_id & pop_valid | _GEN_19780; // @[lut_35.scala 4409:78 lut_35.scala 4445:40]
  wire [31:0] _GEN_19804 = read_stack18_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_19782; // @[lut_35.scala 4409:78 lut_35.scala 4447:38]
  wire [31:0] _GEN_19805 = read_stack18_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_19783; // @[lut_35.scala 4409:78 lut_35.scala 4448:41]
  wire  _GEN_19808 = read_stack17_pop == pop_ray_id & pop_valid ? 1'h0 : _T_805; // @[lut_35.scala 4369:78 lut_35.scala 4388:45]
  wire  _GEN_19809 = read_stack17_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19786; // @[lut_35.scala 4369:78 lut_35.scala 4389:45]
  wire  _GEN_19810 = read_stack17_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19787; // @[lut_35.scala 4369:78 lut_35.scala 4390:45]
  wire  _GEN_19811 = read_stack17_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19788; // @[lut_35.scala 4369:78 lut_35.scala 4391:45]
  wire  _GEN_19812 = read_stack17_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19789; // @[lut_35.scala 4369:78 lut_35.scala 4392:45]
  wire  _GEN_19813 = read_stack17_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19790; // @[lut_35.scala 4369:78 lut_35.scala 4393:45]
  wire  _GEN_19814 = read_stack17_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19791; // @[lut_35.scala 4369:78 lut_35.scala 4394:45]
  wire  _GEN_19815 = read_stack17_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19792; // @[lut_35.scala 4369:78 lut_35.scala 4395:45]
  wire  _GEN_19816 = read_stack17_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19793; // @[lut_35.scala 4369:78 lut_35.scala 4396:45]
  wire  _GEN_19817 = read_stack17_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19794; // @[lut_35.scala 4369:78 lut_35.scala 4397:45]
  wire  _GEN_19818 = read_stack17_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19795; // @[lut_35.scala 4369:78 lut_35.scala 4398:45]
  wire  _GEN_19819 = read_stack17_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19796; // @[lut_35.scala 4369:78 lut_35.scala 4399:45]
  wire  _GEN_19820 = read_stack17_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19797; // @[lut_35.scala 4369:78 lut_35.scala 4400:45]
  wire  _GEN_19821 = read_stack17_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19798; // @[lut_35.scala 4369:78 lut_35.scala 4401:45]
  wire  _GEN_19822 = read_stack17_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19799; // @[lut_35.scala 4369:78 lut_35.scala 4402:45]
  wire  _GEN_19823 = read_stack17_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19800; // @[lut_35.scala 4369:78 lut_35.scala 4403:45]
  wire  _GEN_19824 = read_stack17_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19801; // @[lut_35.scala 4369:78 lut_35.scala 4404:45]
  wire  _GEN_19825 = read_stack17_pop == pop_ray_id & pop_valid | _GEN_19802; // @[lut_35.scala 4369:78 lut_35.scala 4405:40]
  wire [31:0] _GEN_19827 = read_stack17_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_19804; // @[lut_35.scala 4369:78 lut_35.scala 4407:38]
  wire [31:0] _GEN_19828 = read_stack17_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_19805; // @[lut_35.scala 4369:78 lut_35.scala 4408:41]
  wire  _GEN_19831 = read_stack16_pop == pop_ray_id & pop_valid ? 1'h0 : _T_802; // @[lut_35.scala 4329:78 lut_35.scala 4347:45]
  wire  _GEN_19832 = read_stack16_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19808; // @[lut_35.scala 4329:78 lut_35.scala 4348:45]
  wire  _GEN_19833 = read_stack16_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19809; // @[lut_35.scala 4329:78 lut_35.scala 4349:45]
  wire  _GEN_19834 = read_stack16_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19810; // @[lut_35.scala 4329:78 lut_35.scala 4350:45]
  wire  _GEN_19835 = read_stack16_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19811; // @[lut_35.scala 4329:78 lut_35.scala 4351:45]
  wire  _GEN_19836 = read_stack16_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19812; // @[lut_35.scala 4329:78 lut_35.scala 4352:45]
  wire  _GEN_19837 = read_stack16_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19813; // @[lut_35.scala 4329:78 lut_35.scala 4353:45]
  wire  _GEN_19838 = read_stack16_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19814; // @[lut_35.scala 4329:78 lut_35.scala 4354:45]
  wire  _GEN_19839 = read_stack16_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19815; // @[lut_35.scala 4329:78 lut_35.scala 4355:45]
  wire  _GEN_19840 = read_stack16_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19816; // @[lut_35.scala 4329:78 lut_35.scala 4356:45]
  wire  _GEN_19841 = read_stack16_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19817; // @[lut_35.scala 4329:78 lut_35.scala 4357:45]
  wire  _GEN_19842 = read_stack16_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19818; // @[lut_35.scala 4329:78 lut_35.scala 4358:45]
  wire  _GEN_19843 = read_stack16_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19819; // @[lut_35.scala 4329:78 lut_35.scala 4359:45]
  wire  _GEN_19844 = read_stack16_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19820; // @[lut_35.scala 4329:78 lut_35.scala 4360:45]
  wire  _GEN_19845 = read_stack16_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19821; // @[lut_35.scala 4329:78 lut_35.scala 4361:45]
  wire  _GEN_19846 = read_stack16_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19822; // @[lut_35.scala 4329:78 lut_35.scala 4362:45]
  wire  _GEN_19847 = read_stack16_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19823; // @[lut_35.scala 4329:78 lut_35.scala 4363:45]
  wire  _GEN_19848 = read_stack16_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19824; // @[lut_35.scala 4329:78 lut_35.scala 4364:45]
  wire  _GEN_19849 = read_stack16_pop == pop_ray_id & pop_valid | _GEN_19825; // @[lut_35.scala 4329:78 lut_35.scala 4365:40]
  wire [31:0] _GEN_19851 = read_stack16_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_19827; // @[lut_35.scala 4329:78 lut_35.scala 4367:38]
  wire [31:0] _GEN_19852 = read_stack16_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_19828; // @[lut_35.scala 4329:78 lut_35.scala 4368:41]
  wire  _GEN_19855 = read_stack15_pop == pop_ray_id & pop_valid ? 1'h0 : _T_799; // @[lut_35.scala 4289:78 lut_35.scala 4306:45]
  wire  _GEN_19856 = read_stack15_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19831; // @[lut_35.scala 4289:78 lut_35.scala 4307:45]
  wire  _GEN_19857 = read_stack15_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19832; // @[lut_35.scala 4289:78 lut_35.scala 4308:45]
  wire  _GEN_19858 = read_stack15_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19833; // @[lut_35.scala 4289:78 lut_35.scala 4309:45]
  wire  _GEN_19859 = read_stack15_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19834; // @[lut_35.scala 4289:78 lut_35.scala 4310:45]
  wire  _GEN_19860 = read_stack15_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19835; // @[lut_35.scala 4289:78 lut_35.scala 4311:45]
  wire  _GEN_19861 = read_stack15_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19836; // @[lut_35.scala 4289:78 lut_35.scala 4312:45]
  wire  _GEN_19862 = read_stack15_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19837; // @[lut_35.scala 4289:78 lut_35.scala 4313:45]
  wire  _GEN_19863 = read_stack15_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19838; // @[lut_35.scala 4289:78 lut_35.scala 4314:45]
  wire  _GEN_19864 = read_stack15_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19839; // @[lut_35.scala 4289:78 lut_35.scala 4315:45]
  wire  _GEN_19865 = read_stack15_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19840; // @[lut_35.scala 4289:78 lut_35.scala 4316:45]
  wire  _GEN_19866 = read_stack15_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19841; // @[lut_35.scala 4289:78 lut_35.scala 4317:45]
  wire  _GEN_19867 = read_stack15_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19842; // @[lut_35.scala 4289:78 lut_35.scala 4318:45]
  wire  _GEN_19868 = read_stack15_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19843; // @[lut_35.scala 4289:78 lut_35.scala 4319:45]
  wire  _GEN_19869 = read_stack15_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19844; // @[lut_35.scala 4289:78 lut_35.scala 4320:45]
  wire  _GEN_19870 = read_stack15_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19845; // @[lut_35.scala 4289:78 lut_35.scala 4321:45]
  wire  _GEN_19871 = read_stack15_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19846; // @[lut_35.scala 4289:78 lut_35.scala 4322:45]
  wire  _GEN_19872 = read_stack15_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19847; // @[lut_35.scala 4289:78 lut_35.scala 4323:45]
  wire  _GEN_19873 = read_stack15_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19848; // @[lut_35.scala 4289:78 lut_35.scala 4324:45]
  wire  _GEN_19874 = read_stack15_pop == pop_ray_id & pop_valid | _GEN_19849; // @[lut_35.scala 4289:78 lut_35.scala 4325:40]
  wire [31:0] _GEN_19876 = read_stack15_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_19851; // @[lut_35.scala 4289:78 lut_35.scala 4327:38]
  wire [31:0] _GEN_19877 = read_stack15_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_19852; // @[lut_35.scala 4289:78 lut_35.scala 4328:41]
  wire  _GEN_19880 = read_stack14_pop == pop_ray_id & pop_valid ? 1'h0 : _T_796; // @[lut_35.scala 4249:78 lut_35.scala 4265:45]
  wire  _GEN_19881 = read_stack14_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19855; // @[lut_35.scala 4249:78 lut_35.scala 4266:45]
  wire  _GEN_19882 = read_stack14_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19856; // @[lut_35.scala 4249:78 lut_35.scala 4267:45]
  wire  _GEN_19883 = read_stack14_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19857; // @[lut_35.scala 4249:78 lut_35.scala 4268:45]
  wire  _GEN_19884 = read_stack14_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19858; // @[lut_35.scala 4249:78 lut_35.scala 4269:45]
  wire  _GEN_19885 = read_stack14_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19859; // @[lut_35.scala 4249:78 lut_35.scala 4270:45]
  wire  _GEN_19886 = read_stack14_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19860; // @[lut_35.scala 4249:78 lut_35.scala 4271:45]
  wire  _GEN_19887 = read_stack14_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19861; // @[lut_35.scala 4249:78 lut_35.scala 4272:45]
  wire  _GEN_19888 = read_stack14_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19862; // @[lut_35.scala 4249:78 lut_35.scala 4273:45]
  wire  _GEN_19889 = read_stack14_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19863; // @[lut_35.scala 4249:78 lut_35.scala 4274:45]
  wire  _GEN_19890 = read_stack14_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19864; // @[lut_35.scala 4249:78 lut_35.scala 4275:45]
  wire  _GEN_19891 = read_stack14_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19865; // @[lut_35.scala 4249:78 lut_35.scala 4276:45]
  wire  _GEN_19892 = read_stack14_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19866; // @[lut_35.scala 4249:78 lut_35.scala 4277:45]
  wire  _GEN_19893 = read_stack14_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19867; // @[lut_35.scala 4249:78 lut_35.scala 4278:45]
  wire  _GEN_19894 = read_stack14_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19868; // @[lut_35.scala 4249:78 lut_35.scala 4279:45]
  wire  _GEN_19895 = read_stack14_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19869; // @[lut_35.scala 4249:78 lut_35.scala 4280:45]
  wire  _GEN_19896 = read_stack14_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19870; // @[lut_35.scala 4249:78 lut_35.scala 4281:45]
  wire  _GEN_19897 = read_stack14_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19871; // @[lut_35.scala 4249:78 lut_35.scala 4282:45]
  wire  _GEN_19898 = read_stack14_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19872; // @[lut_35.scala 4249:78 lut_35.scala 4283:45]
  wire  _GEN_19899 = read_stack14_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19873; // @[lut_35.scala 4249:78 lut_35.scala 4284:45]
  wire  _GEN_19900 = read_stack14_pop == pop_ray_id & pop_valid | _GEN_19874; // @[lut_35.scala 4249:78 lut_35.scala 4285:40]
  wire [31:0] _GEN_19902 = read_stack14_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_19876; // @[lut_35.scala 4249:78 lut_35.scala 4287:38]
  wire [31:0] _GEN_19903 = read_stack14_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_19877; // @[lut_35.scala 4249:78 lut_35.scala 4288:41]
  wire  _GEN_19906 = read_stack13_pop == pop_ray_id & pop_valid ? 1'h0 : _T_793; // @[lut_35.scala 4209:78 lut_35.scala 4224:45]
  wire  _GEN_19907 = read_stack13_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19880; // @[lut_35.scala 4209:78 lut_35.scala 4225:45]
  wire  _GEN_19908 = read_stack13_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19881; // @[lut_35.scala 4209:78 lut_35.scala 4226:45]
  wire  _GEN_19909 = read_stack13_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19882; // @[lut_35.scala 4209:78 lut_35.scala 4227:45]
  wire  _GEN_19910 = read_stack13_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19883; // @[lut_35.scala 4209:78 lut_35.scala 4228:45]
  wire  _GEN_19911 = read_stack13_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19884; // @[lut_35.scala 4209:78 lut_35.scala 4229:45]
  wire  _GEN_19912 = read_stack13_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19885; // @[lut_35.scala 4209:78 lut_35.scala 4230:45]
  wire  _GEN_19913 = read_stack13_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19886; // @[lut_35.scala 4209:78 lut_35.scala 4231:45]
  wire  _GEN_19914 = read_stack13_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19887; // @[lut_35.scala 4209:78 lut_35.scala 4232:45]
  wire  _GEN_19915 = read_stack13_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19888; // @[lut_35.scala 4209:78 lut_35.scala 4233:45]
  wire  _GEN_19916 = read_stack13_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19889; // @[lut_35.scala 4209:78 lut_35.scala 4234:45]
  wire  _GEN_19917 = read_stack13_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19890; // @[lut_35.scala 4209:78 lut_35.scala 4235:45]
  wire  _GEN_19918 = read_stack13_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19891; // @[lut_35.scala 4209:78 lut_35.scala 4236:45]
  wire  _GEN_19919 = read_stack13_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19892; // @[lut_35.scala 4209:78 lut_35.scala 4237:45]
  wire  _GEN_19920 = read_stack13_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19893; // @[lut_35.scala 4209:78 lut_35.scala 4238:45]
  wire  _GEN_19921 = read_stack13_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19894; // @[lut_35.scala 4209:78 lut_35.scala 4239:45]
  wire  _GEN_19922 = read_stack13_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19895; // @[lut_35.scala 4209:78 lut_35.scala 4240:45]
  wire  _GEN_19923 = read_stack13_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19896; // @[lut_35.scala 4209:78 lut_35.scala 4241:45]
  wire  _GEN_19924 = read_stack13_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19897; // @[lut_35.scala 4209:78 lut_35.scala 4242:45]
  wire  _GEN_19925 = read_stack13_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19898; // @[lut_35.scala 4209:78 lut_35.scala 4243:45]
  wire  _GEN_19926 = read_stack13_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19899; // @[lut_35.scala 4209:78 lut_35.scala 4244:45]
  wire  _GEN_19927 = read_stack13_pop == pop_ray_id & pop_valid | _GEN_19900; // @[lut_35.scala 4209:78 lut_35.scala 4245:40]
  wire [31:0] _GEN_19929 = read_stack13_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_19902; // @[lut_35.scala 4209:78 lut_35.scala 4247:38]
  wire [31:0] _GEN_19930 = read_stack13_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_19903; // @[lut_35.scala 4209:78 lut_35.scala 4248:41]
  wire  _GEN_19933 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _T_790; // @[lut_35.scala 4169:78 lut_35.scala 4183:45]
  wire  _GEN_19934 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19906; // @[lut_35.scala 4169:78 lut_35.scala 4184:45]
  wire  _GEN_19935 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19907; // @[lut_35.scala 4169:78 lut_35.scala 4185:45]
  wire  _GEN_19936 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19908; // @[lut_35.scala 4169:78 lut_35.scala 4186:45]
  wire  _GEN_19937 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19909; // @[lut_35.scala 4169:78 lut_35.scala 4187:45]
  wire  _GEN_19938 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19910; // @[lut_35.scala 4169:78 lut_35.scala 4188:45]
  wire  _GEN_19939 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19911; // @[lut_35.scala 4169:78 lut_35.scala 4189:45]
  wire  _GEN_19940 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19912; // @[lut_35.scala 4169:78 lut_35.scala 4190:45]
  wire  _GEN_19941 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19913; // @[lut_35.scala 4169:78 lut_35.scala 4191:45]
  wire  _GEN_19942 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19914; // @[lut_35.scala 4169:78 lut_35.scala 4192:45]
  wire  _GEN_19943 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19915; // @[lut_35.scala 4169:78 lut_35.scala 4193:45]
  wire  _GEN_19944 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19916; // @[lut_35.scala 4169:78 lut_35.scala 4194:45]
  wire  _GEN_19945 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19917; // @[lut_35.scala 4169:78 lut_35.scala 4195:45]
  wire  _GEN_19946 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19918; // @[lut_35.scala 4169:78 lut_35.scala 4196:45]
  wire  _GEN_19947 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19919; // @[lut_35.scala 4169:78 lut_35.scala 4197:45]
  wire  _GEN_19948 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19920; // @[lut_35.scala 4169:78 lut_35.scala 4198:45]
  wire  _GEN_19949 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19921; // @[lut_35.scala 4169:78 lut_35.scala 4199:45]
  wire  _GEN_19950 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19922; // @[lut_35.scala 4169:78 lut_35.scala 4200:45]
  wire  _GEN_19951 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19923; // @[lut_35.scala 4169:78 lut_35.scala 4201:45]
  wire  _GEN_19952 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19924; // @[lut_35.scala 4169:78 lut_35.scala 4202:45]
  wire  _GEN_19953 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19925; // @[lut_35.scala 4169:78 lut_35.scala 4203:45]
  wire  _GEN_19954 = read_stack12_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19926; // @[lut_35.scala 4169:78 lut_35.scala 4204:45]
  wire  _GEN_19955 = read_stack12_pop == pop_ray_id & pop_valid | _GEN_19927; // @[lut_35.scala 4169:78 lut_35.scala 4205:40]
  wire [31:0] _GEN_19957 = read_stack12_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_19929; // @[lut_35.scala 4169:78 lut_35.scala 4207:38]
  wire [31:0] _GEN_19958 = read_stack12_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_19930; // @[lut_35.scala 4169:78 lut_35.scala 4208:41]
  wire  _GEN_19961 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _T_787; // @[lut_35.scala 4129:78 lut_35.scala 4142:45]
  wire  _GEN_19962 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19933; // @[lut_35.scala 4129:78 lut_35.scala 4143:45]
  wire  _GEN_19963 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19934; // @[lut_35.scala 4129:78 lut_35.scala 4144:45]
  wire  _GEN_19964 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19935; // @[lut_35.scala 4129:78 lut_35.scala 4145:45]
  wire  _GEN_19965 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19936; // @[lut_35.scala 4129:78 lut_35.scala 4146:45]
  wire  _GEN_19966 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19937; // @[lut_35.scala 4129:78 lut_35.scala 4147:45]
  wire  _GEN_19967 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19938; // @[lut_35.scala 4129:78 lut_35.scala 4148:45]
  wire  _GEN_19968 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19939; // @[lut_35.scala 4129:78 lut_35.scala 4149:45]
  wire  _GEN_19969 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19940; // @[lut_35.scala 4129:78 lut_35.scala 4150:45]
  wire  _GEN_19970 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19941; // @[lut_35.scala 4129:78 lut_35.scala 4151:45]
  wire  _GEN_19971 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19942; // @[lut_35.scala 4129:78 lut_35.scala 4152:45]
  wire  _GEN_19972 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19943; // @[lut_35.scala 4129:78 lut_35.scala 4153:45]
  wire  _GEN_19973 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19944; // @[lut_35.scala 4129:78 lut_35.scala 4154:45]
  wire  _GEN_19974 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19945; // @[lut_35.scala 4129:78 lut_35.scala 4155:45]
  wire  _GEN_19975 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19946; // @[lut_35.scala 4129:78 lut_35.scala 4156:45]
  wire  _GEN_19976 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19947; // @[lut_35.scala 4129:78 lut_35.scala 4157:45]
  wire  _GEN_19977 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19948; // @[lut_35.scala 4129:78 lut_35.scala 4158:45]
  wire  _GEN_19978 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19949; // @[lut_35.scala 4129:78 lut_35.scala 4159:45]
  wire  _GEN_19979 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19950; // @[lut_35.scala 4129:78 lut_35.scala 4160:45]
  wire  _GEN_19980 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19951; // @[lut_35.scala 4129:78 lut_35.scala 4161:45]
  wire  _GEN_19981 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19952; // @[lut_35.scala 4129:78 lut_35.scala 4162:45]
  wire  _GEN_19982 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19953; // @[lut_35.scala 4129:78 lut_35.scala 4163:45]
  wire  _GEN_19983 = read_stack11_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19954; // @[lut_35.scala 4129:78 lut_35.scala 4164:45]
  wire  _GEN_19984 = read_stack11_pop == pop_ray_id & pop_valid | _GEN_19955; // @[lut_35.scala 4129:78 lut_35.scala 4165:40]
  wire [31:0] _GEN_19986 = read_stack11_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_19957; // @[lut_35.scala 4129:78 lut_35.scala 4167:38]
  wire [31:0] _GEN_19987 = read_stack11_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_19958; // @[lut_35.scala 4129:78 lut_35.scala 4168:41]
  wire  _GEN_19990 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _T_784; // @[lut_35.scala 4089:78 lut_35.scala 4101:45]
  wire  _GEN_19991 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19961; // @[lut_35.scala 4089:78 lut_35.scala 4102:45]
  wire  _GEN_19992 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19962; // @[lut_35.scala 4089:78 lut_35.scala 4103:45]
  wire  _GEN_19993 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19963; // @[lut_35.scala 4089:78 lut_35.scala 4104:45]
  wire  _GEN_19994 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19964; // @[lut_35.scala 4089:78 lut_35.scala 4105:45]
  wire  _GEN_19995 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19965; // @[lut_35.scala 4089:78 lut_35.scala 4106:45]
  wire  _GEN_19996 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19966; // @[lut_35.scala 4089:78 lut_35.scala 4107:45]
  wire  _GEN_19997 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19967; // @[lut_35.scala 4089:78 lut_35.scala 4108:45]
  wire  _GEN_19998 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19968; // @[lut_35.scala 4089:78 lut_35.scala 4109:45]
  wire  _GEN_19999 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19969; // @[lut_35.scala 4089:78 lut_35.scala 4110:45]
  wire  _GEN_20000 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19970; // @[lut_35.scala 4089:78 lut_35.scala 4111:45]
  wire  _GEN_20001 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19971; // @[lut_35.scala 4089:78 lut_35.scala 4112:45]
  wire  _GEN_20002 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19972; // @[lut_35.scala 4089:78 lut_35.scala 4113:45]
  wire  _GEN_20003 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19973; // @[lut_35.scala 4089:78 lut_35.scala 4114:45]
  wire  _GEN_20004 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19974; // @[lut_35.scala 4089:78 lut_35.scala 4115:45]
  wire  _GEN_20005 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19975; // @[lut_35.scala 4089:78 lut_35.scala 4116:45]
  wire  _GEN_20006 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19976; // @[lut_35.scala 4089:78 lut_35.scala 4117:45]
  wire  _GEN_20007 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19977; // @[lut_35.scala 4089:78 lut_35.scala 4118:45]
  wire  _GEN_20008 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19978; // @[lut_35.scala 4089:78 lut_35.scala 4119:45]
  wire  _GEN_20009 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19979; // @[lut_35.scala 4089:78 lut_35.scala 4120:45]
  wire  _GEN_20010 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19980; // @[lut_35.scala 4089:78 lut_35.scala 4121:45]
  wire  _GEN_20011 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19981; // @[lut_35.scala 4089:78 lut_35.scala 4122:45]
  wire  _GEN_20012 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19982; // @[lut_35.scala 4089:78 lut_35.scala 4123:45]
  wire  _GEN_20013 = read_stack10_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19983; // @[lut_35.scala 4089:78 lut_35.scala 4124:45]
  wire  _GEN_20014 = read_stack10_pop == pop_ray_id & pop_valid | _GEN_19984; // @[lut_35.scala 4089:78 lut_35.scala 4125:40]
  wire [31:0] _GEN_20016 = read_stack10_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_19986; // @[lut_35.scala 4089:78 lut_35.scala 4127:38]
  wire [31:0] _GEN_20017 = read_stack10_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_19987; // @[lut_35.scala 4089:78 lut_35.scala 4128:41]
  wire  _GEN_20020 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _T_781; // @[lut_35.scala 4049:77 lut_35.scala 4060:45]
  wire  _GEN_20021 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19990; // @[lut_35.scala 4049:77 lut_35.scala 4061:45]
  wire  _GEN_20022 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19991; // @[lut_35.scala 4049:77 lut_35.scala 4062:45]
  wire  _GEN_20023 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19992; // @[lut_35.scala 4049:77 lut_35.scala 4063:45]
  wire  _GEN_20024 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19993; // @[lut_35.scala 4049:77 lut_35.scala 4064:45]
  wire  _GEN_20025 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19994; // @[lut_35.scala 4049:77 lut_35.scala 4065:45]
  wire  _GEN_20026 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19995; // @[lut_35.scala 4049:77 lut_35.scala 4066:45]
  wire  _GEN_20027 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19996; // @[lut_35.scala 4049:77 lut_35.scala 4067:45]
  wire  _GEN_20028 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19997; // @[lut_35.scala 4049:77 lut_35.scala 4068:45]
  wire  _GEN_20029 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19998; // @[lut_35.scala 4049:77 lut_35.scala 4069:45]
  wire  _GEN_20030 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_19999; // @[lut_35.scala 4049:77 lut_35.scala 4070:45]
  wire  _GEN_20031 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20000; // @[lut_35.scala 4049:77 lut_35.scala 4071:45]
  wire  _GEN_20032 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20001; // @[lut_35.scala 4049:77 lut_35.scala 4072:45]
  wire  _GEN_20033 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20002; // @[lut_35.scala 4049:77 lut_35.scala 4073:45]
  wire  _GEN_20034 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20003; // @[lut_35.scala 4049:77 lut_35.scala 4074:45]
  wire  _GEN_20035 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20004; // @[lut_35.scala 4049:77 lut_35.scala 4075:45]
  wire  _GEN_20036 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20005; // @[lut_35.scala 4049:77 lut_35.scala 4076:45]
  wire  _GEN_20037 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20006; // @[lut_35.scala 4049:77 lut_35.scala 4077:45]
  wire  _GEN_20038 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20007; // @[lut_35.scala 4049:77 lut_35.scala 4078:45]
  wire  _GEN_20039 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20008; // @[lut_35.scala 4049:77 lut_35.scala 4079:45]
  wire  _GEN_20040 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20009; // @[lut_35.scala 4049:77 lut_35.scala 4080:45]
  wire  _GEN_20041 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20010; // @[lut_35.scala 4049:77 lut_35.scala 4081:45]
  wire  _GEN_20042 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20011; // @[lut_35.scala 4049:77 lut_35.scala 4082:45]
  wire  _GEN_20043 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20012; // @[lut_35.scala 4049:77 lut_35.scala 4083:45]
  wire  _GEN_20044 = read_stack9_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20013; // @[lut_35.scala 4049:77 lut_35.scala 4084:45]
  wire  _GEN_20045 = read_stack9_pop == pop_ray_id & pop_valid | _GEN_20014; // @[lut_35.scala 4049:77 lut_35.scala 4085:40]
  wire [31:0] _GEN_20047 = read_stack9_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_20016; // @[lut_35.scala 4049:77 lut_35.scala 4087:38]
  wire [31:0] _GEN_20048 = read_stack9_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_20017; // @[lut_35.scala 4049:77 lut_35.scala 4088:41]
  wire  _GEN_20051 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _T_778; // @[lut_35.scala 4008:77 lut_35.scala 4018:44]
  wire  _GEN_20052 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20020; // @[lut_35.scala 4008:77 lut_35.scala 4019:45]
  wire  _GEN_20053 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20021; // @[lut_35.scala 4008:77 lut_35.scala 4020:45]
  wire  _GEN_20054 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20022; // @[lut_35.scala 4008:77 lut_35.scala 4021:45]
  wire  _GEN_20055 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20023; // @[lut_35.scala 4008:77 lut_35.scala 4022:45]
  wire  _GEN_20056 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20024; // @[lut_35.scala 4008:77 lut_35.scala 4023:45]
  wire  _GEN_20057 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20025; // @[lut_35.scala 4008:77 lut_35.scala 4024:45]
  wire  _GEN_20058 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20026; // @[lut_35.scala 4008:77 lut_35.scala 4025:45]
  wire  _GEN_20059 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20027; // @[lut_35.scala 4008:77 lut_35.scala 4026:45]
  wire  _GEN_20060 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20028; // @[lut_35.scala 4008:77 lut_35.scala 4027:45]
  wire  _GEN_20061 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20029; // @[lut_35.scala 4008:77 lut_35.scala 4028:45]
  wire  _GEN_20062 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20030; // @[lut_35.scala 4008:77 lut_35.scala 4029:45]
  wire  _GEN_20063 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20031; // @[lut_35.scala 4008:77 lut_35.scala 4030:45]
  wire  _GEN_20064 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20032; // @[lut_35.scala 4008:77 lut_35.scala 4031:45]
  wire  _GEN_20065 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20033; // @[lut_35.scala 4008:77 lut_35.scala 4032:45]
  wire  _GEN_20066 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20034; // @[lut_35.scala 4008:77 lut_35.scala 4033:45]
  wire  _GEN_20067 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20035; // @[lut_35.scala 4008:77 lut_35.scala 4034:45]
  wire  _GEN_20068 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20036; // @[lut_35.scala 4008:77 lut_35.scala 4035:45]
  wire  _GEN_20069 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20037; // @[lut_35.scala 4008:77 lut_35.scala 4036:45]
  wire  _GEN_20070 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20038; // @[lut_35.scala 4008:77 lut_35.scala 4037:45]
  wire  _GEN_20071 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20039; // @[lut_35.scala 4008:77 lut_35.scala 4038:45]
  wire  _GEN_20072 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20040; // @[lut_35.scala 4008:77 lut_35.scala 4039:45]
  wire  _GEN_20073 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20041; // @[lut_35.scala 4008:77 lut_35.scala 4040:45]
  wire  _GEN_20074 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20042; // @[lut_35.scala 4008:77 lut_35.scala 4041:45]
  wire  _GEN_20075 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20043; // @[lut_35.scala 4008:77 lut_35.scala 4042:45]
  wire  _GEN_20076 = read_stack8_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20044; // @[lut_35.scala 4008:77 lut_35.scala 4043:45]
  wire  _GEN_20077 = read_stack8_pop == pop_ray_id & pop_valid | _GEN_20045; // @[lut_35.scala 4008:77 lut_35.scala 4044:40]
  wire [31:0] _GEN_20079 = read_stack8_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_20047; // @[lut_35.scala 4008:77 lut_35.scala 4046:38]
  wire [31:0] _GEN_20080 = read_stack8_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_20048; // @[lut_35.scala 4008:77 lut_35.scala 4047:41]
  wire  _GEN_20083 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _T_775; // @[lut_35.scala 3968:77 lut_35.scala 3977:44]
  wire  _GEN_20084 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20051; // @[lut_35.scala 3968:77 lut_35.scala 3978:44]
  wire  _GEN_20085 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20052; // @[lut_35.scala 3968:77 lut_35.scala 3979:45]
  wire  _GEN_20086 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20053; // @[lut_35.scala 3968:77 lut_35.scala 3980:45]
  wire  _GEN_20087 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20054; // @[lut_35.scala 3968:77 lut_35.scala 3981:45]
  wire  _GEN_20088 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20055; // @[lut_35.scala 3968:77 lut_35.scala 3982:45]
  wire  _GEN_20089 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20056; // @[lut_35.scala 3968:77 lut_35.scala 3983:45]
  wire  _GEN_20090 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20057; // @[lut_35.scala 3968:77 lut_35.scala 3984:45]
  wire  _GEN_20091 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20058; // @[lut_35.scala 3968:77 lut_35.scala 3985:45]
  wire  _GEN_20092 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20059; // @[lut_35.scala 3968:77 lut_35.scala 3986:45]
  wire  _GEN_20093 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20060; // @[lut_35.scala 3968:77 lut_35.scala 3987:45]
  wire  _GEN_20094 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20061; // @[lut_35.scala 3968:77 lut_35.scala 3988:45]
  wire  _GEN_20095 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20062; // @[lut_35.scala 3968:77 lut_35.scala 3989:45]
  wire  _GEN_20096 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20063; // @[lut_35.scala 3968:77 lut_35.scala 3990:45]
  wire  _GEN_20097 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20064; // @[lut_35.scala 3968:77 lut_35.scala 3991:45]
  wire  _GEN_20098 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20065; // @[lut_35.scala 3968:77 lut_35.scala 3992:45]
  wire  _GEN_20099 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20066; // @[lut_35.scala 3968:77 lut_35.scala 3993:45]
  wire  _GEN_20100 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20067; // @[lut_35.scala 3968:77 lut_35.scala 3994:45]
  wire  _GEN_20101 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20068; // @[lut_35.scala 3968:77 lut_35.scala 3995:45]
  wire  _GEN_20102 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20069; // @[lut_35.scala 3968:77 lut_35.scala 3996:45]
  wire  _GEN_20103 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20070; // @[lut_35.scala 3968:77 lut_35.scala 3997:45]
  wire  _GEN_20104 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20071; // @[lut_35.scala 3968:77 lut_35.scala 3998:45]
  wire  _GEN_20105 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20072; // @[lut_35.scala 3968:77 lut_35.scala 3999:45]
  wire  _GEN_20106 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20073; // @[lut_35.scala 3968:77 lut_35.scala 4000:45]
  wire  _GEN_20107 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20074; // @[lut_35.scala 3968:77 lut_35.scala 4001:45]
  wire  _GEN_20108 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20075; // @[lut_35.scala 3968:77 lut_35.scala 4002:45]
  wire  _GEN_20109 = read_stack7_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20076; // @[lut_35.scala 3968:77 lut_35.scala 4003:45]
  wire  _GEN_20110 = read_stack7_pop == pop_ray_id & pop_valid | _GEN_20077; // @[lut_35.scala 3968:77 lut_35.scala 4004:40]
  wire [31:0] _GEN_20112 = read_stack7_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_20079; // @[lut_35.scala 3968:77 lut_35.scala 4006:38]
  wire [31:0] _GEN_20113 = read_stack7_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_20080; // @[lut_35.scala 3968:77 lut_35.scala 4007:41]
  wire  _GEN_20116 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _T_772; // @[lut_35.scala 3928:77 lut_35.scala 3936:44]
  wire  _GEN_20117 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20083; // @[lut_35.scala 3928:77 lut_35.scala 3937:44]
  wire  _GEN_20118 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20084; // @[lut_35.scala 3928:77 lut_35.scala 3938:44]
  wire  _GEN_20119 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20085; // @[lut_35.scala 3928:77 lut_35.scala 3939:45]
  wire  _GEN_20120 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20086; // @[lut_35.scala 3928:77 lut_35.scala 3940:45]
  wire  _GEN_20121 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20087; // @[lut_35.scala 3928:77 lut_35.scala 3941:45]
  wire  _GEN_20122 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20088; // @[lut_35.scala 3928:77 lut_35.scala 3942:45]
  wire  _GEN_20123 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20089; // @[lut_35.scala 3928:77 lut_35.scala 3943:45]
  wire  _GEN_20124 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20090; // @[lut_35.scala 3928:77 lut_35.scala 3944:45]
  wire  _GEN_20125 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20091; // @[lut_35.scala 3928:77 lut_35.scala 3945:45]
  wire  _GEN_20126 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20092; // @[lut_35.scala 3928:77 lut_35.scala 3946:45]
  wire  _GEN_20127 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20093; // @[lut_35.scala 3928:77 lut_35.scala 3947:45]
  wire  _GEN_20128 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20094; // @[lut_35.scala 3928:77 lut_35.scala 3948:45]
  wire  _GEN_20129 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20095; // @[lut_35.scala 3928:77 lut_35.scala 3949:45]
  wire  _GEN_20130 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20096; // @[lut_35.scala 3928:77 lut_35.scala 3950:45]
  wire  _GEN_20131 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20097; // @[lut_35.scala 3928:77 lut_35.scala 3951:45]
  wire  _GEN_20132 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20098; // @[lut_35.scala 3928:77 lut_35.scala 3952:45]
  wire  _GEN_20133 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20099; // @[lut_35.scala 3928:77 lut_35.scala 3953:45]
  wire  _GEN_20134 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20100; // @[lut_35.scala 3928:77 lut_35.scala 3954:45]
  wire  _GEN_20135 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20101; // @[lut_35.scala 3928:77 lut_35.scala 3955:45]
  wire  _GEN_20136 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20102; // @[lut_35.scala 3928:77 lut_35.scala 3956:45]
  wire  _GEN_20137 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20103; // @[lut_35.scala 3928:77 lut_35.scala 3957:45]
  wire  _GEN_20138 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20104; // @[lut_35.scala 3928:77 lut_35.scala 3958:45]
  wire  _GEN_20139 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20105; // @[lut_35.scala 3928:77 lut_35.scala 3959:45]
  wire  _GEN_20140 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20106; // @[lut_35.scala 3928:77 lut_35.scala 3960:45]
  wire  _GEN_20141 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20107; // @[lut_35.scala 3928:77 lut_35.scala 3961:45]
  wire  _GEN_20142 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20108; // @[lut_35.scala 3928:77 lut_35.scala 3962:45]
  wire  _GEN_20143 = read_stack6_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20109; // @[lut_35.scala 3928:77 lut_35.scala 3963:45]
  wire  _GEN_20144 = read_stack6_pop == pop_ray_id & pop_valid | _GEN_20110; // @[lut_35.scala 3928:77 lut_35.scala 3964:40]
  wire [31:0] _GEN_20146 = read_stack6_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_20112; // @[lut_35.scala 3928:77 lut_35.scala 3966:38]
  wire [31:0] _GEN_20147 = read_stack6_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_20113; // @[lut_35.scala 3928:77 lut_35.scala 3967:41]
  wire  _GEN_20150 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _T_769; // @[lut_35.scala 3888:77 lut_35.scala 3895:44]
  wire  _GEN_20151 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20116; // @[lut_35.scala 3888:77 lut_35.scala 3896:44]
  wire  _GEN_20152 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20117; // @[lut_35.scala 3888:77 lut_35.scala 3897:44]
  wire  _GEN_20153 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20118; // @[lut_35.scala 3888:77 lut_35.scala 3898:44]
  wire  _GEN_20154 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20119; // @[lut_35.scala 3888:77 lut_35.scala 3899:45]
  wire  _GEN_20155 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20120; // @[lut_35.scala 3888:77 lut_35.scala 3900:45]
  wire  _GEN_20156 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20121; // @[lut_35.scala 3888:77 lut_35.scala 3901:45]
  wire  _GEN_20157 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20122; // @[lut_35.scala 3888:77 lut_35.scala 3902:45]
  wire  _GEN_20158 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20123; // @[lut_35.scala 3888:77 lut_35.scala 3903:45]
  wire  _GEN_20159 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20124; // @[lut_35.scala 3888:77 lut_35.scala 3904:45]
  wire  _GEN_20160 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20125; // @[lut_35.scala 3888:77 lut_35.scala 3905:45]
  wire  _GEN_20161 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20126; // @[lut_35.scala 3888:77 lut_35.scala 3906:45]
  wire  _GEN_20162 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20127; // @[lut_35.scala 3888:77 lut_35.scala 3907:45]
  wire  _GEN_20163 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20128; // @[lut_35.scala 3888:77 lut_35.scala 3908:45]
  wire  _GEN_20164 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20129; // @[lut_35.scala 3888:77 lut_35.scala 3909:45]
  wire  _GEN_20165 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20130; // @[lut_35.scala 3888:77 lut_35.scala 3910:45]
  wire  _GEN_20166 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20131; // @[lut_35.scala 3888:77 lut_35.scala 3911:45]
  wire  _GEN_20167 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20132; // @[lut_35.scala 3888:77 lut_35.scala 3912:45]
  wire  _GEN_20168 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20133; // @[lut_35.scala 3888:77 lut_35.scala 3913:45]
  wire  _GEN_20169 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20134; // @[lut_35.scala 3888:77 lut_35.scala 3914:45]
  wire  _GEN_20170 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20135; // @[lut_35.scala 3888:77 lut_35.scala 3915:45]
  wire  _GEN_20171 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20136; // @[lut_35.scala 3888:77 lut_35.scala 3916:45]
  wire  _GEN_20172 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20137; // @[lut_35.scala 3888:77 lut_35.scala 3917:45]
  wire  _GEN_20173 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20138; // @[lut_35.scala 3888:77 lut_35.scala 3918:45]
  wire  _GEN_20174 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20139; // @[lut_35.scala 3888:77 lut_35.scala 3919:45]
  wire  _GEN_20175 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20140; // @[lut_35.scala 3888:77 lut_35.scala 3920:45]
  wire  _GEN_20176 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20141; // @[lut_35.scala 3888:77 lut_35.scala 3921:45]
  wire  _GEN_20177 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20142; // @[lut_35.scala 3888:77 lut_35.scala 3922:45]
  wire  _GEN_20178 = read_stack5_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20143; // @[lut_35.scala 3888:77 lut_35.scala 3923:45]
  wire  _GEN_20179 = read_stack5_pop == pop_ray_id & pop_valid | _GEN_20144; // @[lut_35.scala 3888:77 lut_35.scala 3924:40]
  wire [31:0] _GEN_20181 = read_stack5_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_20146; // @[lut_35.scala 3888:77 lut_35.scala 3926:38]
  wire [31:0] _GEN_20182 = read_stack5_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_20147; // @[lut_35.scala 3888:77 lut_35.scala 3927:41]
  wire  _GEN_20185 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _T_766; // @[lut_35.scala 3848:77 lut_35.scala 3854:44]
  wire  _GEN_20186 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20150; // @[lut_35.scala 3848:77 lut_35.scala 3855:44]
  wire  _GEN_20187 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20151; // @[lut_35.scala 3848:77 lut_35.scala 3856:44]
  wire  _GEN_20188 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20152; // @[lut_35.scala 3848:77 lut_35.scala 3857:44]
  wire  _GEN_20189 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20153; // @[lut_35.scala 3848:77 lut_35.scala 3858:44]
  wire  _GEN_20190 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20154; // @[lut_35.scala 3848:77 lut_35.scala 3859:45]
  wire  _GEN_20191 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20155; // @[lut_35.scala 3848:77 lut_35.scala 3860:45]
  wire  _GEN_20192 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20156; // @[lut_35.scala 3848:77 lut_35.scala 3861:45]
  wire  _GEN_20193 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20157; // @[lut_35.scala 3848:77 lut_35.scala 3862:45]
  wire  _GEN_20194 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20158; // @[lut_35.scala 3848:77 lut_35.scala 3863:45]
  wire  _GEN_20195 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20159; // @[lut_35.scala 3848:77 lut_35.scala 3864:45]
  wire  _GEN_20196 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20160; // @[lut_35.scala 3848:77 lut_35.scala 3865:45]
  wire  _GEN_20197 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20161; // @[lut_35.scala 3848:77 lut_35.scala 3866:45]
  wire  _GEN_20198 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20162; // @[lut_35.scala 3848:77 lut_35.scala 3867:45]
  wire  _GEN_20199 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20163; // @[lut_35.scala 3848:77 lut_35.scala 3868:45]
  wire  _GEN_20200 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20164; // @[lut_35.scala 3848:77 lut_35.scala 3869:45]
  wire  _GEN_20201 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20165; // @[lut_35.scala 3848:77 lut_35.scala 3870:45]
  wire  _GEN_20202 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20166; // @[lut_35.scala 3848:77 lut_35.scala 3871:45]
  wire  _GEN_20203 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20167; // @[lut_35.scala 3848:77 lut_35.scala 3872:45]
  wire  _GEN_20204 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20168; // @[lut_35.scala 3848:77 lut_35.scala 3873:45]
  wire  _GEN_20205 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20169; // @[lut_35.scala 3848:77 lut_35.scala 3874:45]
  wire  _GEN_20206 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20170; // @[lut_35.scala 3848:77 lut_35.scala 3875:45]
  wire  _GEN_20207 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20171; // @[lut_35.scala 3848:77 lut_35.scala 3876:45]
  wire  _GEN_20208 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20172; // @[lut_35.scala 3848:77 lut_35.scala 3877:45]
  wire  _GEN_20209 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20173; // @[lut_35.scala 3848:77 lut_35.scala 3878:45]
  wire  _GEN_20210 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20174; // @[lut_35.scala 3848:77 lut_35.scala 3879:45]
  wire  _GEN_20211 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20175; // @[lut_35.scala 3848:77 lut_35.scala 3880:45]
  wire  _GEN_20212 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20176; // @[lut_35.scala 3848:77 lut_35.scala 3881:45]
  wire  _GEN_20213 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20177; // @[lut_35.scala 3848:77 lut_35.scala 3882:45]
  wire  _GEN_20214 = read_stack4_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20178; // @[lut_35.scala 3848:77 lut_35.scala 3883:45]
  wire  _GEN_20215 = read_stack4_pop == pop_ray_id & pop_valid | _GEN_20179; // @[lut_35.scala 3848:77 lut_35.scala 3884:40]
  wire [31:0] _GEN_20217 = read_stack4_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_20181; // @[lut_35.scala 3848:77 lut_35.scala 3886:38]
  wire [31:0] _GEN_20218 = read_stack4_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_20182; // @[lut_35.scala 3848:77 lut_35.scala 3887:41]
  wire  _GEN_20221 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _T_763; // @[lut_35.scala 3808:77 lut_35.scala 3813:44]
  wire  _GEN_20222 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20185; // @[lut_35.scala 3808:77 lut_35.scala 3814:44]
  wire  _GEN_20223 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20186; // @[lut_35.scala 3808:77 lut_35.scala 3815:44]
  wire  _GEN_20224 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20187; // @[lut_35.scala 3808:77 lut_35.scala 3816:44]
  wire  _GEN_20225 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20188; // @[lut_35.scala 3808:77 lut_35.scala 3817:44]
  wire  _GEN_20226 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20189; // @[lut_35.scala 3808:77 lut_35.scala 3818:44]
  wire  _GEN_20227 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20190; // @[lut_35.scala 3808:77 lut_35.scala 3819:45]
  wire  _GEN_20228 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20191; // @[lut_35.scala 3808:77 lut_35.scala 3820:45]
  wire  _GEN_20229 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20192; // @[lut_35.scala 3808:77 lut_35.scala 3821:45]
  wire  _GEN_20230 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20193; // @[lut_35.scala 3808:77 lut_35.scala 3822:45]
  wire  _GEN_20231 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20194; // @[lut_35.scala 3808:77 lut_35.scala 3823:45]
  wire  _GEN_20232 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20195; // @[lut_35.scala 3808:77 lut_35.scala 3824:45]
  wire  _GEN_20233 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20196; // @[lut_35.scala 3808:77 lut_35.scala 3825:45]
  wire  _GEN_20234 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20197; // @[lut_35.scala 3808:77 lut_35.scala 3826:45]
  wire  _GEN_20235 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20198; // @[lut_35.scala 3808:77 lut_35.scala 3827:45]
  wire  _GEN_20236 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20199; // @[lut_35.scala 3808:77 lut_35.scala 3828:45]
  wire  _GEN_20237 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20200; // @[lut_35.scala 3808:77 lut_35.scala 3829:45]
  wire  _GEN_20238 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20201; // @[lut_35.scala 3808:77 lut_35.scala 3830:45]
  wire  _GEN_20239 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20202; // @[lut_35.scala 3808:77 lut_35.scala 3831:45]
  wire  _GEN_20240 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20203; // @[lut_35.scala 3808:77 lut_35.scala 3832:45]
  wire  _GEN_20241 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20204; // @[lut_35.scala 3808:77 lut_35.scala 3833:45]
  wire  _GEN_20242 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20205; // @[lut_35.scala 3808:77 lut_35.scala 3834:45]
  wire  _GEN_20243 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20206; // @[lut_35.scala 3808:77 lut_35.scala 3835:45]
  wire  _GEN_20244 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20207; // @[lut_35.scala 3808:77 lut_35.scala 3836:45]
  wire  _GEN_20245 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20208; // @[lut_35.scala 3808:77 lut_35.scala 3837:45]
  wire  _GEN_20246 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20209; // @[lut_35.scala 3808:77 lut_35.scala 3838:45]
  wire  _GEN_20247 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20210; // @[lut_35.scala 3808:77 lut_35.scala 3839:45]
  wire  _GEN_20248 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20211; // @[lut_35.scala 3808:77 lut_35.scala 3840:45]
  wire  _GEN_20249 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20212; // @[lut_35.scala 3808:77 lut_35.scala 3841:45]
  wire  _GEN_20250 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20213; // @[lut_35.scala 3808:77 lut_35.scala 3842:45]
  wire  _GEN_20251 = read_stack3_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20214; // @[lut_35.scala 3808:77 lut_35.scala 3843:45]
  wire  _GEN_20252 = read_stack3_pop == pop_ray_id & pop_valid | _GEN_20215; // @[lut_35.scala 3808:77 lut_35.scala 3844:40]
  wire [31:0] _GEN_20254 = read_stack3_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_20217; // @[lut_35.scala 3808:77 lut_35.scala 3846:38]
  wire [31:0] _GEN_20255 = read_stack3_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_20218; // @[lut_35.scala 3808:77 lut_35.scala 3847:41]
  wire  _GEN_20258 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _T_760; // @[lut_35.scala 3768:77 lut_35.scala 3772:44]
  wire  _GEN_20259 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20221; // @[lut_35.scala 3768:77 lut_35.scala 3773:44]
  wire  _GEN_20260 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20222; // @[lut_35.scala 3768:77 lut_35.scala 3774:44]
  wire  _GEN_20261 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20223; // @[lut_35.scala 3768:77 lut_35.scala 3775:44]
  wire  _GEN_20262 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20224; // @[lut_35.scala 3768:77 lut_35.scala 3776:44]
  wire  _GEN_20263 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20225; // @[lut_35.scala 3768:77 lut_35.scala 3777:44]
  wire  _GEN_20264 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20226; // @[lut_35.scala 3768:77 lut_35.scala 3778:44]
  wire  _GEN_20265 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20227; // @[lut_35.scala 3768:77 lut_35.scala 3779:45]
  wire  _GEN_20266 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20228; // @[lut_35.scala 3768:77 lut_35.scala 3780:45]
  wire  _GEN_20267 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20229; // @[lut_35.scala 3768:77 lut_35.scala 3781:45]
  wire  _GEN_20268 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20230; // @[lut_35.scala 3768:77 lut_35.scala 3782:45]
  wire  _GEN_20269 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20231; // @[lut_35.scala 3768:77 lut_35.scala 3783:45]
  wire  _GEN_20270 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20232; // @[lut_35.scala 3768:77 lut_35.scala 3784:45]
  wire  _GEN_20271 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20233; // @[lut_35.scala 3768:77 lut_35.scala 3785:45]
  wire  _GEN_20272 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20234; // @[lut_35.scala 3768:77 lut_35.scala 3786:45]
  wire  _GEN_20273 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20235; // @[lut_35.scala 3768:77 lut_35.scala 3787:45]
  wire  _GEN_20274 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20236; // @[lut_35.scala 3768:77 lut_35.scala 3788:45]
  wire  _GEN_20275 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20237; // @[lut_35.scala 3768:77 lut_35.scala 3789:45]
  wire  _GEN_20276 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20238; // @[lut_35.scala 3768:77 lut_35.scala 3790:45]
  wire  _GEN_20277 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20239; // @[lut_35.scala 3768:77 lut_35.scala 3791:45]
  wire  _GEN_20278 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20240; // @[lut_35.scala 3768:77 lut_35.scala 3792:45]
  wire  _GEN_20279 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20241; // @[lut_35.scala 3768:77 lut_35.scala 3793:45]
  wire  _GEN_20280 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20242; // @[lut_35.scala 3768:77 lut_35.scala 3794:45]
  wire  _GEN_20281 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20243; // @[lut_35.scala 3768:77 lut_35.scala 3795:45]
  wire  _GEN_20282 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20244; // @[lut_35.scala 3768:77 lut_35.scala 3796:45]
  wire  _GEN_20283 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20245; // @[lut_35.scala 3768:77 lut_35.scala 3797:45]
  wire  _GEN_20284 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20246; // @[lut_35.scala 3768:77 lut_35.scala 3798:45]
  wire  _GEN_20285 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20247; // @[lut_35.scala 3768:77 lut_35.scala 3799:45]
  wire  _GEN_20286 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20248; // @[lut_35.scala 3768:77 lut_35.scala 3800:45]
  wire  _GEN_20287 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20249; // @[lut_35.scala 3768:77 lut_35.scala 3801:45]
  wire  _GEN_20288 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20250; // @[lut_35.scala 3768:77 lut_35.scala 3802:45]
  wire  _GEN_20289 = read_stack2_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20251; // @[lut_35.scala 3768:77 lut_35.scala 3803:45]
  wire  _GEN_20290 = read_stack2_pop == pop_ray_id & pop_valid | _GEN_20252; // @[lut_35.scala 3768:77 lut_35.scala 3804:40]
  wire [31:0] _GEN_20292 = read_stack2_pop == pop_ray_id & pop_valid ? pop_ray_id : _GEN_20254; // @[lut_35.scala 3768:77 lut_35.scala 3806:38]
  wire [31:0] _GEN_20293 = read_stack2_pop == pop_ray_id & pop_valid ? pop_hitT_1 : _GEN_20255; // @[lut_35.scala 3768:77 lut_35.scala 3807:41]
  wire  _GEN_20296 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _T_757; // @[lut_35.scala 3728:77 lut_35.scala 3731:44]
  wire  _GEN_20297 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20258; // @[lut_35.scala 3728:77 lut_35.scala 3732:44]
  wire  _GEN_20298 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20259; // @[lut_35.scala 3728:77 lut_35.scala 3733:44]
  wire  _GEN_20299 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20260; // @[lut_35.scala 3728:77 lut_35.scala 3734:44]
  wire  _GEN_20300 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20261; // @[lut_35.scala 3728:77 lut_35.scala 3735:44]
  wire  _GEN_20301 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20262; // @[lut_35.scala 3728:77 lut_35.scala 3736:44]
  wire  _GEN_20302 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20263; // @[lut_35.scala 3728:77 lut_35.scala 3737:44]
  wire  _GEN_20303 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20264; // @[lut_35.scala 3728:77 lut_35.scala 3738:44]
  wire  _GEN_20304 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20265; // @[lut_35.scala 3728:77 lut_35.scala 3739:45]
  wire  _GEN_20305 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20266; // @[lut_35.scala 3728:77 lut_35.scala 3740:45]
  wire  _GEN_20306 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20267; // @[lut_35.scala 3728:77 lut_35.scala 3741:45]
  wire  _GEN_20307 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20268; // @[lut_35.scala 3728:77 lut_35.scala 3742:45]
  wire  _GEN_20308 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20269; // @[lut_35.scala 3728:77 lut_35.scala 3743:45]
  wire  _GEN_20309 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20270; // @[lut_35.scala 3728:77 lut_35.scala 3744:45]
  wire  _GEN_20310 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20271; // @[lut_35.scala 3728:77 lut_35.scala 3745:45]
  wire  _GEN_20311 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20272; // @[lut_35.scala 3728:77 lut_35.scala 3746:45]
  wire  _GEN_20312 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20273; // @[lut_35.scala 3728:77 lut_35.scala 3747:45]
  wire  _GEN_20313 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20274; // @[lut_35.scala 3728:77 lut_35.scala 3748:45]
  wire  _GEN_20314 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20275; // @[lut_35.scala 3728:77 lut_35.scala 3749:45]
  wire  _GEN_20315 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20276; // @[lut_35.scala 3728:77 lut_35.scala 3750:45]
  wire  _GEN_20316 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20277; // @[lut_35.scala 3728:77 lut_35.scala 3751:45]
  wire  _GEN_20317 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20278; // @[lut_35.scala 3728:77 lut_35.scala 3752:45]
  wire  _GEN_20318 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20279; // @[lut_35.scala 3728:77 lut_35.scala 3753:45]
  wire  _GEN_20319 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20280; // @[lut_35.scala 3728:77 lut_35.scala 3754:45]
  wire  _GEN_20320 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20281; // @[lut_35.scala 3728:77 lut_35.scala 3755:45]
  wire  _GEN_20321 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20282; // @[lut_35.scala 3728:77 lut_35.scala 3756:45]
  wire  _GEN_20322 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20283; // @[lut_35.scala 3728:77 lut_35.scala 3757:45]
  wire  _GEN_20323 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20284; // @[lut_35.scala 3728:77 lut_35.scala 3758:45]
  wire  _GEN_20324 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20285; // @[lut_35.scala 3728:77 lut_35.scala 3759:45]
  wire  _GEN_20325 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20286; // @[lut_35.scala 3728:77 lut_35.scala 3760:45]
  wire  _GEN_20326 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20287; // @[lut_35.scala 3728:77 lut_35.scala 3761:45]
  wire  _GEN_20327 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20288; // @[lut_35.scala 3728:77 lut_35.scala 3762:45]
  wire  _GEN_20328 = read_stack1_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20289; // @[lut_35.scala 3728:77 lut_35.scala 3763:45]
  wire  _GEN_20329 = read_stack1_pop == pop_ray_id & pop_valid | _GEN_20290; // @[lut_35.scala 3728:77 lut_35.scala 3764:40]
  wire  _GEN_20334 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _T_754; // @[lut_35.scala 3688:67 lut_35.scala 3690:40]
  wire  _GEN_20335 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20296; // @[lut_35.scala 3688:67 lut_35.scala 3691:40]
  wire  _GEN_20336 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20297; // @[lut_35.scala 3688:67 lut_35.scala 3692:40]
  wire  _GEN_20337 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20298; // @[lut_35.scala 3688:67 lut_35.scala 3693:40]
  wire  _GEN_20338 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20299; // @[lut_35.scala 3688:67 lut_35.scala 3694:40]
  wire  _GEN_20339 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20300; // @[lut_35.scala 3688:67 lut_35.scala 3695:40]
  wire  _GEN_20340 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20301; // @[lut_35.scala 3688:67 lut_35.scala 3696:40]
  wire  _GEN_20341 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20302; // @[lut_35.scala 3688:67 lut_35.scala 3697:40]
  wire  _GEN_20342 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20303; // @[lut_35.scala 3688:67 lut_35.scala 3698:40]
  wire  _GEN_20343 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20304; // @[lut_35.scala 3688:67 lut_35.scala 3699:41]
  wire  _GEN_20344 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20305; // @[lut_35.scala 3688:67 lut_35.scala 3700:41]
  wire  _GEN_20345 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20306; // @[lut_35.scala 3688:67 lut_35.scala 3701:41]
  wire  _GEN_20346 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20307; // @[lut_35.scala 3688:67 lut_35.scala 3702:41]
  wire  _GEN_20347 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20308; // @[lut_35.scala 3688:67 lut_35.scala 3703:41]
  wire  _GEN_20348 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20309; // @[lut_35.scala 3688:67 lut_35.scala 3704:41]
  wire  _GEN_20349 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20310; // @[lut_35.scala 3688:67 lut_35.scala 3705:41]
  wire  _GEN_20350 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20311; // @[lut_35.scala 3688:67 lut_35.scala 3706:41]
  wire  _GEN_20351 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20312; // @[lut_35.scala 3688:67 lut_35.scala 3707:41]
  wire  _GEN_20352 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20313; // @[lut_35.scala 3688:67 lut_35.scala 3708:41]
  wire  _GEN_20353 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20314; // @[lut_35.scala 3688:67 lut_35.scala 3709:41]
  wire  _GEN_20354 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20315; // @[lut_35.scala 3688:67 lut_35.scala 3710:41]
  wire  _GEN_20355 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20316; // @[lut_35.scala 3688:67 lut_35.scala 3711:41]
  wire  _GEN_20356 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20317; // @[lut_35.scala 3688:67 lut_35.scala 3712:41]
  wire  _GEN_20357 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20318; // @[lut_35.scala 3688:67 lut_35.scala 3713:41]
  wire  _GEN_20358 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20319; // @[lut_35.scala 3688:67 lut_35.scala 3714:41]
  wire  _GEN_20359 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20320; // @[lut_35.scala 3688:67 lut_35.scala 3715:41]
  wire  _GEN_20360 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20321; // @[lut_35.scala 3688:67 lut_35.scala 3716:41]
  wire  _GEN_20361 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20322; // @[lut_35.scala 3688:67 lut_35.scala 3717:41]
  wire  _GEN_20362 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20323; // @[lut_35.scala 3688:67 lut_35.scala 3718:41]
  wire  _GEN_20363 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20324; // @[lut_35.scala 3688:67 lut_35.scala 3719:41]
  wire  _GEN_20364 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20325; // @[lut_35.scala 3688:67 lut_35.scala 3720:41]
  wire  _GEN_20365 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20326; // @[lut_35.scala 3688:67 lut_35.scala 3721:41]
  wire  _GEN_20366 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20327; // @[lut_35.scala 3688:67 lut_35.scala 3722:41]
  wire  _GEN_20367 = read_stack0_pop == pop_ray_id & pop_valid ? 1'h0 : _GEN_20328; // @[lut_35.scala 3688:67 lut_35.scala 3723:41]
  wire  _GEN_20368 = read_stack0_pop == pop_ray_id & pop_valid | _GEN_20329; // @[lut_35.scala 3688:67 lut_35.scala 3724:36]
  wire  _GEN_20372 = pop_1 & pop_valid & _T_751; // @[lut_35.scala 3687:46 lut_35.scala 5128:40]
  wire  _GEN_20373 = pop_1 & pop_valid & _GEN_20334; // @[lut_35.scala 3687:46 lut_35.scala 5129:40]
  wire  _GEN_20374 = pop_1 & pop_valid & _GEN_20335; // @[lut_35.scala 3687:46 lut_35.scala 5130:40]
  wire  _GEN_20375 = pop_1 & pop_valid & _GEN_20336; // @[lut_35.scala 3687:46 lut_35.scala 5131:40]
  wire  _GEN_20376 = pop_1 & pop_valid & _GEN_20337; // @[lut_35.scala 3687:46 lut_35.scala 5132:40]
  wire  _GEN_20377 = pop_1 & pop_valid & _GEN_20338; // @[lut_35.scala 3687:46 lut_35.scala 5133:40]
  wire  _GEN_20378 = pop_1 & pop_valid & _GEN_20339; // @[lut_35.scala 3687:46 lut_35.scala 5134:40]
  wire  _GEN_20379 = pop_1 & pop_valid & _GEN_20340; // @[lut_35.scala 3687:46 lut_35.scala 5135:40]
  wire  _GEN_20380 = pop_1 & pop_valid & _GEN_20341; // @[lut_35.scala 3687:46 lut_35.scala 5136:40]
  wire  _GEN_20381 = pop_1 & pop_valid & _GEN_20342; // @[lut_35.scala 3687:46 lut_35.scala 5137:40]
  wire  _GEN_20382 = pop_1 & pop_valid & _GEN_20343; // @[lut_35.scala 3687:46 lut_35.scala 5138:41]
  wire  _GEN_20383 = pop_1 & pop_valid & _GEN_20344; // @[lut_35.scala 3687:46 lut_35.scala 5139:41]
  wire  _GEN_20384 = pop_1 & pop_valid & _GEN_20345; // @[lut_35.scala 3687:46 lut_35.scala 5140:41]
  wire  _GEN_20385 = pop_1 & pop_valid & _GEN_20346; // @[lut_35.scala 3687:46 lut_35.scala 5141:41]
  wire  _GEN_20386 = pop_1 & pop_valid & _GEN_20347; // @[lut_35.scala 3687:46 lut_35.scala 5142:41]
  wire  _GEN_20387 = pop_1 & pop_valid & _GEN_20348; // @[lut_35.scala 3687:46 lut_35.scala 5143:41]
  wire  _GEN_20388 = pop_1 & pop_valid & _GEN_20349; // @[lut_35.scala 3687:46 lut_35.scala 5144:41]
  wire  _GEN_20389 = pop_1 & pop_valid & _GEN_20350; // @[lut_35.scala 3687:46 lut_35.scala 5145:41]
  wire  _GEN_20390 = pop_1 & pop_valid & _GEN_20351; // @[lut_35.scala 3687:46 lut_35.scala 5146:41]
  wire  _GEN_20391 = pop_1 & pop_valid & _GEN_20352; // @[lut_35.scala 3687:46 lut_35.scala 5147:41]
  wire  _GEN_20392 = pop_1 & pop_valid & _GEN_20353; // @[lut_35.scala 3687:46 lut_35.scala 5148:41]
  wire  _GEN_20393 = pop_1 & pop_valid & _GEN_20354; // @[lut_35.scala 3687:46 lut_35.scala 5149:41]
  wire  _GEN_20394 = pop_1 & pop_valid & _GEN_20355; // @[lut_35.scala 3687:46 lut_35.scala 5150:41]
  wire  _GEN_20395 = pop_1 & pop_valid & _GEN_20356; // @[lut_35.scala 3687:46 lut_35.scala 5151:41]
  wire  _GEN_20396 = pop_1 & pop_valid & _GEN_20357; // @[lut_35.scala 3687:46 lut_35.scala 5152:41]
  wire  _GEN_20397 = pop_1 & pop_valid & _GEN_20358; // @[lut_35.scala 3687:46 lut_35.scala 5153:41]
  wire  _GEN_20398 = pop_1 & pop_valid & _GEN_20359; // @[lut_35.scala 3687:46 lut_35.scala 5154:41]
  wire  _GEN_20399 = pop_1 & pop_valid & _GEN_20360; // @[lut_35.scala 3687:46 lut_35.scala 5155:41]
  wire  _GEN_20400 = pop_1 & pop_valid & _GEN_20361; // @[lut_35.scala 3687:46 lut_35.scala 5156:41]
  wire  _GEN_20401 = pop_1 & pop_valid & _GEN_20362; // @[lut_35.scala 3687:46 lut_35.scala 5157:41]
  wire  _GEN_20402 = pop_1 & pop_valid & _GEN_20363; // @[lut_35.scala 3687:46 lut_35.scala 5158:41]
  wire  _GEN_20403 = pop_1 & pop_valid & _GEN_20364; // @[lut_35.scala 3687:46 lut_35.scala 5159:41]
  wire  _GEN_20404 = pop_1 & pop_valid & _GEN_20365; // @[lut_35.scala 3687:46 lut_35.scala 5160:41]
  wire  _GEN_20405 = pop_1 & pop_valid & _GEN_20366; // @[lut_35.scala 3687:46 lut_35.scala 5161:41]
  wire  _GEN_20406 = pop_1 & pop_valid & _GEN_20367; // @[lut_35.scala 3687:46 lut_35.scala 5162:41]
  wire  _GEN_20407 = pop_1 & pop_valid & _GEN_20368; // @[lut_35.scala 3687:46 lut_35.scala 5163:37]
  assign LUT_mem_MPORT_1_addr = 6'h0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_1_data = LUT_mem[LUT_mem_MPORT_1_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_1_data = LUT_mem_MPORT_1_addr >= 6'h23 ? _RAND_1[32:0] : LUT_mem[LUT_mem_MPORT_1_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_3_addr = 6'h0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_3_data = LUT_mem[LUT_mem_MPORT_3_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_3_data = LUT_mem_MPORT_3_addr >= 6'h23 ? _RAND_2[32:0] : LUT_mem[LUT_mem_MPORT_3_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_5_addr = 6'h1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_5_data = LUT_mem[LUT_mem_MPORT_5_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_5_data = LUT_mem_MPORT_5_addr >= 6'h23 ? _RAND_3[32:0] : LUT_mem[LUT_mem_MPORT_5_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_7_addr = 6'h1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_7_data = LUT_mem[LUT_mem_MPORT_7_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_7_data = LUT_mem_MPORT_7_addr >= 6'h23 ? _RAND_4[32:0] : LUT_mem[LUT_mem_MPORT_7_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_9_addr = 6'h2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_9_data = LUT_mem[LUT_mem_MPORT_9_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_9_data = LUT_mem_MPORT_9_addr >= 6'h23 ? _RAND_5[32:0] : LUT_mem[LUT_mem_MPORT_9_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_11_addr = 6'h2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_11_data = LUT_mem[LUT_mem_MPORT_11_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_11_data = LUT_mem_MPORT_11_addr >= 6'h23 ? _RAND_6[32:0] : LUT_mem[LUT_mem_MPORT_11_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_13_addr = 6'h3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_13_data = LUT_mem[LUT_mem_MPORT_13_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_13_data = LUT_mem_MPORT_13_addr >= 6'h23 ? _RAND_7[32:0] : LUT_mem[LUT_mem_MPORT_13_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_15_addr = 6'h3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_15_data = LUT_mem[LUT_mem_MPORT_15_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_15_data = LUT_mem_MPORT_15_addr >= 6'h23 ? _RAND_8[32:0] : LUT_mem[LUT_mem_MPORT_15_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_17_addr = 6'h4;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_17_data = LUT_mem[LUT_mem_MPORT_17_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_17_data = LUT_mem_MPORT_17_addr >= 6'h23 ? _RAND_9[32:0] : LUT_mem[LUT_mem_MPORT_17_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_19_addr = 6'h4;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_19_data = LUT_mem[LUT_mem_MPORT_19_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_19_data = LUT_mem_MPORT_19_addr >= 6'h23 ? _RAND_10[32:0] : LUT_mem[LUT_mem_MPORT_19_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_21_addr = 6'h5;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_21_data = LUT_mem[LUT_mem_MPORT_21_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_21_data = LUT_mem_MPORT_21_addr >= 6'h23 ? _RAND_11[32:0] : LUT_mem[LUT_mem_MPORT_21_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_23_addr = 6'h5;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_23_data = LUT_mem[LUT_mem_MPORT_23_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_23_data = LUT_mem_MPORT_23_addr >= 6'h23 ? _RAND_12[32:0] : LUT_mem[LUT_mem_MPORT_23_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_25_addr = 6'h6;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_25_data = LUT_mem[LUT_mem_MPORT_25_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_25_data = LUT_mem_MPORT_25_addr >= 6'h23 ? _RAND_13[32:0] : LUT_mem[LUT_mem_MPORT_25_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_27_addr = 6'h6;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_27_data = LUT_mem[LUT_mem_MPORT_27_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_27_data = LUT_mem_MPORT_27_addr >= 6'h23 ? _RAND_14[32:0] : LUT_mem[LUT_mem_MPORT_27_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_29_addr = 6'h7;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_29_data = LUT_mem[LUT_mem_MPORT_29_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_29_data = LUT_mem_MPORT_29_addr >= 6'h23 ? _RAND_15[32:0] : LUT_mem[LUT_mem_MPORT_29_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_31_addr = 6'h7;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_31_data = LUT_mem[LUT_mem_MPORT_31_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_31_data = LUT_mem_MPORT_31_addr >= 6'h23 ? _RAND_16[32:0] : LUT_mem[LUT_mem_MPORT_31_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_33_addr = 6'h8;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_33_data = LUT_mem[LUT_mem_MPORT_33_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_33_data = LUT_mem_MPORT_33_addr >= 6'h23 ? _RAND_17[32:0] : LUT_mem[LUT_mem_MPORT_33_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_35_addr = 6'h8;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_35_data = LUT_mem[LUT_mem_MPORT_35_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_35_data = LUT_mem_MPORT_35_addr >= 6'h23 ? _RAND_18[32:0] : LUT_mem[LUT_mem_MPORT_35_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_37_addr = 6'h9;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_37_data = LUT_mem[LUT_mem_MPORT_37_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_37_data = LUT_mem_MPORT_37_addr >= 6'h23 ? _RAND_19[32:0] : LUT_mem[LUT_mem_MPORT_37_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_39_addr = 6'h9;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_39_data = LUT_mem[LUT_mem_MPORT_39_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_39_data = LUT_mem_MPORT_39_addr >= 6'h23 ? _RAND_20[32:0] : LUT_mem[LUT_mem_MPORT_39_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_41_addr = 6'ha;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_41_data = LUT_mem[LUT_mem_MPORT_41_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_41_data = LUT_mem_MPORT_41_addr >= 6'h23 ? _RAND_21[32:0] : LUT_mem[LUT_mem_MPORT_41_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_43_addr = 6'ha;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_43_data = LUT_mem[LUT_mem_MPORT_43_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_43_data = LUT_mem_MPORT_43_addr >= 6'h23 ? _RAND_22[32:0] : LUT_mem[LUT_mem_MPORT_43_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_45_addr = 6'hb;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_45_data = LUT_mem[LUT_mem_MPORT_45_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_45_data = LUT_mem_MPORT_45_addr >= 6'h23 ? _RAND_23[32:0] : LUT_mem[LUT_mem_MPORT_45_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_47_addr = 6'hb;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_47_data = LUT_mem[LUT_mem_MPORT_47_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_47_data = LUT_mem_MPORT_47_addr >= 6'h23 ? _RAND_24[32:0] : LUT_mem[LUT_mem_MPORT_47_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_49_addr = 6'hc;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_49_data = LUT_mem[LUT_mem_MPORT_49_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_49_data = LUT_mem_MPORT_49_addr >= 6'h23 ? _RAND_25[32:0] : LUT_mem[LUT_mem_MPORT_49_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_51_addr = 6'hc;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_51_data = LUT_mem[LUT_mem_MPORT_51_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_51_data = LUT_mem_MPORT_51_addr >= 6'h23 ? _RAND_26[32:0] : LUT_mem[LUT_mem_MPORT_51_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_53_addr = 6'hd;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_53_data = LUT_mem[LUT_mem_MPORT_53_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_53_data = LUT_mem_MPORT_53_addr >= 6'h23 ? _RAND_27[32:0] : LUT_mem[LUT_mem_MPORT_53_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_55_addr = 6'hd;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_55_data = LUT_mem[LUT_mem_MPORT_55_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_55_data = LUT_mem_MPORT_55_addr >= 6'h23 ? _RAND_28[32:0] : LUT_mem[LUT_mem_MPORT_55_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_57_addr = 6'he;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_57_data = LUT_mem[LUT_mem_MPORT_57_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_57_data = LUT_mem_MPORT_57_addr >= 6'h23 ? _RAND_29[32:0] : LUT_mem[LUT_mem_MPORT_57_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_59_addr = 6'he;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_59_data = LUT_mem[LUT_mem_MPORT_59_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_59_data = LUT_mem_MPORT_59_addr >= 6'h23 ? _RAND_30[32:0] : LUT_mem[LUT_mem_MPORT_59_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_61_addr = 6'hf;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_61_data = LUT_mem[LUT_mem_MPORT_61_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_61_data = LUT_mem_MPORT_61_addr >= 6'h23 ? _RAND_31[32:0] : LUT_mem[LUT_mem_MPORT_61_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_63_addr = 6'hf;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_63_data = LUT_mem[LUT_mem_MPORT_63_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_63_data = LUT_mem_MPORT_63_addr >= 6'h23 ? _RAND_32[32:0] : LUT_mem[LUT_mem_MPORT_63_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_65_addr = 6'h10;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_65_data = LUT_mem[LUT_mem_MPORT_65_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_65_data = LUT_mem_MPORT_65_addr >= 6'h23 ? _RAND_33[32:0] : LUT_mem[LUT_mem_MPORT_65_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_67_addr = 6'h10;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_67_data = LUT_mem[LUT_mem_MPORT_67_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_67_data = LUT_mem_MPORT_67_addr >= 6'h23 ? _RAND_34[32:0] : LUT_mem[LUT_mem_MPORT_67_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_69_addr = 6'h11;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_69_data = LUT_mem[LUT_mem_MPORT_69_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_69_data = LUT_mem_MPORT_69_addr >= 6'h23 ? _RAND_35[32:0] : LUT_mem[LUT_mem_MPORT_69_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_71_addr = 6'h11;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_71_data = LUT_mem[LUT_mem_MPORT_71_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_71_data = LUT_mem_MPORT_71_addr >= 6'h23 ? _RAND_36[32:0] : LUT_mem[LUT_mem_MPORT_71_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_73_addr = 6'h12;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_73_data = LUT_mem[LUT_mem_MPORT_73_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_73_data = LUT_mem_MPORT_73_addr >= 6'h23 ? _RAND_37[32:0] : LUT_mem[LUT_mem_MPORT_73_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_75_addr = 6'h12;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_75_data = LUT_mem[LUT_mem_MPORT_75_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_75_data = LUT_mem_MPORT_75_addr >= 6'h23 ? _RAND_38[32:0] : LUT_mem[LUT_mem_MPORT_75_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_77_addr = 6'h13;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_77_data = LUT_mem[LUT_mem_MPORT_77_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_77_data = LUT_mem_MPORT_77_addr >= 6'h23 ? _RAND_39[32:0] : LUT_mem[LUT_mem_MPORT_77_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_79_addr = 6'h13;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_79_data = LUT_mem[LUT_mem_MPORT_79_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_79_data = LUT_mem_MPORT_79_addr >= 6'h23 ? _RAND_40[32:0] : LUT_mem[LUT_mem_MPORT_79_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_81_addr = 6'h14;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_81_data = LUT_mem[LUT_mem_MPORT_81_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_81_data = LUT_mem_MPORT_81_addr >= 6'h23 ? _RAND_41[32:0] : LUT_mem[LUT_mem_MPORT_81_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_83_addr = 6'h14;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_83_data = LUT_mem[LUT_mem_MPORT_83_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_83_data = LUT_mem_MPORT_83_addr >= 6'h23 ? _RAND_42[32:0] : LUT_mem[LUT_mem_MPORT_83_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_85_addr = 6'h15;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_85_data = LUT_mem[LUT_mem_MPORT_85_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_85_data = LUT_mem_MPORT_85_addr >= 6'h23 ? _RAND_43[32:0] : LUT_mem[LUT_mem_MPORT_85_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_87_addr = 6'h15;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_87_data = LUT_mem[LUT_mem_MPORT_87_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_87_data = LUT_mem_MPORT_87_addr >= 6'h23 ? _RAND_44[32:0] : LUT_mem[LUT_mem_MPORT_87_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_89_addr = 6'h16;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_89_data = LUT_mem[LUT_mem_MPORT_89_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_89_data = LUT_mem_MPORT_89_addr >= 6'h23 ? _RAND_45[32:0] : LUT_mem[LUT_mem_MPORT_89_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_91_addr = 6'h16;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_91_data = LUT_mem[LUT_mem_MPORT_91_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_91_data = LUT_mem_MPORT_91_addr >= 6'h23 ? _RAND_46[32:0] : LUT_mem[LUT_mem_MPORT_91_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_93_addr = 6'h17;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_93_data = LUT_mem[LUT_mem_MPORT_93_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_93_data = LUT_mem_MPORT_93_addr >= 6'h23 ? _RAND_47[32:0] : LUT_mem[LUT_mem_MPORT_93_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_95_addr = 6'h17;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_95_data = LUT_mem[LUT_mem_MPORT_95_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_95_data = LUT_mem_MPORT_95_addr >= 6'h23 ? _RAND_48[32:0] : LUT_mem[LUT_mem_MPORT_95_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_97_addr = 6'h18;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_97_data = LUT_mem[LUT_mem_MPORT_97_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_97_data = LUT_mem_MPORT_97_addr >= 6'h23 ? _RAND_49[32:0] : LUT_mem[LUT_mem_MPORT_97_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_99_addr = 6'h18;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_99_data = LUT_mem[LUT_mem_MPORT_99_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_99_data = LUT_mem_MPORT_99_addr >= 6'h23 ? _RAND_50[32:0] : LUT_mem[LUT_mem_MPORT_99_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_101_addr = 6'h19;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_101_data = LUT_mem[LUT_mem_MPORT_101_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_101_data = LUT_mem_MPORT_101_addr >= 6'h23 ? _RAND_51[32:0] : LUT_mem[LUT_mem_MPORT_101_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_103_addr = 6'h19;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_103_data = LUT_mem[LUT_mem_MPORT_103_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_103_data = LUT_mem_MPORT_103_addr >= 6'h23 ? _RAND_52[32:0] : LUT_mem[LUT_mem_MPORT_103_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_105_addr = 6'h1a;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_105_data = LUT_mem[LUT_mem_MPORT_105_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_105_data = LUT_mem_MPORT_105_addr >= 6'h23 ? _RAND_53[32:0] : LUT_mem[LUT_mem_MPORT_105_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_107_addr = 6'h1a;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_107_data = LUT_mem[LUT_mem_MPORT_107_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_107_data = LUT_mem_MPORT_107_addr >= 6'h23 ? _RAND_54[32:0] : LUT_mem[LUT_mem_MPORT_107_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_109_addr = 6'h1b;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_109_data = LUT_mem[LUT_mem_MPORT_109_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_109_data = LUT_mem_MPORT_109_addr >= 6'h23 ? _RAND_55[32:0] : LUT_mem[LUT_mem_MPORT_109_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_111_addr = 6'h1b;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_111_data = LUT_mem[LUT_mem_MPORT_111_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_111_data = LUT_mem_MPORT_111_addr >= 6'h23 ? _RAND_56[32:0] : LUT_mem[LUT_mem_MPORT_111_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_113_addr = 6'h1c;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_113_data = LUT_mem[LUT_mem_MPORT_113_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_113_data = LUT_mem_MPORT_113_addr >= 6'h23 ? _RAND_57[32:0] : LUT_mem[LUT_mem_MPORT_113_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_115_addr = 6'h1c;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_115_data = LUT_mem[LUT_mem_MPORT_115_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_115_data = LUT_mem_MPORT_115_addr >= 6'h23 ? _RAND_58[32:0] : LUT_mem[LUT_mem_MPORT_115_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_117_addr = 6'h1d;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_117_data = LUT_mem[LUT_mem_MPORT_117_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_117_data = LUT_mem_MPORT_117_addr >= 6'h23 ? _RAND_59[32:0] : LUT_mem[LUT_mem_MPORT_117_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_119_addr = 6'h1d;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_119_data = LUT_mem[LUT_mem_MPORT_119_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_119_data = LUT_mem_MPORT_119_addr >= 6'h23 ? _RAND_60[32:0] : LUT_mem[LUT_mem_MPORT_119_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_121_addr = 6'h1e;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_121_data = LUT_mem[LUT_mem_MPORT_121_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_121_data = LUT_mem_MPORT_121_addr >= 6'h23 ? _RAND_61[32:0] : LUT_mem[LUT_mem_MPORT_121_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_123_addr = 6'h1e;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_123_data = LUT_mem[LUT_mem_MPORT_123_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_123_data = LUT_mem_MPORT_123_addr >= 6'h23 ? _RAND_62[32:0] : LUT_mem[LUT_mem_MPORT_123_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_125_addr = 6'h1f;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_125_data = LUT_mem[LUT_mem_MPORT_125_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_125_data = LUT_mem_MPORT_125_addr >= 6'h23 ? _RAND_63[32:0] : LUT_mem[LUT_mem_MPORT_125_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_127_addr = 6'h1f;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_127_data = LUT_mem[LUT_mem_MPORT_127_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_127_data = LUT_mem_MPORT_127_addr >= 6'h23 ? _RAND_64[32:0] : LUT_mem[LUT_mem_MPORT_127_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_129_addr = 6'h20;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_129_data = LUT_mem[LUT_mem_MPORT_129_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_129_data = LUT_mem_MPORT_129_addr >= 6'h23 ? _RAND_65[32:0] : LUT_mem[LUT_mem_MPORT_129_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_131_addr = 6'h20;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_131_data = LUT_mem[LUT_mem_MPORT_131_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_131_data = LUT_mem_MPORT_131_addr >= 6'h23 ? _RAND_66[32:0] : LUT_mem[LUT_mem_MPORT_131_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_133_addr = 6'h21;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_133_data = LUT_mem[LUT_mem_MPORT_133_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_133_data = LUT_mem_MPORT_133_addr >= 6'h23 ? _RAND_67[32:0] : LUT_mem[LUT_mem_MPORT_133_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_135_addr = 6'h21;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_135_data = LUT_mem[LUT_mem_MPORT_135_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_135_data = LUT_mem_MPORT_135_addr >= 6'h23 ? _RAND_68[32:0] : LUT_mem[LUT_mem_MPORT_135_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_137_addr = 6'h22;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_137_data = LUT_mem[LUT_mem_MPORT_137_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_137_data = LUT_mem_MPORT_137_addr >= 6'h23 ? _RAND_69[32:0] : LUT_mem[LUT_mem_MPORT_137_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_139_addr = 6'h22;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_139_data = LUT_mem[LUT_mem_MPORT_139_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_139_data = LUT_mem_MPORT_139_addr >= 6'h23 ? _RAND_70[32:0] : LUT_mem[LUT_mem_MPORT_139_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_140_addr = 6'h0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_140_data = LUT_mem[LUT_mem_MPORT_140_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_140_data = LUT_mem_MPORT_140_addr >= 6'h23 ? _RAND_71[32:0] : LUT_mem[LUT_mem_MPORT_140_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_141_addr = 6'h1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_141_data = LUT_mem[LUT_mem_MPORT_141_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_141_data = LUT_mem_MPORT_141_addr >= 6'h23 ? _RAND_72[32:0] : LUT_mem[LUT_mem_MPORT_141_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_142_addr = 6'h2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_142_data = LUT_mem[LUT_mem_MPORT_142_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_142_data = LUT_mem_MPORT_142_addr >= 6'h23 ? _RAND_73[32:0] : LUT_mem[LUT_mem_MPORT_142_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_143_addr = 6'h3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_143_data = LUT_mem[LUT_mem_MPORT_143_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_143_data = LUT_mem_MPORT_143_addr >= 6'h23 ? _RAND_74[32:0] : LUT_mem[LUT_mem_MPORT_143_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_144_addr = 6'h4;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_144_data = LUT_mem[LUT_mem_MPORT_144_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_144_data = LUT_mem_MPORT_144_addr >= 6'h23 ? _RAND_75[32:0] : LUT_mem[LUT_mem_MPORT_144_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_145_addr = 6'h5;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_145_data = LUT_mem[LUT_mem_MPORT_145_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_145_data = LUT_mem_MPORT_145_addr >= 6'h23 ? _RAND_76[32:0] : LUT_mem[LUT_mem_MPORT_145_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_146_addr = 6'h6;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_146_data = LUT_mem[LUT_mem_MPORT_146_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_146_data = LUT_mem_MPORT_146_addr >= 6'h23 ? _RAND_77[32:0] : LUT_mem[LUT_mem_MPORT_146_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_147_addr = 6'h7;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_147_data = LUT_mem[LUT_mem_MPORT_147_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_147_data = LUT_mem_MPORT_147_addr >= 6'h23 ? _RAND_78[32:0] : LUT_mem[LUT_mem_MPORT_147_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_148_addr = 6'h8;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_148_data = LUT_mem[LUT_mem_MPORT_148_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_148_data = LUT_mem_MPORT_148_addr >= 6'h23 ? _RAND_79[32:0] : LUT_mem[LUT_mem_MPORT_148_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_149_addr = 6'h9;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_149_data = LUT_mem[LUT_mem_MPORT_149_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_149_data = LUT_mem_MPORT_149_addr >= 6'h23 ? _RAND_80[32:0] : LUT_mem[LUT_mem_MPORT_149_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_150_addr = 6'ha;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_150_data = LUT_mem[LUT_mem_MPORT_150_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_150_data = LUT_mem_MPORT_150_addr >= 6'h23 ? _RAND_81[32:0] : LUT_mem[LUT_mem_MPORT_150_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_151_addr = 6'hb;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_151_data = LUT_mem[LUT_mem_MPORT_151_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_151_data = LUT_mem_MPORT_151_addr >= 6'h23 ? _RAND_82[32:0] : LUT_mem[LUT_mem_MPORT_151_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_152_addr = 6'hc;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_152_data = LUT_mem[LUT_mem_MPORT_152_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_152_data = LUT_mem_MPORT_152_addr >= 6'h23 ? _RAND_83[32:0] : LUT_mem[LUT_mem_MPORT_152_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_153_addr = 6'hd;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_153_data = LUT_mem[LUT_mem_MPORT_153_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_153_data = LUT_mem_MPORT_153_addr >= 6'h23 ? _RAND_84[32:0] : LUT_mem[LUT_mem_MPORT_153_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_154_addr = 6'he;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_154_data = LUT_mem[LUT_mem_MPORT_154_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_154_data = LUT_mem_MPORT_154_addr >= 6'h23 ? _RAND_85[32:0] : LUT_mem[LUT_mem_MPORT_154_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_155_addr = 6'hf;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_155_data = LUT_mem[LUT_mem_MPORT_155_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_155_data = LUT_mem_MPORT_155_addr >= 6'h23 ? _RAND_86[32:0] : LUT_mem[LUT_mem_MPORT_155_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_156_addr = 6'h10;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_156_data = LUT_mem[LUT_mem_MPORT_156_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_156_data = LUT_mem_MPORT_156_addr >= 6'h23 ? _RAND_87[32:0] : LUT_mem[LUT_mem_MPORT_156_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_157_addr = 6'h11;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_157_data = LUT_mem[LUT_mem_MPORT_157_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_157_data = LUT_mem_MPORT_157_addr >= 6'h23 ? _RAND_88[32:0] : LUT_mem[LUT_mem_MPORT_157_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_158_addr = 6'h12;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_158_data = LUT_mem[LUT_mem_MPORT_158_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_158_data = LUT_mem_MPORT_158_addr >= 6'h23 ? _RAND_89[32:0] : LUT_mem[LUT_mem_MPORT_158_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_159_addr = 6'h13;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_159_data = LUT_mem[LUT_mem_MPORT_159_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_159_data = LUT_mem_MPORT_159_addr >= 6'h23 ? _RAND_90[32:0] : LUT_mem[LUT_mem_MPORT_159_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_160_addr = 6'h14;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_160_data = LUT_mem[LUT_mem_MPORT_160_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_160_data = LUT_mem_MPORT_160_addr >= 6'h23 ? _RAND_91[32:0] : LUT_mem[LUT_mem_MPORT_160_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_161_addr = 6'h15;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_161_data = LUT_mem[LUT_mem_MPORT_161_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_161_data = LUT_mem_MPORT_161_addr >= 6'h23 ? _RAND_92[32:0] : LUT_mem[LUT_mem_MPORT_161_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_162_addr = 6'h16;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_162_data = LUT_mem[LUT_mem_MPORT_162_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_162_data = LUT_mem_MPORT_162_addr >= 6'h23 ? _RAND_93[32:0] : LUT_mem[LUT_mem_MPORT_162_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_163_addr = 6'h17;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_163_data = LUT_mem[LUT_mem_MPORT_163_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_163_data = LUT_mem_MPORT_163_addr >= 6'h23 ? _RAND_94[32:0] : LUT_mem[LUT_mem_MPORT_163_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_164_addr = 6'h18;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_164_data = LUT_mem[LUT_mem_MPORT_164_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_164_data = LUT_mem_MPORT_164_addr >= 6'h23 ? _RAND_95[32:0] : LUT_mem[LUT_mem_MPORT_164_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_165_addr = 6'h19;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_165_data = LUT_mem[LUT_mem_MPORT_165_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_165_data = LUT_mem_MPORT_165_addr >= 6'h23 ? _RAND_96[32:0] : LUT_mem[LUT_mem_MPORT_165_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_166_addr = 6'h1a;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_166_data = LUT_mem[LUT_mem_MPORT_166_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_166_data = LUT_mem_MPORT_166_addr >= 6'h23 ? _RAND_97[32:0] : LUT_mem[LUT_mem_MPORT_166_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_167_addr = 6'h1b;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_167_data = LUT_mem[LUT_mem_MPORT_167_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_167_data = LUT_mem_MPORT_167_addr >= 6'h23 ? _RAND_98[32:0] : LUT_mem[LUT_mem_MPORT_167_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_168_addr = 6'h1c;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_168_data = LUT_mem[LUT_mem_MPORT_168_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_168_data = LUT_mem_MPORT_168_addr >= 6'h23 ? _RAND_99[32:0] : LUT_mem[LUT_mem_MPORT_168_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_169_addr = 6'h1d;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_169_data = LUT_mem[LUT_mem_MPORT_169_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_169_data = LUT_mem_MPORT_169_addr >= 6'h23 ? _RAND_100[32:0] : LUT_mem[LUT_mem_MPORT_169_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_170_addr = 6'h1e;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_170_data = LUT_mem[LUT_mem_MPORT_170_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_170_data = LUT_mem_MPORT_170_addr >= 6'h23 ? _RAND_101[32:0] : LUT_mem[LUT_mem_MPORT_170_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_171_addr = 6'h1f;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_171_data = LUT_mem[LUT_mem_MPORT_171_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_171_data = LUT_mem_MPORT_171_addr >= 6'h23 ? _RAND_102[32:0] : LUT_mem[LUT_mem_MPORT_171_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_172_addr = 6'h20;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_172_data = LUT_mem[LUT_mem_MPORT_172_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_172_data = LUT_mem_MPORT_172_addr >= 6'h23 ? _RAND_103[32:0] : LUT_mem[LUT_mem_MPORT_172_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_173_addr = 6'h21;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_173_data = LUT_mem[LUT_mem_MPORT_173_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_173_data = LUT_mem_MPORT_173_addr >= 6'h23 ? _RAND_104[32:0] : LUT_mem[LUT_mem_MPORT_173_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_174_addr = 6'h22;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_174_data = LUT_mem[LUT_mem_MPORT_174_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_174_data = LUT_mem_MPORT_174_addr >= 6'h23 ? _RAND_105[32:0] : LUT_mem[LUT_mem_MPORT_174_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_175_addr = 6'h0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_175_data = LUT_mem[LUT_mem_MPORT_175_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_175_data = LUT_mem_MPORT_175_addr >= 6'h23 ? _RAND_106[32:0] : LUT_mem[LUT_mem_MPORT_175_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_176_addr = 6'h1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_176_data = LUT_mem[LUT_mem_MPORT_176_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_176_data = LUT_mem_MPORT_176_addr >= 6'h23 ? _RAND_107[32:0] : LUT_mem[LUT_mem_MPORT_176_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_177_addr = 6'h2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_177_data = LUT_mem[LUT_mem_MPORT_177_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_177_data = LUT_mem_MPORT_177_addr >= 6'h23 ? _RAND_108[32:0] : LUT_mem[LUT_mem_MPORT_177_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_178_addr = 6'h3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_178_data = LUT_mem[LUT_mem_MPORT_178_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_178_data = LUT_mem_MPORT_178_addr >= 6'h23 ? _RAND_109[32:0] : LUT_mem[LUT_mem_MPORT_178_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_179_addr = 6'h4;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_179_data = LUT_mem[LUT_mem_MPORT_179_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_179_data = LUT_mem_MPORT_179_addr >= 6'h23 ? _RAND_110[32:0] : LUT_mem[LUT_mem_MPORT_179_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_180_addr = 6'h5;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_180_data = LUT_mem[LUT_mem_MPORT_180_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_180_data = LUT_mem_MPORT_180_addr >= 6'h23 ? _RAND_111[32:0] : LUT_mem[LUT_mem_MPORT_180_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_181_addr = 6'h6;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_181_data = LUT_mem[LUT_mem_MPORT_181_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_181_data = LUT_mem_MPORT_181_addr >= 6'h23 ? _RAND_112[32:0] : LUT_mem[LUT_mem_MPORT_181_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_182_addr = 6'h7;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_182_data = LUT_mem[LUT_mem_MPORT_182_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_182_data = LUT_mem_MPORT_182_addr >= 6'h23 ? _RAND_113[32:0] : LUT_mem[LUT_mem_MPORT_182_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_183_addr = 6'h8;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_183_data = LUT_mem[LUT_mem_MPORT_183_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_183_data = LUT_mem_MPORT_183_addr >= 6'h23 ? _RAND_114[32:0] : LUT_mem[LUT_mem_MPORT_183_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_184_addr = 6'h9;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_184_data = LUT_mem[LUT_mem_MPORT_184_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_184_data = LUT_mem_MPORT_184_addr >= 6'h23 ? _RAND_115[32:0] : LUT_mem[LUT_mem_MPORT_184_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_185_addr = 6'ha;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_185_data = LUT_mem[LUT_mem_MPORT_185_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_185_data = LUT_mem_MPORT_185_addr >= 6'h23 ? _RAND_116[32:0] : LUT_mem[LUT_mem_MPORT_185_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_186_addr = 6'hb;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_186_data = LUT_mem[LUT_mem_MPORT_186_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_186_data = LUT_mem_MPORT_186_addr >= 6'h23 ? _RAND_117[32:0] : LUT_mem[LUT_mem_MPORT_186_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_187_addr = 6'hc;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_187_data = LUT_mem[LUT_mem_MPORT_187_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_187_data = LUT_mem_MPORT_187_addr >= 6'h23 ? _RAND_118[32:0] : LUT_mem[LUT_mem_MPORT_187_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_188_addr = 6'hd;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_188_data = LUT_mem[LUT_mem_MPORT_188_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_188_data = LUT_mem_MPORT_188_addr >= 6'h23 ? _RAND_119[32:0] : LUT_mem[LUT_mem_MPORT_188_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_189_addr = 6'he;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_189_data = LUT_mem[LUT_mem_MPORT_189_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_189_data = LUT_mem_MPORT_189_addr >= 6'h23 ? _RAND_120[32:0] : LUT_mem[LUT_mem_MPORT_189_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_190_addr = 6'hf;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_190_data = LUT_mem[LUT_mem_MPORT_190_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_190_data = LUT_mem_MPORT_190_addr >= 6'h23 ? _RAND_121[32:0] : LUT_mem[LUT_mem_MPORT_190_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_191_addr = 6'h10;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_191_data = LUT_mem[LUT_mem_MPORT_191_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_191_data = LUT_mem_MPORT_191_addr >= 6'h23 ? _RAND_122[32:0] : LUT_mem[LUT_mem_MPORT_191_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_192_addr = 6'h11;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_192_data = LUT_mem[LUT_mem_MPORT_192_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_192_data = LUT_mem_MPORT_192_addr >= 6'h23 ? _RAND_123[32:0] : LUT_mem[LUT_mem_MPORT_192_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_193_addr = 6'h12;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_193_data = LUT_mem[LUT_mem_MPORT_193_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_193_data = LUT_mem_MPORT_193_addr >= 6'h23 ? _RAND_124[32:0] : LUT_mem[LUT_mem_MPORT_193_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_194_addr = 6'h13;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_194_data = LUT_mem[LUT_mem_MPORT_194_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_194_data = LUT_mem_MPORT_194_addr >= 6'h23 ? _RAND_125[32:0] : LUT_mem[LUT_mem_MPORT_194_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_195_addr = 6'h14;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_195_data = LUT_mem[LUT_mem_MPORT_195_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_195_data = LUT_mem_MPORT_195_addr >= 6'h23 ? _RAND_126[32:0] : LUT_mem[LUT_mem_MPORT_195_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_196_addr = 6'h15;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_196_data = LUT_mem[LUT_mem_MPORT_196_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_196_data = LUT_mem_MPORT_196_addr >= 6'h23 ? _RAND_127[32:0] : LUT_mem[LUT_mem_MPORT_196_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_197_addr = 6'h16;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_197_data = LUT_mem[LUT_mem_MPORT_197_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_197_data = LUT_mem_MPORT_197_addr >= 6'h23 ? _RAND_128[32:0] : LUT_mem[LUT_mem_MPORT_197_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_198_addr = 6'h17;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_198_data = LUT_mem[LUT_mem_MPORT_198_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_198_data = LUT_mem_MPORT_198_addr >= 6'h23 ? _RAND_129[32:0] : LUT_mem[LUT_mem_MPORT_198_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_199_addr = 6'h18;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_199_data = LUT_mem[LUT_mem_MPORT_199_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_199_data = LUT_mem_MPORT_199_addr >= 6'h23 ? _RAND_130[32:0] : LUT_mem[LUT_mem_MPORT_199_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_200_addr = 6'h19;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_200_data = LUT_mem[LUT_mem_MPORT_200_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_200_data = LUT_mem_MPORT_200_addr >= 6'h23 ? _RAND_131[32:0] : LUT_mem[LUT_mem_MPORT_200_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_201_addr = 6'h1a;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_201_data = LUT_mem[LUT_mem_MPORT_201_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_201_data = LUT_mem_MPORT_201_addr >= 6'h23 ? _RAND_132[32:0] : LUT_mem[LUT_mem_MPORT_201_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_202_addr = 6'h1b;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_202_data = LUT_mem[LUT_mem_MPORT_202_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_202_data = LUT_mem_MPORT_202_addr >= 6'h23 ? _RAND_133[32:0] : LUT_mem[LUT_mem_MPORT_202_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_203_addr = 6'h1c;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_203_data = LUT_mem[LUT_mem_MPORT_203_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_203_data = LUT_mem_MPORT_203_addr >= 6'h23 ? _RAND_134[32:0] : LUT_mem[LUT_mem_MPORT_203_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_204_addr = 6'h1d;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_204_data = LUT_mem[LUT_mem_MPORT_204_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_204_data = LUT_mem_MPORT_204_addr >= 6'h23 ? _RAND_135[32:0] : LUT_mem[LUT_mem_MPORT_204_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_205_addr = 6'h1e;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_205_data = LUT_mem[LUT_mem_MPORT_205_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_205_data = LUT_mem_MPORT_205_addr >= 6'h23 ? _RAND_136[32:0] : LUT_mem[LUT_mem_MPORT_205_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_206_addr = 6'h1f;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_206_data = LUT_mem[LUT_mem_MPORT_206_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_206_data = LUT_mem_MPORT_206_addr >= 6'h23 ? _RAND_137[32:0] : LUT_mem[LUT_mem_MPORT_206_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_207_addr = 6'h20;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_207_data = LUT_mem[LUT_mem_MPORT_207_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_207_data = LUT_mem_MPORT_207_addr >= 6'h23 ? _RAND_138[32:0] : LUT_mem[LUT_mem_MPORT_207_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_208_addr = 6'h21;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_208_data = LUT_mem[LUT_mem_MPORT_208_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_208_data = LUT_mem_MPORT_208_addr >= 6'h23 ? _RAND_139[32:0] : LUT_mem[LUT_mem_MPORT_208_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_209_addr = 6'h22;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_209_data = LUT_mem[LUT_mem_MPORT_209_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_209_data = LUT_mem_MPORT_209_addr >= 6'h23 ? _RAND_140[32:0] : LUT_mem[LUT_mem_MPORT_209_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_210_addr = 6'h0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_210_data = LUT_mem[LUT_mem_MPORT_210_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_210_data = LUT_mem_MPORT_210_addr >= 6'h23 ? _RAND_141[32:0] : LUT_mem[LUT_mem_MPORT_210_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_212_addr = 6'h1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_212_data = LUT_mem[LUT_mem_MPORT_212_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_212_data = LUT_mem_MPORT_212_addr >= 6'h23 ? _RAND_142[32:0] : LUT_mem[LUT_mem_MPORT_212_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_214_addr = 6'h2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_214_data = LUT_mem[LUT_mem_MPORT_214_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_214_data = LUT_mem_MPORT_214_addr >= 6'h23 ? _RAND_143[32:0] : LUT_mem[LUT_mem_MPORT_214_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_216_addr = 6'h3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_216_data = LUT_mem[LUT_mem_MPORT_216_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_216_data = LUT_mem_MPORT_216_addr >= 6'h23 ? _RAND_144[32:0] : LUT_mem[LUT_mem_MPORT_216_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_218_addr = 6'h4;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_218_data = LUT_mem[LUT_mem_MPORT_218_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_218_data = LUT_mem_MPORT_218_addr >= 6'h23 ? _RAND_145[32:0] : LUT_mem[LUT_mem_MPORT_218_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_220_addr = 6'h5;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_220_data = LUT_mem[LUT_mem_MPORT_220_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_220_data = LUT_mem_MPORT_220_addr >= 6'h23 ? _RAND_146[32:0] : LUT_mem[LUT_mem_MPORT_220_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_222_addr = 6'h6;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_222_data = LUT_mem[LUT_mem_MPORT_222_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_222_data = LUT_mem_MPORT_222_addr >= 6'h23 ? _RAND_147[32:0] : LUT_mem[LUT_mem_MPORT_222_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_224_addr = 6'h7;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_224_data = LUT_mem[LUT_mem_MPORT_224_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_224_data = LUT_mem_MPORT_224_addr >= 6'h23 ? _RAND_148[32:0] : LUT_mem[LUT_mem_MPORT_224_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_226_addr = 6'h8;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_226_data = LUT_mem[LUT_mem_MPORT_226_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_226_data = LUT_mem_MPORT_226_addr >= 6'h23 ? _RAND_149[32:0] : LUT_mem[LUT_mem_MPORT_226_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_228_addr = 6'h9;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_228_data = LUT_mem[LUT_mem_MPORT_228_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_228_data = LUT_mem_MPORT_228_addr >= 6'h23 ? _RAND_150[32:0] : LUT_mem[LUT_mem_MPORT_228_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_230_addr = 6'ha;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_230_data = LUT_mem[LUT_mem_MPORT_230_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_230_data = LUT_mem_MPORT_230_addr >= 6'h23 ? _RAND_151[32:0] : LUT_mem[LUT_mem_MPORT_230_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_232_addr = 6'hb;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_232_data = LUT_mem[LUT_mem_MPORT_232_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_232_data = LUT_mem_MPORT_232_addr >= 6'h23 ? _RAND_152[32:0] : LUT_mem[LUT_mem_MPORT_232_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_234_addr = 6'hc;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_234_data = LUT_mem[LUT_mem_MPORT_234_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_234_data = LUT_mem_MPORT_234_addr >= 6'h23 ? _RAND_153[32:0] : LUT_mem[LUT_mem_MPORT_234_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_236_addr = 6'hd;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_236_data = LUT_mem[LUT_mem_MPORT_236_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_236_data = LUT_mem_MPORT_236_addr >= 6'h23 ? _RAND_154[32:0] : LUT_mem[LUT_mem_MPORT_236_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_238_addr = 6'he;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_238_data = LUT_mem[LUT_mem_MPORT_238_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_238_data = LUT_mem_MPORT_238_addr >= 6'h23 ? _RAND_155[32:0] : LUT_mem[LUT_mem_MPORT_238_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_240_addr = 6'hf;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_240_data = LUT_mem[LUT_mem_MPORT_240_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_240_data = LUT_mem_MPORT_240_addr >= 6'h23 ? _RAND_156[32:0] : LUT_mem[LUT_mem_MPORT_240_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_242_addr = 6'h10;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_242_data = LUT_mem[LUT_mem_MPORT_242_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_242_data = LUT_mem_MPORT_242_addr >= 6'h23 ? _RAND_157[32:0] : LUT_mem[LUT_mem_MPORT_242_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_244_addr = 6'h11;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_244_data = LUT_mem[LUT_mem_MPORT_244_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_244_data = LUT_mem_MPORT_244_addr >= 6'h23 ? _RAND_158[32:0] : LUT_mem[LUT_mem_MPORT_244_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_246_addr = 6'h12;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_246_data = LUT_mem[LUT_mem_MPORT_246_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_246_data = LUT_mem_MPORT_246_addr >= 6'h23 ? _RAND_159[32:0] : LUT_mem[LUT_mem_MPORT_246_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_248_addr = 6'h13;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_248_data = LUT_mem[LUT_mem_MPORT_248_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_248_data = LUT_mem_MPORT_248_addr >= 6'h23 ? _RAND_160[32:0] : LUT_mem[LUT_mem_MPORT_248_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_250_addr = 6'h14;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_250_data = LUT_mem[LUT_mem_MPORT_250_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_250_data = LUT_mem_MPORT_250_addr >= 6'h23 ? _RAND_161[32:0] : LUT_mem[LUT_mem_MPORT_250_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_252_addr = 6'h15;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_252_data = LUT_mem[LUT_mem_MPORT_252_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_252_data = LUT_mem_MPORT_252_addr >= 6'h23 ? _RAND_162[32:0] : LUT_mem[LUT_mem_MPORT_252_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_254_addr = 6'h16;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_254_data = LUT_mem[LUT_mem_MPORT_254_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_254_data = LUT_mem_MPORT_254_addr >= 6'h23 ? _RAND_163[32:0] : LUT_mem[LUT_mem_MPORT_254_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_256_addr = 6'h17;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_256_data = LUT_mem[LUT_mem_MPORT_256_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_256_data = LUT_mem_MPORT_256_addr >= 6'h23 ? _RAND_164[32:0] : LUT_mem[LUT_mem_MPORT_256_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_258_addr = 6'h18;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_258_data = LUT_mem[LUT_mem_MPORT_258_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_258_data = LUT_mem_MPORT_258_addr >= 6'h23 ? _RAND_165[32:0] : LUT_mem[LUT_mem_MPORT_258_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_260_addr = 6'h19;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_260_data = LUT_mem[LUT_mem_MPORT_260_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_260_data = LUT_mem_MPORT_260_addr >= 6'h23 ? _RAND_166[32:0] : LUT_mem[LUT_mem_MPORT_260_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_262_addr = 6'h1a;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_262_data = LUT_mem[LUT_mem_MPORT_262_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_262_data = LUT_mem_MPORT_262_addr >= 6'h23 ? _RAND_167[32:0] : LUT_mem[LUT_mem_MPORT_262_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_264_addr = 6'h1b;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_264_data = LUT_mem[LUT_mem_MPORT_264_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_264_data = LUT_mem_MPORT_264_addr >= 6'h23 ? _RAND_168[32:0] : LUT_mem[LUT_mem_MPORT_264_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_266_addr = 6'h1c;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_266_data = LUT_mem[LUT_mem_MPORT_266_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_266_data = LUT_mem_MPORT_266_addr >= 6'h23 ? _RAND_169[32:0] : LUT_mem[LUT_mem_MPORT_266_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_268_addr = 6'h1d;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_268_data = LUT_mem[LUT_mem_MPORT_268_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_268_data = LUT_mem_MPORT_268_addr >= 6'h23 ? _RAND_170[32:0] : LUT_mem[LUT_mem_MPORT_268_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_270_addr = 6'h1e;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_270_data = LUT_mem[LUT_mem_MPORT_270_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_270_data = LUT_mem_MPORT_270_addr >= 6'h23 ? _RAND_171[32:0] : LUT_mem[LUT_mem_MPORT_270_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_272_addr = 6'h1f;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_272_data = LUT_mem[LUT_mem_MPORT_272_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_272_data = LUT_mem_MPORT_272_addr >= 6'h23 ? _RAND_172[32:0] : LUT_mem[LUT_mem_MPORT_272_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_274_addr = 6'h20;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_274_data = LUT_mem[LUT_mem_MPORT_274_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_274_data = LUT_mem_MPORT_274_addr >= 6'h23 ? _RAND_173[32:0] : LUT_mem[LUT_mem_MPORT_274_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_276_addr = 6'h21;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_276_data = LUT_mem[LUT_mem_MPORT_276_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_276_data = LUT_mem_MPORT_276_addr >= 6'h23 ? _RAND_174[32:0] : LUT_mem[LUT_mem_MPORT_276_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_278_addr = 6'h22;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_278_data = LUT_mem[LUT_mem_MPORT_278_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_278_data = LUT_mem_MPORT_278_addr >= 6'h23 ? _RAND_175[32:0] : LUT_mem[LUT_mem_MPORT_278_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_280_addr = 6'h0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_280_data = LUT_mem[LUT_mem_MPORT_280_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_280_data = LUT_mem_MPORT_280_addr >= 6'h23 ? _RAND_176[32:0] : LUT_mem[LUT_mem_MPORT_280_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_281_addr = 6'h1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_281_data = LUT_mem[LUT_mem_MPORT_281_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_281_data = LUT_mem_MPORT_281_addr >= 6'h23 ? _RAND_177[32:0] : LUT_mem[LUT_mem_MPORT_281_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_282_addr = 6'h2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_282_data = LUT_mem[LUT_mem_MPORT_282_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_282_data = LUT_mem_MPORT_282_addr >= 6'h23 ? _RAND_178[32:0] : LUT_mem[LUT_mem_MPORT_282_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_283_addr = 6'h3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_283_data = LUT_mem[LUT_mem_MPORT_283_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_283_data = LUT_mem_MPORT_283_addr >= 6'h23 ? _RAND_179[32:0] : LUT_mem[LUT_mem_MPORT_283_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_284_addr = 6'h4;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_284_data = LUT_mem[LUT_mem_MPORT_284_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_284_data = LUT_mem_MPORT_284_addr >= 6'h23 ? _RAND_180[32:0] : LUT_mem[LUT_mem_MPORT_284_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_285_addr = 6'h5;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_285_data = LUT_mem[LUT_mem_MPORT_285_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_285_data = LUT_mem_MPORT_285_addr >= 6'h23 ? _RAND_181[32:0] : LUT_mem[LUT_mem_MPORT_285_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_286_addr = 6'h6;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_286_data = LUT_mem[LUT_mem_MPORT_286_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_286_data = LUT_mem_MPORT_286_addr >= 6'h23 ? _RAND_182[32:0] : LUT_mem[LUT_mem_MPORT_286_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_287_addr = 6'h7;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_287_data = LUT_mem[LUT_mem_MPORT_287_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_287_data = LUT_mem_MPORT_287_addr >= 6'h23 ? _RAND_183[32:0] : LUT_mem[LUT_mem_MPORT_287_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_288_addr = 6'h8;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_288_data = LUT_mem[LUT_mem_MPORT_288_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_288_data = LUT_mem_MPORT_288_addr >= 6'h23 ? _RAND_184[32:0] : LUT_mem[LUT_mem_MPORT_288_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_289_addr = 6'h9;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_289_data = LUT_mem[LUT_mem_MPORT_289_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_289_data = LUT_mem_MPORT_289_addr >= 6'h23 ? _RAND_185[32:0] : LUT_mem[LUT_mem_MPORT_289_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_290_addr = 6'ha;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_290_data = LUT_mem[LUT_mem_MPORT_290_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_290_data = LUT_mem_MPORT_290_addr >= 6'h23 ? _RAND_186[32:0] : LUT_mem[LUT_mem_MPORT_290_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_291_addr = 6'hb;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_291_data = LUT_mem[LUT_mem_MPORT_291_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_291_data = LUT_mem_MPORT_291_addr >= 6'h23 ? _RAND_187[32:0] : LUT_mem[LUT_mem_MPORT_291_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_292_addr = 6'hc;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_292_data = LUT_mem[LUT_mem_MPORT_292_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_292_data = LUT_mem_MPORT_292_addr >= 6'h23 ? _RAND_188[32:0] : LUT_mem[LUT_mem_MPORT_292_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_293_addr = 6'hd;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_293_data = LUT_mem[LUT_mem_MPORT_293_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_293_data = LUT_mem_MPORT_293_addr >= 6'h23 ? _RAND_189[32:0] : LUT_mem[LUT_mem_MPORT_293_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_294_addr = 6'he;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_294_data = LUT_mem[LUT_mem_MPORT_294_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_294_data = LUT_mem_MPORT_294_addr >= 6'h23 ? _RAND_190[32:0] : LUT_mem[LUT_mem_MPORT_294_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_295_addr = 6'hf;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_295_data = LUT_mem[LUT_mem_MPORT_295_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_295_data = LUT_mem_MPORT_295_addr >= 6'h23 ? _RAND_191[32:0] : LUT_mem[LUT_mem_MPORT_295_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_296_addr = 6'h10;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_296_data = LUT_mem[LUT_mem_MPORT_296_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_296_data = LUT_mem_MPORT_296_addr >= 6'h23 ? _RAND_192[32:0] : LUT_mem[LUT_mem_MPORT_296_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_297_addr = 6'h11;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_297_data = LUT_mem[LUT_mem_MPORT_297_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_297_data = LUT_mem_MPORT_297_addr >= 6'h23 ? _RAND_193[32:0] : LUT_mem[LUT_mem_MPORT_297_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_298_addr = 6'h12;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_298_data = LUT_mem[LUT_mem_MPORT_298_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_298_data = LUT_mem_MPORT_298_addr >= 6'h23 ? _RAND_194[32:0] : LUT_mem[LUT_mem_MPORT_298_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_299_addr = 6'h13;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_299_data = LUT_mem[LUT_mem_MPORT_299_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_299_data = LUT_mem_MPORT_299_addr >= 6'h23 ? _RAND_195[32:0] : LUT_mem[LUT_mem_MPORT_299_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_300_addr = 6'h14;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_300_data = LUT_mem[LUT_mem_MPORT_300_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_300_data = LUT_mem_MPORT_300_addr >= 6'h23 ? _RAND_196[32:0] : LUT_mem[LUT_mem_MPORT_300_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_301_addr = 6'h15;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_301_data = LUT_mem[LUT_mem_MPORT_301_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_301_data = LUT_mem_MPORT_301_addr >= 6'h23 ? _RAND_197[32:0] : LUT_mem[LUT_mem_MPORT_301_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_302_addr = 6'h16;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_302_data = LUT_mem[LUT_mem_MPORT_302_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_302_data = LUT_mem_MPORT_302_addr >= 6'h23 ? _RAND_198[32:0] : LUT_mem[LUT_mem_MPORT_302_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_303_addr = 6'h17;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_303_data = LUT_mem[LUT_mem_MPORT_303_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_303_data = LUT_mem_MPORT_303_addr >= 6'h23 ? _RAND_199[32:0] : LUT_mem[LUT_mem_MPORT_303_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_304_addr = 6'h18;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_304_data = LUT_mem[LUT_mem_MPORT_304_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_304_data = LUT_mem_MPORT_304_addr >= 6'h23 ? _RAND_200[32:0] : LUT_mem[LUT_mem_MPORT_304_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_305_addr = 6'h19;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_305_data = LUT_mem[LUT_mem_MPORT_305_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_305_data = LUT_mem_MPORT_305_addr >= 6'h23 ? _RAND_201[32:0] : LUT_mem[LUT_mem_MPORT_305_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_306_addr = 6'h1a;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_306_data = LUT_mem[LUT_mem_MPORT_306_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_306_data = LUT_mem_MPORT_306_addr >= 6'h23 ? _RAND_202[32:0] : LUT_mem[LUT_mem_MPORT_306_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_307_addr = 6'h1b;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_307_data = LUT_mem[LUT_mem_MPORT_307_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_307_data = LUT_mem_MPORT_307_addr >= 6'h23 ? _RAND_203[32:0] : LUT_mem[LUT_mem_MPORT_307_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_308_addr = 6'h1c;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_308_data = LUT_mem[LUT_mem_MPORT_308_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_308_data = LUT_mem_MPORT_308_addr >= 6'h23 ? _RAND_204[32:0] : LUT_mem[LUT_mem_MPORT_308_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_309_addr = 6'h1d;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_309_data = LUT_mem[LUT_mem_MPORT_309_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_309_data = LUT_mem_MPORT_309_addr >= 6'h23 ? _RAND_205[32:0] : LUT_mem[LUT_mem_MPORT_309_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_310_addr = 6'h1e;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_310_data = LUT_mem[LUT_mem_MPORT_310_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_310_data = LUT_mem_MPORT_310_addr >= 6'h23 ? _RAND_206[32:0] : LUT_mem[LUT_mem_MPORT_310_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_311_addr = 6'h1f;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_311_data = LUT_mem[LUT_mem_MPORT_311_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_311_data = LUT_mem_MPORT_311_addr >= 6'h23 ? _RAND_207[32:0] : LUT_mem[LUT_mem_MPORT_311_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_312_addr = 6'h20;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_312_data = LUT_mem[LUT_mem_MPORT_312_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_312_data = LUT_mem_MPORT_312_addr >= 6'h23 ? _RAND_208[32:0] : LUT_mem[LUT_mem_MPORT_312_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_313_addr = 6'h21;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_313_data = LUT_mem[LUT_mem_MPORT_313_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_313_data = LUT_mem_MPORT_313_addr >= 6'h23 ? _RAND_209[32:0] : LUT_mem[LUT_mem_MPORT_313_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_314_addr = 6'h22;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_314_data = LUT_mem[LUT_mem_MPORT_314_addr]; // @[lut_35.scala 177:26]
  `else
  assign LUT_mem_MPORT_314_data = LUT_mem_MPORT_314_addr >= 6'h23 ? _RAND_210[32:0] : LUT_mem[LUT_mem_MPORT_314_addr]; // @[lut_35.scala 177:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign LUT_mem_MPORT_data = {1'h0,lo};
  assign LUT_mem_MPORT_addr = 6'h0;
  assign LUT_mem_MPORT_mask = 1'h1;
  assign LUT_mem_MPORT_en = io_dispatch_0;
  assign LUT_mem_MPORT_2_data = LUT_mem_MPORT_3_data;
  assign LUT_mem_MPORT_2_addr = 6'h0;
  assign LUT_mem_MPORT_2_mask = 1'h1;
  assign LUT_mem_MPORT_2_en = io_dispatch_0 ? 1'h0 : 1'h1;
  assign LUT_mem_MPORT_4_data = {1'h0,lo_1};
  assign LUT_mem_MPORT_4_addr = 6'h1;
  assign LUT_mem_MPORT_4_mask = 1'h1;
  assign LUT_mem_MPORT_4_en = io_dispatch_1;
  assign LUT_mem_MPORT_6_data = LUT_mem_MPORT_7_data;
  assign LUT_mem_MPORT_6_addr = 6'h1;
  assign LUT_mem_MPORT_6_mask = 1'h1;
  assign LUT_mem_MPORT_6_en = io_dispatch_1 ? 1'h0 : 1'h1;
  assign LUT_mem_MPORT_8_data = {1'h0,lo_2};
  assign LUT_mem_MPORT_8_addr = 6'h2;
  assign LUT_mem_MPORT_8_mask = 1'h1;
  assign LUT_mem_MPORT_8_en = io_dispatch_2;
  assign LUT_mem_MPORT_10_data = LUT_mem_MPORT_11_data;
  assign LUT_mem_MPORT_10_addr = 6'h2;
  assign LUT_mem_MPORT_10_mask = 1'h1;
  assign LUT_mem_MPORT_10_en = io_dispatch_2 ? 1'h0 : 1'h1;
  assign LUT_mem_MPORT_12_data = {1'h0,lo_3};
  assign LUT_mem_MPORT_12_addr = 6'h3;
  assign LUT_mem_MPORT_12_mask = 1'h1;
  assign LUT_mem_MPORT_12_en = io_dispatch_3;
  assign LUT_mem_MPORT_14_data = LUT_mem_MPORT_15_data;
  assign LUT_mem_MPORT_14_addr = 6'h3;
  assign LUT_mem_MPORT_14_mask = 1'h1;
  assign LUT_mem_MPORT_14_en = io_dispatch_3 ? 1'h0 : 1'h1;
  assign LUT_mem_MPORT_16_data = {1'h0,lo_4};
  assign LUT_mem_MPORT_16_addr = 6'h4;
  assign LUT_mem_MPORT_16_mask = 1'h1;
  assign LUT_mem_MPORT_16_en = io_dispatch_4;
  assign LUT_mem_MPORT_18_data = LUT_mem_MPORT_19_data;
  assign LUT_mem_MPORT_18_addr = 6'h4;
  assign LUT_mem_MPORT_18_mask = 1'h1;
  assign LUT_mem_MPORT_18_en = io_dispatch_4 ? 1'h0 : 1'h1;
  assign LUT_mem_MPORT_20_data = {1'h0,lo_5};
  assign LUT_mem_MPORT_20_addr = 6'h5;
  assign LUT_mem_MPORT_20_mask = 1'h1;
  assign LUT_mem_MPORT_20_en = io_dispatch_5;
  assign LUT_mem_MPORT_22_data = LUT_mem_MPORT_23_data;
  assign LUT_mem_MPORT_22_addr = 6'h5;
  assign LUT_mem_MPORT_22_mask = 1'h1;
  assign LUT_mem_MPORT_22_en = io_dispatch_5 ? 1'h0 : 1'h1;
  assign LUT_mem_MPORT_24_data = {1'h0,lo_6};
  assign LUT_mem_MPORT_24_addr = 6'h6;
  assign LUT_mem_MPORT_24_mask = 1'h1;
  assign LUT_mem_MPORT_24_en = io_dispatch_6;
  assign LUT_mem_MPORT_26_data = LUT_mem_MPORT_27_data;
  assign LUT_mem_MPORT_26_addr = 6'h6;
  assign LUT_mem_MPORT_26_mask = 1'h1;
  assign LUT_mem_MPORT_26_en = io_dispatch_6 ? 1'h0 : 1'h1;
  assign LUT_mem_MPORT_28_data = {1'h0,lo_7};
  assign LUT_mem_MPORT_28_addr = 6'h7;
  assign LUT_mem_MPORT_28_mask = 1'h1;
  assign LUT_mem_MPORT_28_en = io_dispatch_7;
  assign LUT_mem_MPORT_30_data = LUT_mem_MPORT_31_data;
  assign LUT_mem_MPORT_30_addr = 6'h7;
  assign LUT_mem_MPORT_30_mask = 1'h1;
  assign LUT_mem_MPORT_30_en = io_dispatch_7 ? 1'h0 : 1'h1;
  assign LUT_mem_MPORT_32_data = {1'h0,lo_8};
  assign LUT_mem_MPORT_32_addr = 6'h8;
  assign LUT_mem_MPORT_32_mask = 1'h1;
  assign LUT_mem_MPORT_32_en = io_dispatch_8;
  assign LUT_mem_MPORT_34_data = LUT_mem_MPORT_35_data;
  assign LUT_mem_MPORT_34_addr = 6'h8;
  assign LUT_mem_MPORT_34_mask = 1'h1;
  assign LUT_mem_MPORT_34_en = io_dispatch_8 ? 1'h0 : 1'h1;
  assign LUT_mem_MPORT_36_data = {1'h0,lo_9};
  assign LUT_mem_MPORT_36_addr = 6'h9;
  assign LUT_mem_MPORT_36_mask = 1'h1;
  assign LUT_mem_MPORT_36_en = io_dispatch_9;
  assign LUT_mem_MPORT_38_data = LUT_mem_MPORT_39_data;
  assign LUT_mem_MPORT_38_addr = 6'h9;
  assign LUT_mem_MPORT_38_mask = 1'h1;
  assign LUT_mem_MPORT_38_en = io_dispatch_9 ? 1'h0 : 1'h1;
  assign LUT_mem_MPORT_40_data = {1'h0,lo_10};
  assign LUT_mem_MPORT_40_addr = 6'ha;
  assign LUT_mem_MPORT_40_mask = 1'h1;
  assign LUT_mem_MPORT_40_en = io_dispatch_10;
  assign LUT_mem_MPORT_42_data = LUT_mem_MPORT_43_data;
  assign LUT_mem_MPORT_42_addr = 6'ha;
  assign LUT_mem_MPORT_42_mask = 1'h1;
  assign LUT_mem_MPORT_42_en = io_dispatch_10 ? 1'h0 : 1'h1;
  assign LUT_mem_MPORT_44_data = {1'h0,lo_11};
  assign LUT_mem_MPORT_44_addr = 6'hb;
  assign LUT_mem_MPORT_44_mask = 1'h1;
  assign LUT_mem_MPORT_44_en = io_dispatch_11;
  assign LUT_mem_MPORT_46_data = LUT_mem_MPORT_47_data;
  assign LUT_mem_MPORT_46_addr = 6'hb;
  assign LUT_mem_MPORT_46_mask = 1'h1;
  assign LUT_mem_MPORT_46_en = io_dispatch_11 ? 1'h0 : 1'h1;
  assign LUT_mem_MPORT_48_data = {1'h0,lo_12};
  assign LUT_mem_MPORT_48_addr = 6'hc;
  assign LUT_mem_MPORT_48_mask = 1'h1;
  assign LUT_mem_MPORT_48_en = io_dispatch_12;
  assign LUT_mem_MPORT_50_data = LUT_mem_MPORT_51_data;
  assign LUT_mem_MPORT_50_addr = 6'hc;
  assign LUT_mem_MPORT_50_mask = 1'h1;
  assign LUT_mem_MPORT_50_en = io_dispatch_12 ? 1'h0 : 1'h1;
  assign LUT_mem_MPORT_52_data = {1'h0,lo_13};
  assign LUT_mem_MPORT_52_addr = 6'hd;
  assign LUT_mem_MPORT_52_mask = 1'h1;
  assign LUT_mem_MPORT_52_en = io_dispatch_13;
  assign LUT_mem_MPORT_54_data = LUT_mem_MPORT_55_data;
  assign LUT_mem_MPORT_54_addr = 6'hd;
  assign LUT_mem_MPORT_54_mask = 1'h1;
  assign LUT_mem_MPORT_54_en = io_dispatch_13 ? 1'h0 : 1'h1;
  assign LUT_mem_MPORT_56_data = {1'h0,lo_14};
  assign LUT_mem_MPORT_56_addr = 6'he;
  assign LUT_mem_MPORT_56_mask = 1'h1;
  assign LUT_mem_MPORT_56_en = io_dispatch_14;
  assign LUT_mem_MPORT_58_data = LUT_mem_MPORT_59_data;
  assign LUT_mem_MPORT_58_addr = 6'he;
  assign LUT_mem_MPORT_58_mask = 1'h1;
  assign LUT_mem_MPORT_58_en = io_dispatch_14 ? 1'h0 : 1'h1;
  assign LUT_mem_MPORT_60_data = {1'h0,lo_15};
  assign LUT_mem_MPORT_60_addr = 6'hf;
  assign LUT_mem_MPORT_60_mask = 1'h1;
  assign LUT_mem_MPORT_60_en = io_dispatch_15;
  assign LUT_mem_MPORT_62_data = LUT_mem_MPORT_63_data;
  assign LUT_mem_MPORT_62_addr = 6'hf;
  assign LUT_mem_MPORT_62_mask = 1'h1;
  assign LUT_mem_MPORT_62_en = io_dispatch_15 ? 1'h0 : 1'h1;
  assign LUT_mem_MPORT_64_data = {1'h0,lo_16};
  assign LUT_mem_MPORT_64_addr = 6'h10;
  assign LUT_mem_MPORT_64_mask = 1'h1;
  assign LUT_mem_MPORT_64_en = io_dispatch_16;
  assign LUT_mem_MPORT_66_data = LUT_mem_MPORT_67_data;
  assign LUT_mem_MPORT_66_addr = 6'h10;
  assign LUT_mem_MPORT_66_mask = 1'h1;
  assign LUT_mem_MPORT_66_en = io_dispatch_16 ? 1'h0 : 1'h1;
  assign LUT_mem_MPORT_68_data = {1'h0,lo_17};
  assign LUT_mem_MPORT_68_addr = 6'h11;
  assign LUT_mem_MPORT_68_mask = 1'h1;
  assign LUT_mem_MPORT_68_en = io_dispatch_17;
  assign LUT_mem_MPORT_70_data = LUT_mem_MPORT_71_data;
  assign LUT_mem_MPORT_70_addr = 6'h11;
  assign LUT_mem_MPORT_70_mask = 1'h1;
  assign LUT_mem_MPORT_70_en = io_dispatch_17 ? 1'h0 : 1'h1;
  assign LUT_mem_MPORT_72_data = {1'h0,lo_18};
  assign LUT_mem_MPORT_72_addr = 6'h12;
  assign LUT_mem_MPORT_72_mask = 1'h1;
  assign LUT_mem_MPORT_72_en = io_dispatch_18;
  assign LUT_mem_MPORT_74_data = LUT_mem_MPORT_75_data;
  assign LUT_mem_MPORT_74_addr = 6'h12;
  assign LUT_mem_MPORT_74_mask = 1'h1;
  assign LUT_mem_MPORT_74_en = io_dispatch_18 ? 1'h0 : 1'h1;
  assign LUT_mem_MPORT_76_data = {1'h0,lo_19};
  assign LUT_mem_MPORT_76_addr = 6'h13;
  assign LUT_mem_MPORT_76_mask = 1'h1;
  assign LUT_mem_MPORT_76_en = io_dispatch_19;
  assign LUT_mem_MPORT_78_data = LUT_mem_MPORT_79_data;
  assign LUT_mem_MPORT_78_addr = 6'h13;
  assign LUT_mem_MPORT_78_mask = 1'h1;
  assign LUT_mem_MPORT_78_en = io_dispatch_19 ? 1'h0 : 1'h1;
  assign LUT_mem_MPORT_80_data = {1'h0,lo_20};
  assign LUT_mem_MPORT_80_addr = 6'h14;
  assign LUT_mem_MPORT_80_mask = 1'h1;
  assign LUT_mem_MPORT_80_en = io_dispatch_20;
  assign LUT_mem_MPORT_82_data = LUT_mem_MPORT_83_data;
  assign LUT_mem_MPORT_82_addr = 6'h14;
  assign LUT_mem_MPORT_82_mask = 1'h1;
  assign LUT_mem_MPORT_82_en = io_dispatch_20 ? 1'h0 : 1'h1;
  assign LUT_mem_MPORT_84_data = {1'h0,lo_21};
  assign LUT_mem_MPORT_84_addr = 6'h15;
  assign LUT_mem_MPORT_84_mask = 1'h1;
  assign LUT_mem_MPORT_84_en = io_dispatch_21;
  assign LUT_mem_MPORT_86_data = LUT_mem_MPORT_87_data;
  assign LUT_mem_MPORT_86_addr = 6'h15;
  assign LUT_mem_MPORT_86_mask = 1'h1;
  assign LUT_mem_MPORT_86_en = io_dispatch_21 ? 1'h0 : 1'h1;
  assign LUT_mem_MPORT_88_data = {1'h0,lo_22};
  assign LUT_mem_MPORT_88_addr = 6'h16;
  assign LUT_mem_MPORT_88_mask = 1'h1;
  assign LUT_mem_MPORT_88_en = io_dispatch_22;
  assign LUT_mem_MPORT_90_data = LUT_mem_MPORT_91_data;
  assign LUT_mem_MPORT_90_addr = 6'h16;
  assign LUT_mem_MPORT_90_mask = 1'h1;
  assign LUT_mem_MPORT_90_en = io_dispatch_22 ? 1'h0 : 1'h1;
  assign LUT_mem_MPORT_92_data = {1'h0,lo_23};
  assign LUT_mem_MPORT_92_addr = 6'h17;
  assign LUT_mem_MPORT_92_mask = 1'h1;
  assign LUT_mem_MPORT_92_en = io_dispatch_23;
  assign LUT_mem_MPORT_94_data = LUT_mem_MPORT_95_data;
  assign LUT_mem_MPORT_94_addr = 6'h17;
  assign LUT_mem_MPORT_94_mask = 1'h1;
  assign LUT_mem_MPORT_94_en = io_dispatch_23 ? 1'h0 : 1'h1;
  assign LUT_mem_MPORT_96_data = {1'h0,lo_24};
  assign LUT_mem_MPORT_96_addr = 6'h18;
  assign LUT_mem_MPORT_96_mask = 1'h1;
  assign LUT_mem_MPORT_96_en = io_dispatch_24;
  assign LUT_mem_MPORT_98_data = LUT_mem_MPORT_99_data;
  assign LUT_mem_MPORT_98_addr = 6'h18;
  assign LUT_mem_MPORT_98_mask = 1'h1;
  assign LUT_mem_MPORT_98_en = io_dispatch_24 ? 1'h0 : 1'h1;
  assign LUT_mem_MPORT_100_data = {1'h0,lo_25};
  assign LUT_mem_MPORT_100_addr = 6'h19;
  assign LUT_mem_MPORT_100_mask = 1'h1;
  assign LUT_mem_MPORT_100_en = io_dispatch_25;
  assign LUT_mem_MPORT_102_data = LUT_mem_MPORT_103_data;
  assign LUT_mem_MPORT_102_addr = 6'h19;
  assign LUT_mem_MPORT_102_mask = 1'h1;
  assign LUT_mem_MPORT_102_en = io_dispatch_25 ? 1'h0 : 1'h1;
  assign LUT_mem_MPORT_104_data = {1'h0,lo_26};
  assign LUT_mem_MPORT_104_addr = 6'h1a;
  assign LUT_mem_MPORT_104_mask = 1'h1;
  assign LUT_mem_MPORT_104_en = io_dispatch_26;
  assign LUT_mem_MPORT_106_data = LUT_mem_MPORT_107_data;
  assign LUT_mem_MPORT_106_addr = 6'h1a;
  assign LUT_mem_MPORT_106_mask = 1'h1;
  assign LUT_mem_MPORT_106_en = io_dispatch_26 ? 1'h0 : 1'h1;
  assign LUT_mem_MPORT_108_data = {1'h0,lo_27};
  assign LUT_mem_MPORT_108_addr = 6'h1b;
  assign LUT_mem_MPORT_108_mask = 1'h1;
  assign LUT_mem_MPORT_108_en = io_dispatch_27;
  assign LUT_mem_MPORT_110_data = LUT_mem_MPORT_111_data;
  assign LUT_mem_MPORT_110_addr = 6'h1b;
  assign LUT_mem_MPORT_110_mask = 1'h1;
  assign LUT_mem_MPORT_110_en = io_dispatch_27 ? 1'h0 : 1'h1;
  assign LUT_mem_MPORT_112_data = {1'h0,lo_28};
  assign LUT_mem_MPORT_112_addr = 6'h1c;
  assign LUT_mem_MPORT_112_mask = 1'h1;
  assign LUT_mem_MPORT_112_en = io_dispatch_28;
  assign LUT_mem_MPORT_114_data = LUT_mem_MPORT_115_data;
  assign LUT_mem_MPORT_114_addr = 6'h1c;
  assign LUT_mem_MPORT_114_mask = 1'h1;
  assign LUT_mem_MPORT_114_en = io_dispatch_28 ? 1'h0 : 1'h1;
  assign LUT_mem_MPORT_116_data = {1'h0,lo_29};
  assign LUT_mem_MPORT_116_addr = 6'h1d;
  assign LUT_mem_MPORT_116_mask = 1'h1;
  assign LUT_mem_MPORT_116_en = io_dispatch_29;
  assign LUT_mem_MPORT_118_data = LUT_mem_MPORT_119_data;
  assign LUT_mem_MPORT_118_addr = 6'h1d;
  assign LUT_mem_MPORT_118_mask = 1'h1;
  assign LUT_mem_MPORT_118_en = io_dispatch_29 ? 1'h0 : 1'h1;
  assign LUT_mem_MPORT_120_data = {1'h0,lo_30};
  assign LUT_mem_MPORT_120_addr = 6'h1e;
  assign LUT_mem_MPORT_120_mask = 1'h1;
  assign LUT_mem_MPORT_120_en = io_dispatch_30;
  assign LUT_mem_MPORT_122_data = LUT_mem_MPORT_123_data;
  assign LUT_mem_MPORT_122_addr = 6'h1e;
  assign LUT_mem_MPORT_122_mask = 1'h1;
  assign LUT_mem_MPORT_122_en = io_dispatch_30 ? 1'h0 : 1'h1;
  assign LUT_mem_MPORT_124_data = {1'h0,lo_31};
  assign LUT_mem_MPORT_124_addr = 6'h1f;
  assign LUT_mem_MPORT_124_mask = 1'h1;
  assign LUT_mem_MPORT_124_en = io_dispatch_31;
  assign LUT_mem_MPORT_126_data = LUT_mem_MPORT_127_data;
  assign LUT_mem_MPORT_126_addr = 6'h1f;
  assign LUT_mem_MPORT_126_mask = 1'h1;
  assign LUT_mem_MPORT_126_en = io_dispatch_31 ? 1'h0 : 1'h1;
  assign LUT_mem_MPORT_128_data = {1'h0,lo_32};
  assign LUT_mem_MPORT_128_addr = 6'h20;
  assign LUT_mem_MPORT_128_mask = 1'h1;
  assign LUT_mem_MPORT_128_en = io_dispatch_32;
  assign LUT_mem_MPORT_130_data = LUT_mem_MPORT_131_data;
  assign LUT_mem_MPORT_130_addr = 6'h20;
  assign LUT_mem_MPORT_130_mask = 1'h1;
  assign LUT_mem_MPORT_130_en = io_dispatch_32 ? 1'h0 : 1'h1;
  assign LUT_mem_MPORT_132_data = {1'h0,lo_33};
  assign LUT_mem_MPORT_132_addr = 6'h21;
  assign LUT_mem_MPORT_132_mask = 1'h1;
  assign LUT_mem_MPORT_132_en = io_dispatch_33;
  assign LUT_mem_MPORT_134_data = LUT_mem_MPORT_135_data;
  assign LUT_mem_MPORT_134_addr = 6'h21;
  assign LUT_mem_MPORT_134_mask = 1'h1;
  assign LUT_mem_MPORT_134_en = io_dispatch_33 ? 1'h0 : 1'h1;
  assign LUT_mem_MPORT_136_data = {1'h0,lo_34};
  assign LUT_mem_MPORT_136_addr = 6'h22;
  assign LUT_mem_MPORT_136_mask = 1'h1;
  assign LUT_mem_MPORT_136_en = io_dispatch_34;
  assign LUT_mem_MPORT_138_data = LUT_mem_MPORT_139_data;
  assign LUT_mem_MPORT_138_addr = 6'h22;
  assign LUT_mem_MPORT_138_mask = 1'h1;
  assign LUT_mem_MPORT_138_en = io_dispatch_34 ? 1'h0 : 1'h1;
  assign LUT_mem_MPORT_211_data = {1'h1,push_ray_id};
  assign LUT_mem_MPORT_211_addr = 6'h0;
  assign LUT_mem_MPORT_211_mask = 1'h1;
  assign LUT_mem_MPORT_211_en = _T_109 & _GEN_18869;
  assign LUT_mem_MPORT_213_data = {1'h1,push_ray_id};
  assign LUT_mem_MPORT_213_addr = 6'h1;
  assign LUT_mem_MPORT_213_mask = 1'h1;
  assign LUT_mem_MPORT_213_en = _T_109 & _GEN_18877;
  assign LUT_mem_MPORT_215_data = {1'h1,push_ray_id};
  assign LUT_mem_MPORT_215_addr = 6'h2;
  assign LUT_mem_MPORT_215_mask = 1'h1;
  assign LUT_mem_MPORT_215_en = _T_109 & _GEN_18884;
  assign LUT_mem_MPORT_217_data = {1'h1,push_ray_id};
  assign LUT_mem_MPORT_217_addr = 6'h3;
  assign LUT_mem_MPORT_217_mask = 1'h1;
  assign LUT_mem_MPORT_217_en = _T_109 & _GEN_18892;
  assign LUT_mem_MPORT_219_data = {1'h1,push_ray_id};
  assign LUT_mem_MPORT_219_addr = 6'h4;
  assign LUT_mem_MPORT_219_mask = 1'h1;
  assign LUT_mem_MPORT_219_en = _T_109 & _GEN_18900;
  assign LUT_mem_MPORT_221_data = {1'h1,push_ray_id};
  assign LUT_mem_MPORT_221_addr = 6'h5;
  assign LUT_mem_MPORT_221_mask = 1'h1;
  assign LUT_mem_MPORT_221_en = _T_109 & _GEN_18908;
  assign LUT_mem_MPORT_223_data = {1'h1,push_ray_id};
  assign LUT_mem_MPORT_223_addr = 6'h6;
  assign LUT_mem_MPORT_223_mask = 1'h1;
  assign LUT_mem_MPORT_223_en = _T_109 & _GEN_18916;
  assign LUT_mem_MPORT_225_data = {1'h1,push_ray_id};
  assign LUT_mem_MPORT_225_addr = 6'h7;
  assign LUT_mem_MPORT_225_mask = 1'h1;
  assign LUT_mem_MPORT_225_en = _T_109 & _GEN_18924;
  assign LUT_mem_MPORT_227_data = {1'h1,push_ray_id};
  assign LUT_mem_MPORT_227_addr = 6'h8;
  assign LUT_mem_MPORT_227_mask = 1'h1;
  assign LUT_mem_MPORT_227_en = _T_109 & _GEN_18932;
  assign LUT_mem_MPORT_229_data = {1'h1,push_ray_id};
  assign LUT_mem_MPORT_229_addr = 6'h9;
  assign LUT_mem_MPORT_229_mask = 1'h1;
  assign LUT_mem_MPORT_229_en = _T_109 & _GEN_18940;
  assign LUT_mem_MPORT_231_data = {1'h1,push_ray_id};
  assign LUT_mem_MPORT_231_addr = 6'ha;
  assign LUT_mem_MPORT_231_mask = 1'h1;
  assign LUT_mem_MPORT_231_en = _T_109 & _GEN_18948;
  assign LUT_mem_MPORT_233_data = {1'h1,push_ray_id};
  assign LUT_mem_MPORT_233_addr = 6'hb;
  assign LUT_mem_MPORT_233_mask = 1'h1;
  assign LUT_mem_MPORT_233_en = _T_109 & _GEN_18956;
  assign LUT_mem_MPORT_235_data = {1'h1,push_ray_id};
  assign LUT_mem_MPORT_235_addr = 6'hc;
  assign LUT_mem_MPORT_235_mask = 1'h1;
  assign LUT_mem_MPORT_235_en = _T_109 & _GEN_18964;
  assign LUT_mem_MPORT_237_data = {1'h1,push_ray_id};
  assign LUT_mem_MPORT_237_addr = 6'hd;
  assign LUT_mem_MPORT_237_mask = 1'h1;
  assign LUT_mem_MPORT_237_en = _T_109 & _GEN_18972;
  assign LUT_mem_MPORT_239_data = {1'h1,push_ray_id};
  assign LUT_mem_MPORT_239_addr = 6'he;
  assign LUT_mem_MPORT_239_mask = 1'h1;
  assign LUT_mem_MPORT_239_en = _T_109 & _GEN_18980;
  assign LUT_mem_MPORT_241_data = {1'h1,push_ray_id};
  assign LUT_mem_MPORT_241_addr = 6'hf;
  assign LUT_mem_MPORT_241_mask = 1'h1;
  assign LUT_mem_MPORT_241_en = _T_109 & _GEN_18988;
  assign LUT_mem_MPORT_243_data = {1'h1,push_ray_id};
  assign LUT_mem_MPORT_243_addr = 6'h10;
  assign LUT_mem_MPORT_243_mask = 1'h1;
  assign LUT_mem_MPORT_243_en = _T_109 & _GEN_18996;
  assign LUT_mem_MPORT_245_data = {1'h1,push_ray_id};
  assign LUT_mem_MPORT_245_addr = 6'h11;
  assign LUT_mem_MPORT_245_mask = 1'h1;
  assign LUT_mem_MPORT_245_en = _T_109 & _GEN_19004;
  assign LUT_mem_MPORT_247_data = {1'h1,push_ray_id};
  assign LUT_mem_MPORT_247_addr = 6'h12;
  assign LUT_mem_MPORT_247_mask = 1'h1;
  assign LUT_mem_MPORT_247_en = _T_109 & _GEN_19012;
  assign LUT_mem_MPORT_249_data = {1'h1,push_ray_id};
  assign LUT_mem_MPORT_249_addr = 6'h13;
  assign LUT_mem_MPORT_249_mask = 1'h1;
  assign LUT_mem_MPORT_249_en = _T_109 & _GEN_19020;
  assign LUT_mem_MPORT_251_data = {1'h1,push_ray_id};
  assign LUT_mem_MPORT_251_addr = 6'h14;
  assign LUT_mem_MPORT_251_mask = 1'h1;
  assign LUT_mem_MPORT_251_en = _T_109 & _GEN_19028;
  assign LUT_mem_MPORT_253_data = {1'h1,push_ray_id};
  assign LUT_mem_MPORT_253_addr = 6'h15;
  assign LUT_mem_MPORT_253_mask = 1'h1;
  assign LUT_mem_MPORT_253_en = _T_109 & _GEN_19036;
  assign LUT_mem_MPORT_255_data = {1'h1,push_ray_id};
  assign LUT_mem_MPORT_255_addr = 6'h16;
  assign LUT_mem_MPORT_255_mask = 1'h1;
  assign LUT_mem_MPORT_255_en = _T_109 & _GEN_19044;
  assign LUT_mem_MPORT_257_data = {1'h1,push_ray_id};
  assign LUT_mem_MPORT_257_addr = 6'h17;
  assign LUT_mem_MPORT_257_mask = 1'h1;
  assign LUT_mem_MPORT_257_en = _T_109 & _GEN_19052;
  assign LUT_mem_MPORT_259_data = {1'h1,push_ray_id};
  assign LUT_mem_MPORT_259_addr = 6'h18;
  assign LUT_mem_MPORT_259_mask = 1'h1;
  assign LUT_mem_MPORT_259_en = _T_109 & _GEN_19060;
  assign LUT_mem_MPORT_261_data = {1'h1,push_ray_id};
  assign LUT_mem_MPORT_261_addr = 6'h19;
  assign LUT_mem_MPORT_261_mask = 1'h1;
  assign LUT_mem_MPORT_261_en = _T_109 & _GEN_19068;
  assign LUT_mem_MPORT_263_data = {1'h1,push_ray_id};
  assign LUT_mem_MPORT_263_addr = 6'h1a;
  assign LUT_mem_MPORT_263_mask = 1'h1;
  assign LUT_mem_MPORT_263_en = _T_109 & _GEN_19076;
  assign LUT_mem_MPORT_265_data = {1'h1,push_ray_id};
  assign LUT_mem_MPORT_265_addr = 6'h1b;
  assign LUT_mem_MPORT_265_mask = 1'h1;
  assign LUT_mem_MPORT_265_en = _T_109 & _GEN_19084;
  assign LUT_mem_MPORT_267_data = {1'h1,push_ray_id};
  assign LUT_mem_MPORT_267_addr = 6'h1c;
  assign LUT_mem_MPORT_267_mask = 1'h1;
  assign LUT_mem_MPORT_267_en = _T_109 & _GEN_19092;
  assign LUT_mem_MPORT_269_data = {1'h1,push_ray_id};
  assign LUT_mem_MPORT_269_addr = 6'h1d;
  assign LUT_mem_MPORT_269_mask = 1'h1;
  assign LUT_mem_MPORT_269_en = _T_109 & _GEN_19100;
  assign LUT_mem_MPORT_271_data = {1'h1,push_ray_id};
  assign LUT_mem_MPORT_271_addr = 6'h1e;
  assign LUT_mem_MPORT_271_mask = 1'h1;
  assign LUT_mem_MPORT_271_en = _T_109 & _GEN_19108;
  assign LUT_mem_MPORT_273_data = {1'h1,push_ray_id};
  assign LUT_mem_MPORT_273_addr = 6'h1f;
  assign LUT_mem_MPORT_273_mask = 1'h1;
  assign LUT_mem_MPORT_273_en = _T_109 & _GEN_19116;
  assign LUT_mem_MPORT_275_data = {1'h1,push_ray_id};
  assign LUT_mem_MPORT_275_addr = 6'h20;
  assign LUT_mem_MPORT_275_mask = 1'h1;
  assign LUT_mem_MPORT_275_en = _T_109 & _GEN_19124;
  assign LUT_mem_MPORT_277_data = {1'h1,push_ray_id};
  assign LUT_mem_MPORT_277_addr = 6'h21;
  assign LUT_mem_MPORT_277_mask = 1'h1;
  assign LUT_mem_MPORT_277_en = _T_109 & _GEN_19132;
  assign LUT_mem_MPORT_279_data = {1'h1,push_ray_id};
  assign LUT_mem_MPORT_279_addr = 6'h22;
  assign LUT_mem_MPORT_279_mask = 1'h1;
  assign LUT_mem_MPORT_279_en = _T_109 & _GEN_19140;
  assign io_ray_id_pop_out = pop_ray_id_2; // @[lut_35.scala 5208:46]
  assign io_hitT_out = pop_hitT_2; // @[lut_35.scala 5209:56]
  assign io_pop_0 = pop_0_1; // @[lut_35.scala 5166:57]
  assign io_pop_1 = pop_1_1; // @[lut_35.scala 5167:57]
  assign io_pop_2 = pop_2_1; // @[lut_35.scala 5168:57]
  assign io_pop_3 = pop_3_1; // @[lut_35.scala 5169:57]
  assign io_pop_4 = pop_4_1; // @[lut_35.scala 5170:57]
  assign io_pop_5 = pop_5_1; // @[lut_35.scala 5171:57]
  assign io_pop_6 = pop_6_1; // @[lut_35.scala 5172:57]
  assign io_pop_7 = pop_7_1; // @[lut_35.scala 5173:57]
  assign io_pop_8 = pop_8_1; // @[lut_35.scala 5174:57]
  assign io_pop_9 = pop_9_1; // @[lut_35.scala 5175:57]
  assign io_pop_10 = pop_10_1; // @[lut_35.scala 5177:58]
  assign io_pop_11 = pop_11_1; // @[lut_35.scala 5178:58]
  assign io_pop_12 = pop_12_1; // @[lut_35.scala 5179:58]
  assign io_pop_13 = pop_13_1; // @[lut_35.scala 5180:58]
  assign io_pop_14 = pop_14_1; // @[lut_35.scala 5181:58]
  assign io_pop_15 = pop_15_1; // @[lut_35.scala 5182:58]
  assign io_pop_16 = pop_16_1; // @[lut_35.scala 5183:58]
  assign io_pop_17 = pop_17_1; // @[lut_35.scala 5184:58]
  assign io_pop_18 = pop_18_1; // @[lut_35.scala 5185:58]
  assign io_pop_19 = pop_19_1; // @[lut_35.scala 5186:58]
  assign io_pop_20 = pop_20_1; // @[lut_35.scala 5188:58]
  assign io_pop_21 = pop_21_1; // @[lut_35.scala 5189:58]
  assign io_pop_22 = pop_22_1; // @[lut_35.scala 5190:58]
  assign io_pop_23 = pop_23_1; // @[lut_35.scala 5191:58]
  assign io_pop_24 = pop_24_1; // @[lut_35.scala 5192:58]
  assign io_pop_25 = pop_25_1; // @[lut_35.scala 5193:58]
  assign io_pop_26 = pop_26_1; // @[lut_35.scala 5194:58]
  assign io_pop_27 = pop_27_1; // @[lut_35.scala 5195:58]
  assign io_pop_28 = pop_28_1; // @[lut_35.scala 5196:58]
  assign io_pop_29 = pop_29_1; // @[lut_35.scala 5197:58]
  assign io_pop_30 = pop_30_1; // @[lut_35.scala 5199:58]
  assign io_pop_31 = pop_31_1; // @[lut_35.scala 5200:58]
  assign io_pop_32 = pop_32_1; // @[lut_35.scala 5201:58]
  assign io_pop_33 = pop_33_1; // @[lut_35.scala 5202:58]
  assign io_pop_34 = pop_34_1; // @[lut_35.scala 5203:58]
  assign io_pop_en = pop_valid_2; // @[lut_35.scala 5207:55]
  assign io_push_0 = push_0_1; // @[lut_35.scala 3493:51]
  assign io_push_1 = push_1_1; // @[lut_35.scala 3494:51]
  assign io_push_2 = push_2_1; // @[lut_35.scala 3495:51]
  assign io_push_3 = push_3_1; // @[lut_35.scala 3496:51]
  assign io_push_4 = push_4_1; // @[lut_35.scala 3497:51]
  assign io_push_5 = push_5_1; // @[lut_35.scala 3498:51]
  assign io_push_6 = push_6_1; // @[lut_35.scala 3499:51]
  assign io_push_7 = push_7_1; // @[lut_35.scala 3500:51]
  assign io_push_8 = push_8_1; // @[lut_35.scala 3501:51]
  assign io_push_9 = push_9_1; // @[lut_35.scala 3502:51]
  assign io_push_10 = push_10_1; // @[lut_35.scala 3503:52]
  assign io_push_11 = push_11_1; // @[lut_35.scala 3504:52]
  assign io_push_12 = push_12_1; // @[lut_35.scala 3505:52]
  assign io_push_13 = push_13_1; // @[lut_35.scala 3506:52]
  assign io_push_14 = push_14_1; // @[lut_35.scala 3507:52]
  assign io_push_15 = push_15_1; // @[lut_35.scala 3508:52]
  assign io_push_16 = push_16_1; // @[lut_35.scala 3509:52]
  assign io_push_17 = push_17_1; // @[lut_35.scala 3510:52]
  assign io_push_18 = push_18_1; // @[lut_35.scala 3511:52]
  assign io_push_19 = push_19_1; // @[lut_35.scala 3512:52]
  assign io_push_20 = push_20_1; // @[lut_35.scala 3513:52]
  assign io_push_21 = push_21_1; // @[lut_35.scala 3514:52]
  assign io_push_22 = push_22_1; // @[lut_35.scala 3515:52]
  assign io_push_23 = push_23_1; // @[lut_35.scala 3516:52]
  assign io_push_24 = push_24_1; // @[lut_35.scala 3517:52]
  assign io_push_25 = push_25_1; // @[lut_35.scala 3518:52]
  assign io_push_26 = push_26_1; // @[lut_35.scala 3519:52]
  assign io_push_27 = push_27_1; // @[lut_35.scala 3520:52]
  assign io_push_28 = push_28_1; // @[lut_35.scala 3521:52]
  assign io_push_29 = push_29_1; // @[lut_35.scala 3522:52]
  assign io_push_30 = push_30_1; // @[lut_35.scala 3523:52]
  assign io_push_31 = push_31_1; // @[lut_35.scala 3524:52]
  assign io_push_32 = push_32_1; // @[lut_35.scala 3525:52]
  assign io_push_33 = push_33_1; // @[lut_35.scala 3526:52]
  assign io_push_34 = push_34_1; // @[lut_35.scala 3527:52]
  assign io_push_en = push_valid_2; // @[lut_35.scala 3530:50]
  assign io_no_match = no_match_2; // @[lut_35.scala 3686:41]
  always @(posedge clock) begin
    if(LUT_mem_MPORT_en & LUT_mem_MPORT_mask) begin
      LUT_mem[LUT_mem_MPORT_addr] <= LUT_mem_MPORT_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_2_en & LUT_mem_MPORT_2_mask) begin
      LUT_mem[LUT_mem_MPORT_2_addr] <= LUT_mem_MPORT_2_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_4_en & LUT_mem_MPORT_4_mask) begin
      LUT_mem[LUT_mem_MPORT_4_addr] <= LUT_mem_MPORT_4_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_6_en & LUT_mem_MPORT_6_mask) begin
      LUT_mem[LUT_mem_MPORT_6_addr] <= LUT_mem_MPORT_6_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_8_en & LUT_mem_MPORT_8_mask) begin
      LUT_mem[LUT_mem_MPORT_8_addr] <= LUT_mem_MPORT_8_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_10_en & LUT_mem_MPORT_10_mask) begin
      LUT_mem[LUT_mem_MPORT_10_addr] <= LUT_mem_MPORT_10_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_12_en & LUT_mem_MPORT_12_mask) begin
      LUT_mem[LUT_mem_MPORT_12_addr] <= LUT_mem_MPORT_12_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_14_en & LUT_mem_MPORT_14_mask) begin
      LUT_mem[LUT_mem_MPORT_14_addr] <= LUT_mem_MPORT_14_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_16_en & LUT_mem_MPORT_16_mask) begin
      LUT_mem[LUT_mem_MPORT_16_addr] <= LUT_mem_MPORT_16_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_18_en & LUT_mem_MPORT_18_mask) begin
      LUT_mem[LUT_mem_MPORT_18_addr] <= LUT_mem_MPORT_18_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_20_en & LUT_mem_MPORT_20_mask) begin
      LUT_mem[LUT_mem_MPORT_20_addr] <= LUT_mem_MPORT_20_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_22_en & LUT_mem_MPORT_22_mask) begin
      LUT_mem[LUT_mem_MPORT_22_addr] <= LUT_mem_MPORT_22_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_24_en & LUT_mem_MPORT_24_mask) begin
      LUT_mem[LUT_mem_MPORT_24_addr] <= LUT_mem_MPORT_24_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_26_en & LUT_mem_MPORT_26_mask) begin
      LUT_mem[LUT_mem_MPORT_26_addr] <= LUT_mem_MPORT_26_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_28_en & LUT_mem_MPORT_28_mask) begin
      LUT_mem[LUT_mem_MPORT_28_addr] <= LUT_mem_MPORT_28_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_30_en & LUT_mem_MPORT_30_mask) begin
      LUT_mem[LUT_mem_MPORT_30_addr] <= LUT_mem_MPORT_30_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_32_en & LUT_mem_MPORT_32_mask) begin
      LUT_mem[LUT_mem_MPORT_32_addr] <= LUT_mem_MPORT_32_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_34_en & LUT_mem_MPORT_34_mask) begin
      LUT_mem[LUT_mem_MPORT_34_addr] <= LUT_mem_MPORT_34_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_36_en & LUT_mem_MPORT_36_mask) begin
      LUT_mem[LUT_mem_MPORT_36_addr] <= LUT_mem_MPORT_36_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_38_en & LUT_mem_MPORT_38_mask) begin
      LUT_mem[LUT_mem_MPORT_38_addr] <= LUT_mem_MPORT_38_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_40_en & LUT_mem_MPORT_40_mask) begin
      LUT_mem[LUT_mem_MPORT_40_addr] <= LUT_mem_MPORT_40_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_42_en & LUT_mem_MPORT_42_mask) begin
      LUT_mem[LUT_mem_MPORT_42_addr] <= LUT_mem_MPORT_42_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_44_en & LUT_mem_MPORT_44_mask) begin
      LUT_mem[LUT_mem_MPORT_44_addr] <= LUT_mem_MPORT_44_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_46_en & LUT_mem_MPORT_46_mask) begin
      LUT_mem[LUT_mem_MPORT_46_addr] <= LUT_mem_MPORT_46_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_48_en & LUT_mem_MPORT_48_mask) begin
      LUT_mem[LUT_mem_MPORT_48_addr] <= LUT_mem_MPORT_48_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_50_en & LUT_mem_MPORT_50_mask) begin
      LUT_mem[LUT_mem_MPORT_50_addr] <= LUT_mem_MPORT_50_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_52_en & LUT_mem_MPORT_52_mask) begin
      LUT_mem[LUT_mem_MPORT_52_addr] <= LUT_mem_MPORT_52_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_54_en & LUT_mem_MPORT_54_mask) begin
      LUT_mem[LUT_mem_MPORT_54_addr] <= LUT_mem_MPORT_54_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_56_en & LUT_mem_MPORT_56_mask) begin
      LUT_mem[LUT_mem_MPORT_56_addr] <= LUT_mem_MPORT_56_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_58_en & LUT_mem_MPORT_58_mask) begin
      LUT_mem[LUT_mem_MPORT_58_addr] <= LUT_mem_MPORT_58_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_60_en & LUT_mem_MPORT_60_mask) begin
      LUT_mem[LUT_mem_MPORT_60_addr] <= LUT_mem_MPORT_60_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_62_en & LUT_mem_MPORT_62_mask) begin
      LUT_mem[LUT_mem_MPORT_62_addr] <= LUT_mem_MPORT_62_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_64_en & LUT_mem_MPORT_64_mask) begin
      LUT_mem[LUT_mem_MPORT_64_addr] <= LUT_mem_MPORT_64_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_66_en & LUT_mem_MPORT_66_mask) begin
      LUT_mem[LUT_mem_MPORT_66_addr] <= LUT_mem_MPORT_66_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_68_en & LUT_mem_MPORT_68_mask) begin
      LUT_mem[LUT_mem_MPORT_68_addr] <= LUT_mem_MPORT_68_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_70_en & LUT_mem_MPORT_70_mask) begin
      LUT_mem[LUT_mem_MPORT_70_addr] <= LUT_mem_MPORT_70_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_72_en & LUT_mem_MPORT_72_mask) begin
      LUT_mem[LUT_mem_MPORT_72_addr] <= LUT_mem_MPORT_72_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_74_en & LUT_mem_MPORT_74_mask) begin
      LUT_mem[LUT_mem_MPORT_74_addr] <= LUT_mem_MPORT_74_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_76_en & LUT_mem_MPORT_76_mask) begin
      LUT_mem[LUT_mem_MPORT_76_addr] <= LUT_mem_MPORT_76_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_78_en & LUT_mem_MPORT_78_mask) begin
      LUT_mem[LUT_mem_MPORT_78_addr] <= LUT_mem_MPORT_78_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_80_en & LUT_mem_MPORT_80_mask) begin
      LUT_mem[LUT_mem_MPORT_80_addr] <= LUT_mem_MPORT_80_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_82_en & LUT_mem_MPORT_82_mask) begin
      LUT_mem[LUT_mem_MPORT_82_addr] <= LUT_mem_MPORT_82_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_84_en & LUT_mem_MPORT_84_mask) begin
      LUT_mem[LUT_mem_MPORT_84_addr] <= LUT_mem_MPORT_84_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_86_en & LUT_mem_MPORT_86_mask) begin
      LUT_mem[LUT_mem_MPORT_86_addr] <= LUT_mem_MPORT_86_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_88_en & LUT_mem_MPORT_88_mask) begin
      LUT_mem[LUT_mem_MPORT_88_addr] <= LUT_mem_MPORT_88_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_90_en & LUT_mem_MPORT_90_mask) begin
      LUT_mem[LUT_mem_MPORT_90_addr] <= LUT_mem_MPORT_90_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_92_en & LUT_mem_MPORT_92_mask) begin
      LUT_mem[LUT_mem_MPORT_92_addr] <= LUT_mem_MPORT_92_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_94_en & LUT_mem_MPORT_94_mask) begin
      LUT_mem[LUT_mem_MPORT_94_addr] <= LUT_mem_MPORT_94_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_96_en & LUT_mem_MPORT_96_mask) begin
      LUT_mem[LUT_mem_MPORT_96_addr] <= LUT_mem_MPORT_96_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_98_en & LUT_mem_MPORT_98_mask) begin
      LUT_mem[LUT_mem_MPORT_98_addr] <= LUT_mem_MPORT_98_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_100_en & LUT_mem_MPORT_100_mask) begin
      LUT_mem[LUT_mem_MPORT_100_addr] <= LUT_mem_MPORT_100_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_102_en & LUT_mem_MPORT_102_mask) begin
      LUT_mem[LUT_mem_MPORT_102_addr] <= LUT_mem_MPORT_102_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_104_en & LUT_mem_MPORT_104_mask) begin
      LUT_mem[LUT_mem_MPORT_104_addr] <= LUT_mem_MPORT_104_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_106_en & LUT_mem_MPORT_106_mask) begin
      LUT_mem[LUT_mem_MPORT_106_addr] <= LUT_mem_MPORT_106_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_108_en & LUT_mem_MPORT_108_mask) begin
      LUT_mem[LUT_mem_MPORT_108_addr] <= LUT_mem_MPORT_108_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_110_en & LUT_mem_MPORT_110_mask) begin
      LUT_mem[LUT_mem_MPORT_110_addr] <= LUT_mem_MPORT_110_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_112_en & LUT_mem_MPORT_112_mask) begin
      LUT_mem[LUT_mem_MPORT_112_addr] <= LUT_mem_MPORT_112_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_114_en & LUT_mem_MPORT_114_mask) begin
      LUT_mem[LUT_mem_MPORT_114_addr] <= LUT_mem_MPORT_114_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_116_en & LUT_mem_MPORT_116_mask) begin
      LUT_mem[LUT_mem_MPORT_116_addr] <= LUT_mem_MPORT_116_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_118_en & LUT_mem_MPORT_118_mask) begin
      LUT_mem[LUT_mem_MPORT_118_addr] <= LUT_mem_MPORT_118_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_120_en & LUT_mem_MPORT_120_mask) begin
      LUT_mem[LUT_mem_MPORT_120_addr] <= LUT_mem_MPORT_120_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_122_en & LUT_mem_MPORT_122_mask) begin
      LUT_mem[LUT_mem_MPORT_122_addr] <= LUT_mem_MPORT_122_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_124_en & LUT_mem_MPORT_124_mask) begin
      LUT_mem[LUT_mem_MPORT_124_addr] <= LUT_mem_MPORT_124_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_126_en & LUT_mem_MPORT_126_mask) begin
      LUT_mem[LUT_mem_MPORT_126_addr] <= LUT_mem_MPORT_126_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_128_en & LUT_mem_MPORT_128_mask) begin
      LUT_mem[LUT_mem_MPORT_128_addr] <= LUT_mem_MPORT_128_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_130_en & LUT_mem_MPORT_130_mask) begin
      LUT_mem[LUT_mem_MPORT_130_addr] <= LUT_mem_MPORT_130_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_132_en & LUT_mem_MPORT_132_mask) begin
      LUT_mem[LUT_mem_MPORT_132_addr] <= LUT_mem_MPORT_132_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_134_en & LUT_mem_MPORT_134_mask) begin
      LUT_mem[LUT_mem_MPORT_134_addr] <= LUT_mem_MPORT_134_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_136_en & LUT_mem_MPORT_136_mask) begin
      LUT_mem[LUT_mem_MPORT_136_addr] <= LUT_mem_MPORT_136_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_138_en & LUT_mem_MPORT_138_mask) begin
      LUT_mem[LUT_mem_MPORT_138_addr] <= LUT_mem_MPORT_138_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_211_en & LUT_mem_MPORT_211_mask) begin
      LUT_mem[LUT_mem_MPORT_211_addr] <= LUT_mem_MPORT_211_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_213_en & LUT_mem_MPORT_213_mask) begin
      LUT_mem[LUT_mem_MPORT_213_addr] <= LUT_mem_MPORT_213_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_215_en & LUT_mem_MPORT_215_mask) begin
      LUT_mem[LUT_mem_MPORT_215_addr] <= LUT_mem_MPORT_215_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_217_en & LUT_mem_MPORT_217_mask) begin
      LUT_mem[LUT_mem_MPORT_217_addr] <= LUT_mem_MPORT_217_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_219_en & LUT_mem_MPORT_219_mask) begin
      LUT_mem[LUT_mem_MPORT_219_addr] <= LUT_mem_MPORT_219_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_221_en & LUT_mem_MPORT_221_mask) begin
      LUT_mem[LUT_mem_MPORT_221_addr] <= LUT_mem_MPORT_221_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_223_en & LUT_mem_MPORT_223_mask) begin
      LUT_mem[LUT_mem_MPORT_223_addr] <= LUT_mem_MPORT_223_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_225_en & LUT_mem_MPORT_225_mask) begin
      LUT_mem[LUT_mem_MPORT_225_addr] <= LUT_mem_MPORT_225_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_227_en & LUT_mem_MPORT_227_mask) begin
      LUT_mem[LUT_mem_MPORT_227_addr] <= LUT_mem_MPORT_227_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_229_en & LUT_mem_MPORT_229_mask) begin
      LUT_mem[LUT_mem_MPORT_229_addr] <= LUT_mem_MPORT_229_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_231_en & LUT_mem_MPORT_231_mask) begin
      LUT_mem[LUT_mem_MPORT_231_addr] <= LUT_mem_MPORT_231_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_233_en & LUT_mem_MPORT_233_mask) begin
      LUT_mem[LUT_mem_MPORT_233_addr] <= LUT_mem_MPORT_233_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_235_en & LUT_mem_MPORT_235_mask) begin
      LUT_mem[LUT_mem_MPORT_235_addr] <= LUT_mem_MPORT_235_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_237_en & LUT_mem_MPORT_237_mask) begin
      LUT_mem[LUT_mem_MPORT_237_addr] <= LUT_mem_MPORT_237_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_239_en & LUT_mem_MPORT_239_mask) begin
      LUT_mem[LUT_mem_MPORT_239_addr] <= LUT_mem_MPORT_239_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_241_en & LUT_mem_MPORT_241_mask) begin
      LUT_mem[LUT_mem_MPORT_241_addr] <= LUT_mem_MPORT_241_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_243_en & LUT_mem_MPORT_243_mask) begin
      LUT_mem[LUT_mem_MPORT_243_addr] <= LUT_mem_MPORT_243_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_245_en & LUT_mem_MPORT_245_mask) begin
      LUT_mem[LUT_mem_MPORT_245_addr] <= LUT_mem_MPORT_245_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_247_en & LUT_mem_MPORT_247_mask) begin
      LUT_mem[LUT_mem_MPORT_247_addr] <= LUT_mem_MPORT_247_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_249_en & LUT_mem_MPORT_249_mask) begin
      LUT_mem[LUT_mem_MPORT_249_addr] <= LUT_mem_MPORT_249_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_251_en & LUT_mem_MPORT_251_mask) begin
      LUT_mem[LUT_mem_MPORT_251_addr] <= LUT_mem_MPORT_251_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_253_en & LUT_mem_MPORT_253_mask) begin
      LUT_mem[LUT_mem_MPORT_253_addr] <= LUT_mem_MPORT_253_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_255_en & LUT_mem_MPORT_255_mask) begin
      LUT_mem[LUT_mem_MPORT_255_addr] <= LUT_mem_MPORT_255_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_257_en & LUT_mem_MPORT_257_mask) begin
      LUT_mem[LUT_mem_MPORT_257_addr] <= LUT_mem_MPORT_257_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_259_en & LUT_mem_MPORT_259_mask) begin
      LUT_mem[LUT_mem_MPORT_259_addr] <= LUT_mem_MPORT_259_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_261_en & LUT_mem_MPORT_261_mask) begin
      LUT_mem[LUT_mem_MPORT_261_addr] <= LUT_mem_MPORT_261_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_263_en & LUT_mem_MPORT_263_mask) begin
      LUT_mem[LUT_mem_MPORT_263_addr] <= LUT_mem_MPORT_263_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_265_en & LUT_mem_MPORT_265_mask) begin
      LUT_mem[LUT_mem_MPORT_265_addr] <= LUT_mem_MPORT_265_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_267_en & LUT_mem_MPORT_267_mask) begin
      LUT_mem[LUT_mem_MPORT_267_addr] <= LUT_mem_MPORT_267_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_269_en & LUT_mem_MPORT_269_mask) begin
      LUT_mem[LUT_mem_MPORT_269_addr] <= LUT_mem_MPORT_269_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_271_en & LUT_mem_MPORT_271_mask) begin
      LUT_mem[LUT_mem_MPORT_271_addr] <= LUT_mem_MPORT_271_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_273_en & LUT_mem_MPORT_273_mask) begin
      LUT_mem[LUT_mem_MPORT_273_addr] <= LUT_mem_MPORT_273_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_275_en & LUT_mem_MPORT_275_mask) begin
      LUT_mem[LUT_mem_MPORT_275_addr] <= LUT_mem_MPORT_275_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_277_en & LUT_mem_MPORT_277_mask) begin
      LUT_mem[LUT_mem_MPORT_277_addr] <= LUT_mem_MPORT_277_data; // @[lut_35.scala 177:26]
    end
    if(LUT_mem_MPORT_279_en & LUT_mem_MPORT_279_mask) begin
      LUT_mem[LUT_mem_MPORT_279_addr] <= LUT_mem_MPORT_279_data; // @[lut_35.scala 177:26]
    end
    if (reset) begin // @[lut_35.scala 178:30]
      read_stack0 <= 32'h0; // @[lut_35.scala 178:30]
    end else begin
      read_stack0 <= LUT_mem_MPORT_140_data[31:0]; // @[lut_35.scala 550:26]
    end
    if (reset) begin // @[lut_35.scala 179:30]
      read_stack1 <= 32'h0; // @[lut_35.scala 179:30]
    end else begin
      read_stack1 <= LUT_mem_MPORT_141_data[31:0]; // @[lut_35.scala 551:26]
    end
    if (reset) begin // @[lut_35.scala 180:30]
      read_stack2 <= 32'h0; // @[lut_35.scala 180:30]
    end else begin
      read_stack2 <= LUT_mem_MPORT_142_data[31:0]; // @[lut_35.scala 552:26]
    end
    if (reset) begin // @[lut_35.scala 181:30]
      read_stack3 <= 32'h0; // @[lut_35.scala 181:30]
    end else begin
      read_stack3 <= LUT_mem_MPORT_143_data[31:0]; // @[lut_35.scala 553:26]
    end
    if (reset) begin // @[lut_35.scala 182:30]
      read_stack4 <= 32'h0; // @[lut_35.scala 182:30]
    end else begin
      read_stack4 <= LUT_mem_MPORT_144_data[31:0]; // @[lut_35.scala 554:26]
    end
    if (reset) begin // @[lut_35.scala 183:30]
      read_stack5 <= 32'h0; // @[lut_35.scala 183:30]
    end else begin
      read_stack5 <= LUT_mem_MPORT_145_data[31:0]; // @[lut_35.scala 555:26]
    end
    if (reset) begin // @[lut_35.scala 184:30]
      read_stack6 <= 32'h0; // @[lut_35.scala 184:30]
    end else begin
      read_stack6 <= LUT_mem_MPORT_146_data[31:0]; // @[lut_35.scala 556:26]
    end
    if (reset) begin // @[lut_35.scala 185:30]
      read_stack7 <= 32'h0; // @[lut_35.scala 185:30]
    end else begin
      read_stack7 <= LUT_mem_MPORT_147_data[31:0]; // @[lut_35.scala 557:26]
    end
    if (reset) begin // @[lut_35.scala 186:30]
      read_stack8 <= 32'h0; // @[lut_35.scala 186:30]
    end else begin
      read_stack8 <= LUT_mem_MPORT_148_data[31:0]; // @[lut_35.scala 558:26]
    end
    if (reset) begin // @[lut_35.scala 187:30]
      read_stack9 <= 32'h0; // @[lut_35.scala 187:30]
    end else begin
      read_stack9 <= LUT_mem_MPORT_149_data[31:0]; // @[lut_35.scala 559:26]
    end
    if (reset) begin // @[lut_35.scala 188:31]
      read_stack10 <= 32'h0; // @[lut_35.scala 188:31]
    end else begin
      read_stack10 <= LUT_mem_MPORT_150_data[31:0]; // @[lut_35.scala 560:27]
    end
    if (reset) begin // @[lut_35.scala 189:31]
      read_stack11 <= 32'h0; // @[lut_35.scala 189:31]
    end else begin
      read_stack11 <= LUT_mem_MPORT_151_data[31:0]; // @[lut_35.scala 561:27]
    end
    if (reset) begin // @[lut_35.scala 190:31]
      read_stack12 <= 32'h0; // @[lut_35.scala 190:31]
    end else begin
      read_stack12 <= LUT_mem_MPORT_152_data[31:0]; // @[lut_35.scala 562:27]
    end
    if (reset) begin // @[lut_35.scala 191:31]
      read_stack13 <= 32'h0; // @[lut_35.scala 191:31]
    end else begin
      read_stack13 <= LUT_mem_MPORT_153_data[31:0]; // @[lut_35.scala 563:27]
    end
    if (reset) begin // @[lut_35.scala 192:31]
      read_stack14 <= 32'h0; // @[lut_35.scala 192:31]
    end else begin
      read_stack14 <= LUT_mem_MPORT_154_data[31:0]; // @[lut_35.scala 564:27]
    end
    if (reset) begin // @[lut_35.scala 193:31]
      read_stack15 <= 32'h0; // @[lut_35.scala 193:31]
    end else begin
      read_stack15 <= LUT_mem_MPORT_155_data[31:0]; // @[lut_35.scala 565:27]
    end
    if (reset) begin // @[lut_35.scala 194:31]
      read_stack16 <= 32'h0; // @[lut_35.scala 194:31]
    end else begin
      read_stack16 <= LUT_mem_MPORT_156_data[31:0]; // @[lut_35.scala 566:27]
    end
    if (reset) begin // @[lut_35.scala 195:31]
      read_stack17 <= 32'h0; // @[lut_35.scala 195:31]
    end else begin
      read_stack17 <= LUT_mem_MPORT_157_data[31:0]; // @[lut_35.scala 567:27]
    end
    if (reset) begin // @[lut_35.scala 196:31]
      read_stack18 <= 32'h0; // @[lut_35.scala 196:31]
    end else begin
      read_stack18 <= LUT_mem_MPORT_158_data[31:0]; // @[lut_35.scala 568:27]
    end
    if (reset) begin // @[lut_35.scala 197:31]
      read_stack19 <= 32'h0; // @[lut_35.scala 197:31]
    end else begin
      read_stack19 <= LUT_mem_MPORT_159_data[31:0]; // @[lut_35.scala 569:27]
    end
    if (reset) begin // @[lut_35.scala 198:31]
      read_stack20 <= 32'h0; // @[lut_35.scala 198:31]
    end else begin
      read_stack20 <= LUT_mem_MPORT_160_data[31:0]; // @[lut_35.scala 570:27]
    end
    if (reset) begin // @[lut_35.scala 199:31]
      read_stack21 <= 32'h0; // @[lut_35.scala 199:31]
    end else begin
      read_stack21 <= LUT_mem_MPORT_161_data[31:0]; // @[lut_35.scala 571:27]
    end
    if (reset) begin // @[lut_35.scala 200:31]
      read_stack22 <= 32'h0; // @[lut_35.scala 200:31]
    end else begin
      read_stack22 <= LUT_mem_MPORT_162_data[31:0]; // @[lut_35.scala 572:27]
    end
    if (reset) begin // @[lut_35.scala 201:31]
      read_stack23 <= 32'h0; // @[lut_35.scala 201:31]
    end else begin
      read_stack23 <= LUT_mem_MPORT_163_data[31:0]; // @[lut_35.scala 573:27]
    end
    if (reset) begin // @[lut_35.scala 202:31]
      read_stack24 <= 32'h0; // @[lut_35.scala 202:31]
    end else begin
      read_stack24 <= LUT_mem_MPORT_164_data[31:0]; // @[lut_35.scala 574:27]
    end
    if (reset) begin // @[lut_35.scala 203:31]
      read_stack25 <= 32'h0; // @[lut_35.scala 203:31]
    end else begin
      read_stack25 <= LUT_mem_MPORT_165_data[31:0]; // @[lut_35.scala 575:27]
    end
    if (reset) begin // @[lut_35.scala 204:31]
      read_stack26 <= 32'h0; // @[lut_35.scala 204:31]
    end else begin
      read_stack26 <= LUT_mem_MPORT_166_data[31:0]; // @[lut_35.scala 576:27]
    end
    if (reset) begin // @[lut_35.scala 205:31]
      read_stack27 <= 32'h0; // @[lut_35.scala 205:31]
    end else begin
      read_stack27 <= LUT_mem_MPORT_167_data[31:0]; // @[lut_35.scala 577:27]
    end
    if (reset) begin // @[lut_35.scala 206:31]
      read_stack28 <= 32'h0; // @[lut_35.scala 206:31]
    end else begin
      read_stack28 <= LUT_mem_MPORT_168_data[31:0]; // @[lut_35.scala 578:27]
    end
    if (reset) begin // @[lut_35.scala 207:31]
      read_stack29 <= 32'h0; // @[lut_35.scala 207:31]
    end else begin
      read_stack29 <= LUT_mem_MPORT_169_data[31:0]; // @[lut_35.scala 579:27]
    end
    if (reset) begin // @[lut_35.scala 208:31]
      read_stack30 <= 32'h0; // @[lut_35.scala 208:31]
    end else begin
      read_stack30 <= LUT_mem_MPORT_170_data[31:0]; // @[lut_35.scala 580:27]
    end
    if (reset) begin // @[lut_35.scala 209:31]
      read_stack31 <= 32'h0; // @[lut_35.scala 209:31]
    end else begin
      read_stack31 <= LUT_mem_MPORT_171_data[31:0]; // @[lut_35.scala 581:27]
    end
    if (reset) begin // @[lut_35.scala 210:31]
      read_stack32 <= 32'h0; // @[lut_35.scala 210:31]
    end else begin
      read_stack32 <= LUT_mem_MPORT_172_data[31:0]; // @[lut_35.scala 582:27]
    end
    if (reset) begin // @[lut_35.scala 211:31]
      read_stack33 <= 32'h0; // @[lut_35.scala 211:31]
    end else begin
      read_stack33 <= LUT_mem_MPORT_173_data[31:0]; // @[lut_35.scala 583:27]
    end
    if (reset) begin // @[lut_35.scala 212:31]
      read_stack34 <= 32'h0; // @[lut_35.scala 212:31]
    end else begin
      read_stack34 <= LUT_mem_MPORT_174_data[31:0]; // @[lut_35.scala 584:27]
    end
    if (reset) begin // @[lut_35.scala 214:31]
      push_0_1 <= 1'h0; // @[lut_35.scala 214:31]
    end else begin
      push_0_1 <= _GEN_19146;
    end
    if (reset) begin // @[lut_35.scala 215:31]
      push_1_1 <= 1'h0; // @[lut_35.scala 215:31]
    end else begin
      push_1_1 <= _GEN_19147;
    end
    if (reset) begin // @[lut_35.scala 216:31]
      push_2_1 <= 1'h0; // @[lut_35.scala 216:31]
    end else begin
      push_2_1 <= _GEN_19148;
    end
    if (reset) begin // @[lut_35.scala 217:31]
      push_3_1 <= 1'h0; // @[lut_35.scala 217:31]
    end else begin
      push_3_1 <= _GEN_19149;
    end
    if (reset) begin // @[lut_35.scala 218:31]
      push_4_1 <= 1'h0; // @[lut_35.scala 218:31]
    end else begin
      push_4_1 <= _GEN_19150;
    end
    if (reset) begin // @[lut_35.scala 219:31]
      push_5_1 <= 1'h0; // @[lut_35.scala 219:31]
    end else begin
      push_5_1 <= _GEN_19151;
    end
    if (reset) begin // @[lut_35.scala 220:31]
      push_6_1 <= 1'h0; // @[lut_35.scala 220:31]
    end else begin
      push_6_1 <= _GEN_19152;
    end
    if (reset) begin // @[lut_35.scala 221:31]
      push_7_1 <= 1'h0; // @[lut_35.scala 221:31]
    end else begin
      push_7_1 <= _GEN_19153;
    end
    if (reset) begin // @[lut_35.scala 222:31]
      push_8_1 <= 1'h0; // @[lut_35.scala 222:31]
    end else begin
      push_8_1 <= _GEN_19154;
    end
    if (reset) begin // @[lut_35.scala 223:31]
      push_9_1 <= 1'h0; // @[lut_35.scala 223:31]
    end else begin
      push_9_1 <= _GEN_19155;
    end
    if (reset) begin // @[lut_35.scala 224:32]
      push_10_1 <= 1'h0; // @[lut_35.scala 224:32]
    end else begin
      push_10_1 <= _GEN_19156;
    end
    if (reset) begin // @[lut_35.scala 225:32]
      push_11_1 <= 1'h0; // @[lut_35.scala 225:32]
    end else begin
      push_11_1 <= _GEN_19157;
    end
    if (reset) begin // @[lut_35.scala 226:32]
      push_12_1 <= 1'h0; // @[lut_35.scala 226:32]
    end else begin
      push_12_1 <= _GEN_19158;
    end
    if (reset) begin // @[lut_35.scala 227:32]
      push_13_1 <= 1'h0; // @[lut_35.scala 227:32]
    end else begin
      push_13_1 <= _GEN_19159;
    end
    if (reset) begin // @[lut_35.scala 228:32]
      push_14_1 <= 1'h0; // @[lut_35.scala 228:32]
    end else begin
      push_14_1 <= _GEN_19160;
    end
    if (reset) begin // @[lut_35.scala 229:32]
      push_15_1 <= 1'h0; // @[lut_35.scala 229:32]
    end else begin
      push_15_1 <= _GEN_19161;
    end
    if (reset) begin // @[lut_35.scala 230:32]
      push_16_1 <= 1'h0; // @[lut_35.scala 230:32]
    end else begin
      push_16_1 <= _GEN_19162;
    end
    if (reset) begin // @[lut_35.scala 231:32]
      push_17_1 <= 1'h0; // @[lut_35.scala 231:32]
    end else begin
      push_17_1 <= _GEN_19163;
    end
    if (reset) begin // @[lut_35.scala 232:32]
      push_18_1 <= 1'h0; // @[lut_35.scala 232:32]
    end else begin
      push_18_1 <= _GEN_19164;
    end
    if (reset) begin // @[lut_35.scala 233:32]
      push_19_1 <= 1'h0; // @[lut_35.scala 233:32]
    end else begin
      push_19_1 <= _GEN_19165;
    end
    if (reset) begin // @[lut_35.scala 234:32]
      push_20_1 <= 1'h0; // @[lut_35.scala 234:32]
    end else begin
      push_20_1 <= _GEN_19166;
    end
    if (reset) begin // @[lut_35.scala 235:32]
      push_21_1 <= 1'h0; // @[lut_35.scala 235:32]
    end else begin
      push_21_1 <= _GEN_19167;
    end
    if (reset) begin // @[lut_35.scala 236:32]
      push_22_1 <= 1'h0; // @[lut_35.scala 236:32]
    end else begin
      push_22_1 <= _GEN_19168;
    end
    if (reset) begin // @[lut_35.scala 237:32]
      push_23_1 <= 1'h0; // @[lut_35.scala 237:32]
    end else begin
      push_23_1 <= _GEN_19169;
    end
    if (reset) begin // @[lut_35.scala 238:32]
      push_24_1 <= 1'h0; // @[lut_35.scala 238:32]
    end else begin
      push_24_1 <= _GEN_19170;
    end
    if (reset) begin // @[lut_35.scala 239:32]
      push_25_1 <= 1'h0; // @[lut_35.scala 239:32]
    end else begin
      push_25_1 <= _GEN_19171;
    end
    if (reset) begin // @[lut_35.scala 240:32]
      push_26_1 <= 1'h0; // @[lut_35.scala 240:32]
    end else begin
      push_26_1 <= _GEN_19172;
    end
    if (reset) begin // @[lut_35.scala 241:32]
      push_27_1 <= 1'h0; // @[lut_35.scala 241:32]
    end else begin
      push_27_1 <= _GEN_19173;
    end
    if (reset) begin // @[lut_35.scala 242:32]
      push_28_1 <= 1'h0; // @[lut_35.scala 242:32]
    end else begin
      push_28_1 <= _GEN_19174;
    end
    if (reset) begin // @[lut_35.scala 243:32]
      push_29_1 <= 1'h0; // @[lut_35.scala 243:32]
    end else begin
      push_29_1 <= _GEN_19175;
    end
    if (reset) begin // @[lut_35.scala 244:32]
      push_30_1 <= 1'h0; // @[lut_35.scala 244:32]
    end else begin
      push_30_1 <= _GEN_19176;
    end
    if (reset) begin // @[lut_35.scala 245:32]
      push_31_1 <= 1'h0; // @[lut_35.scala 245:32]
    end else begin
      push_31_1 <= _GEN_19177;
    end
    if (reset) begin // @[lut_35.scala 246:32]
      push_32_1 <= 1'h0; // @[lut_35.scala 246:32]
    end else begin
      push_32_1 <= _GEN_19178;
    end
    if (reset) begin // @[lut_35.scala 247:32]
      push_33_1 <= 1'h0; // @[lut_35.scala 247:32]
    end else begin
      push_33_1 <= _GEN_19179;
    end
    if (reset) begin // @[lut_35.scala 248:32]
      push_34_1 <= 1'h0; // @[lut_35.scala 248:32]
    end else begin
      push_34_1 <= _GEN_19180;
    end
    if (reset) begin // @[lut_35.scala 252:40]
      push_1 <= 1'h0; // @[lut_35.scala 252:40]
    end else begin
      push_1 <= _T_106;
    end
    if (reset) begin // @[lut_35.scala 253:41]
      push_valid <= 1'h0; // @[lut_35.scala 253:41]
    end else begin
      push_valid <= _GEN_351;
    end
    if (reset) begin // @[lut_35.scala 255:41]
      push_ray_id <= 32'h0; // @[lut_35.scala 255:41]
    end else if (io_push & io_push_valid) begin // @[lut_35.scala 596:46]
      push_ray_id <= io_ray_id_push; // @[lut_35.scala 600:26]
    end
    if (reset) begin // @[lut_35.scala 295:41]
      push_valid_2 <= 1'h0; // @[lut_35.scala 295:41]
    end else begin
      push_valid_2 <= _GEN_19181;
    end
    if (reset) begin // @[lut_35.scala 3532:50]
      pop_1 <= 1'h0; // @[lut_35.scala 3532:50]
    end else begin
      pop_1 <= _T_672;
    end
    if (reset) begin // @[lut_35.scala 3533:38]
      read_stack0_pop <= 32'h0; // @[lut_35.scala 3533:38]
    end else begin
      read_stack0_pop <= LUT_mem_MPORT_280_data[31:0]; // @[lut_35.scala 3618:30]
    end
    if (reset) begin // @[lut_35.scala 3534:38]
      read_stack1_pop <= 32'h0; // @[lut_35.scala 3534:38]
    end else begin
      read_stack1_pop <= LUT_mem_MPORT_281_data[31:0]; // @[lut_35.scala 3619:30]
    end
    if (reset) begin // @[lut_35.scala 3535:38]
      read_stack2_pop <= 32'h0; // @[lut_35.scala 3535:38]
    end else begin
      read_stack2_pop <= LUT_mem_MPORT_282_data[31:0]; // @[lut_35.scala 3620:30]
    end
    if (reset) begin // @[lut_35.scala 3536:38]
      read_stack3_pop <= 32'h0; // @[lut_35.scala 3536:38]
    end else begin
      read_stack3_pop <= LUT_mem_MPORT_283_data[31:0]; // @[lut_35.scala 3621:30]
    end
    if (reset) begin // @[lut_35.scala 3537:38]
      read_stack4_pop <= 32'h0; // @[lut_35.scala 3537:38]
    end else begin
      read_stack4_pop <= LUT_mem_MPORT_284_data[31:0]; // @[lut_35.scala 3622:30]
    end
    if (reset) begin // @[lut_35.scala 3538:38]
      read_stack5_pop <= 32'h0; // @[lut_35.scala 3538:38]
    end else begin
      read_stack5_pop <= LUT_mem_MPORT_285_data[31:0]; // @[lut_35.scala 3623:30]
    end
    if (reset) begin // @[lut_35.scala 3539:38]
      read_stack6_pop <= 32'h0; // @[lut_35.scala 3539:38]
    end else begin
      read_stack6_pop <= LUT_mem_MPORT_286_data[31:0]; // @[lut_35.scala 3624:30]
    end
    if (reset) begin // @[lut_35.scala 3540:38]
      read_stack7_pop <= 32'h0; // @[lut_35.scala 3540:38]
    end else begin
      read_stack7_pop <= LUT_mem_MPORT_287_data[31:0]; // @[lut_35.scala 3625:30]
    end
    if (reset) begin // @[lut_35.scala 3541:38]
      read_stack8_pop <= 32'h0; // @[lut_35.scala 3541:38]
    end else begin
      read_stack8_pop <= LUT_mem_MPORT_288_data[31:0]; // @[lut_35.scala 3626:30]
    end
    if (reset) begin // @[lut_35.scala 3542:38]
      read_stack9_pop <= 32'h0; // @[lut_35.scala 3542:38]
    end else begin
      read_stack9_pop <= LUT_mem_MPORT_289_data[31:0]; // @[lut_35.scala 3627:30]
    end
    if (reset) begin // @[lut_35.scala 3543:39]
      read_stack10_pop <= 32'h0; // @[lut_35.scala 3543:39]
    end else begin
      read_stack10_pop <= LUT_mem_MPORT_290_data[31:0]; // @[lut_35.scala 3629:31]
    end
    if (reset) begin // @[lut_35.scala 3544:39]
      read_stack11_pop <= 32'h0; // @[lut_35.scala 3544:39]
    end else begin
      read_stack11_pop <= LUT_mem_MPORT_291_data[31:0]; // @[lut_35.scala 3630:31]
    end
    if (reset) begin // @[lut_35.scala 3545:39]
      read_stack12_pop <= 32'h0; // @[lut_35.scala 3545:39]
    end else begin
      read_stack12_pop <= LUT_mem_MPORT_292_data[31:0]; // @[lut_35.scala 3631:31]
    end
    if (reset) begin // @[lut_35.scala 3546:39]
      read_stack13_pop <= 32'h0; // @[lut_35.scala 3546:39]
    end else begin
      read_stack13_pop <= LUT_mem_MPORT_293_data[31:0]; // @[lut_35.scala 3632:31]
    end
    if (reset) begin // @[lut_35.scala 3547:39]
      read_stack14_pop <= 32'h0; // @[lut_35.scala 3547:39]
    end else begin
      read_stack14_pop <= LUT_mem_MPORT_294_data[31:0]; // @[lut_35.scala 3633:31]
    end
    if (reset) begin // @[lut_35.scala 3548:39]
      read_stack15_pop <= 32'h0; // @[lut_35.scala 3548:39]
    end else begin
      read_stack15_pop <= LUT_mem_MPORT_295_data[31:0]; // @[lut_35.scala 3634:31]
    end
    if (reset) begin // @[lut_35.scala 3549:39]
      read_stack16_pop <= 32'h0; // @[lut_35.scala 3549:39]
    end else begin
      read_stack16_pop <= LUT_mem_MPORT_296_data[31:0]; // @[lut_35.scala 3635:31]
    end
    if (reset) begin // @[lut_35.scala 3550:39]
      read_stack17_pop <= 32'h0; // @[lut_35.scala 3550:39]
    end else begin
      read_stack17_pop <= LUT_mem_MPORT_297_data[31:0]; // @[lut_35.scala 3636:31]
    end
    if (reset) begin // @[lut_35.scala 3551:39]
      read_stack18_pop <= 32'h0; // @[lut_35.scala 3551:39]
    end else begin
      read_stack18_pop <= LUT_mem_MPORT_298_data[31:0]; // @[lut_35.scala 3637:31]
    end
    if (reset) begin // @[lut_35.scala 3552:39]
      read_stack19_pop <= 32'h0; // @[lut_35.scala 3552:39]
    end else begin
      read_stack19_pop <= LUT_mem_MPORT_299_data[31:0]; // @[lut_35.scala 3638:31]
    end
    if (reset) begin // @[lut_35.scala 3553:39]
      read_stack20_pop <= 32'h0; // @[lut_35.scala 3553:39]
    end else begin
      read_stack20_pop <= LUT_mem_MPORT_300_data[31:0]; // @[lut_35.scala 3640:31]
    end
    if (reset) begin // @[lut_35.scala 3554:39]
      read_stack21_pop <= 32'h0; // @[lut_35.scala 3554:39]
    end else begin
      read_stack21_pop <= LUT_mem_MPORT_301_data[31:0]; // @[lut_35.scala 3641:31]
    end
    if (reset) begin // @[lut_35.scala 3555:39]
      read_stack22_pop <= 32'h0; // @[lut_35.scala 3555:39]
    end else begin
      read_stack22_pop <= LUT_mem_MPORT_302_data[31:0]; // @[lut_35.scala 3642:31]
    end
    if (reset) begin // @[lut_35.scala 3556:39]
      read_stack23_pop <= 32'h0; // @[lut_35.scala 3556:39]
    end else begin
      read_stack23_pop <= LUT_mem_MPORT_303_data[31:0]; // @[lut_35.scala 3643:31]
    end
    if (reset) begin // @[lut_35.scala 3557:39]
      read_stack24_pop <= 32'h0; // @[lut_35.scala 3557:39]
    end else begin
      read_stack24_pop <= LUT_mem_MPORT_304_data[31:0]; // @[lut_35.scala 3644:31]
    end
    if (reset) begin // @[lut_35.scala 3558:39]
      read_stack25_pop <= 32'h0; // @[lut_35.scala 3558:39]
    end else begin
      read_stack25_pop <= LUT_mem_MPORT_305_data[31:0]; // @[lut_35.scala 3645:31]
    end
    if (reset) begin // @[lut_35.scala 3559:39]
      read_stack26_pop <= 32'h0; // @[lut_35.scala 3559:39]
    end else begin
      read_stack26_pop <= LUT_mem_MPORT_306_data[31:0]; // @[lut_35.scala 3646:31]
    end
    if (reset) begin // @[lut_35.scala 3560:39]
      read_stack27_pop <= 32'h0; // @[lut_35.scala 3560:39]
    end else begin
      read_stack27_pop <= LUT_mem_MPORT_307_data[31:0]; // @[lut_35.scala 3647:31]
    end
    if (reset) begin // @[lut_35.scala 3561:39]
      read_stack28_pop <= 32'h0; // @[lut_35.scala 3561:39]
    end else begin
      read_stack28_pop <= LUT_mem_MPORT_308_data[31:0]; // @[lut_35.scala 3648:31]
    end
    if (reset) begin // @[lut_35.scala 3562:39]
      read_stack29_pop <= 32'h0; // @[lut_35.scala 3562:39]
    end else begin
      read_stack29_pop <= LUT_mem_MPORT_309_data[31:0]; // @[lut_35.scala 3649:31]
    end
    if (reset) begin // @[lut_35.scala 3563:39]
      read_stack30_pop <= 32'h0; // @[lut_35.scala 3563:39]
    end else begin
      read_stack30_pop <= LUT_mem_MPORT_310_data[31:0]; // @[lut_35.scala 3651:31]
    end
    if (reset) begin // @[lut_35.scala 3564:39]
      read_stack31_pop <= 32'h0; // @[lut_35.scala 3564:39]
    end else begin
      read_stack31_pop <= LUT_mem_MPORT_311_data[31:0]; // @[lut_35.scala 3652:31]
    end
    if (reset) begin // @[lut_35.scala 3565:39]
      read_stack32_pop <= 32'h0; // @[lut_35.scala 3565:39]
    end else begin
      read_stack32_pop <= LUT_mem_MPORT_312_data[31:0]; // @[lut_35.scala 3653:31]
    end
    if (reset) begin // @[lut_35.scala 3566:39]
      read_stack33_pop <= 32'h0; // @[lut_35.scala 3566:39]
    end else begin
      read_stack33_pop <= LUT_mem_MPORT_313_data[31:0]; // @[lut_35.scala 3654:31]
    end
    if (reset) begin // @[lut_35.scala 3567:39]
      read_stack34_pop <= 32'h0; // @[lut_35.scala 3567:39]
    end else begin
      read_stack34_pop <= LUT_mem_MPORT_314_data[31:0]; // @[lut_35.scala 3655:31]
    end
    if (reset) begin // @[lut_35.scala 3570:37]
      pop_ray_id <= 32'h0; // @[lut_35.scala 3570:37]
    end else if (io_pop & io_pop_valid) begin // @[lut_35.scala 3657:44]
      pop_ray_id <= io_ray_id_pop; // @[lut_35.scala 3662:26]
    end
    if (reset) begin // @[lut_35.scala 3571:37]
      pop_hitT_1 <= 32'h0; // @[lut_35.scala 3571:37]
    end else if (io_pop & io_pop_valid) begin // @[lut_35.scala 3657:44]
      pop_hitT_1 <= io_hitT_in; // @[lut_35.scala 3663:26]
    end
    if (reset) begin // @[lut_35.scala 3572:36]
      pop_valid <= 1'h0; // @[lut_35.scala 3572:36]
    end else begin
      pop_valid <= _T_672;
    end
    if (reset) begin // @[lut_35.scala 3575:46]
      pop_0_1 <= 1'h0; // @[lut_35.scala 3575:46]
    end else begin
      pop_0_1 <= _GEN_20372;
    end
    if (reset) begin // @[lut_35.scala 3576:46]
      pop_1_1 <= 1'h0; // @[lut_35.scala 3576:46]
    end else begin
      pop_1_1 <= _GEN_20373;
    end
    if (reset) begin // @[lut_35.scala 3577:46]
      pop_2_1 <= 1'h0; // @[lut_35.scala 3577:46]
    end else begin
      pop_2_1 <= _GEN_20374;
    end
    if (reset) begin // @[lut_35.scala 3578:46]
      pop_3_1 <= 1'h0; // @[lut_35.scala 3578:46]
    end else begin
      pop_3_1 <= _GEN_20375;
    end
    if (reset) begin // @[lut_35.scala 3579:46]
      pop_4_1 <= 1'h0; // @[lut_35.scala 3579:46]
    end else begin
      pop_4_1 <= _GEN_20376;
    end
    if (reset) begin // @[lut_35.scala 3580:46]
      pop_5_1 <= 1'h0; // @[lut_35.scala 3580:46]
    end else begin
      pop_5_1 <= _GEN_20377;
    end
    if (reset) begin // @[lut_35.scala 3581:46]
      pop_6_1 <= 1'h0; // @[lut_35.scala 3581:46]
    end else begin
      pop_6_1 <= _GEN_20378;
    end
    if (reset) begin // @[lut_35.scala 3582:46]
      pop_7_1 <= 1'h0; // @[lut_35.scala 3582:46]
    end else begin
      pop_7_1 <= _GEN_20379;
    end
    if (reset) begin // @[lut_35.scala 3583:46]
      pop_8_1 <= 1'h0; // @[lut_35.scala 3583:46]
    end else begin
      pop_8_1 <= _GEN_20380;
    end
    if (reset) begin // @[lut_35.scala 3584:46]
      pop_9_1 <= 1'h0; // @[lut_35.scala 3584:46]
    end else begin
      pop_9_1 <= _GEN_20381;
    end
    if (reset) begin // @[lut_35.scala 3585:47]
      pop_10_1 <= 1'h0; // @[lut_35.scala 3585:47]
    end else begin
      pop_10_1 <= _GEN_20382;
    end
    if (reset) begin // @[lut_35.scala 3586:47]
      pop_11_1 <= 1'h0; // @[lut_35.scala 3586:47]
    end else begin
      pop_11_1 <= _GEN_20383;
    end
    if (reset) begin // @[lut_35.scala 3587:47]
      pop_12_1 <= 1'h0; // @[lut_35.scala 3587:47]
    end else begin
      pop_12_1 <= _GEN_20384;
    end
    if (reset) begin // @[lut_35.scala 3588:47]
      pop_13_1 <= 1'h0; // @[lut_35.scala 3588:47]
    end else begin
      pop_13_1 <= _GEN_20385;
    end
    if (reset) begin // @[lut_35.scala 3589:47]
      pop_14_1 <= 1'h0; // @[lut_35.scala 3589:47]
    end else begin
      pop_14_1 <= _GEN_20386;
    end
    if (reset) begin // @[lut_35.scala 3590:47]
      pop_15_1 <= 1'h0; // @[lut_35.scala 3590:47]
    end else begin
      pop_15_1 <= _GEN_20387;
    end
    if (reset) begin // @[lut_35.scala 3591:47]
      pop_16_1 <= 1'h0; // @[lut_35.scala 3591:47]
    end else begin
      pop_16_1 <= _GEN_20388;
    end
    if (reset) begin // @[lut_35.scala 3592:47]
      pop_17_1 <= 1'h0; // @[lut_35.scala 3592:47]
    end else begin
      pop_17_1 <= _GEN_20389;
    end
    if (reset) begin // @[lut_35.scala 3593:47]
      pop_18_1 <= 1'h0; // @[lut_35.scala 3593:47]
    end else begin
      pop_18_1 <= _GEN_20390;
    end
    if (reset) begin // @[lut_35.scala 3594:47]
      pop_19_1 <= 1'h0; // @[lut_35.scala 3594:47]
    end else begin
      pop_19_1 <= _GEN_20391;
    end
    if (reset) begin // @[lut_35.scala 3595:47]
      pop_20_1 <= 1'h0; // @[lut_35.scala 3595:47]
    end else begin
      pop_20_1 <= _GEN_20392;
    end
    if (reset) begin // @[lut_35.scala 3596:47]
      pop_21_1 <= 1'h0; // @[lut_35.scala 3596:47]
    end else begin
      pop_21_1 <= _GEN_20393;
    end
    if (reset) begin // @[lut_35.scala 3597:47]
      pop_22_1 <= 1'h0; // @[lut_35.scala 3597:47]
    end else begin
      pop_22_1 <= _GEN_20394;
    end
    if (reset) begin // @[lut_35.scala 3598:47]
      pop_23_1 <= 1'h0; // @[lut_35.scala 3598:47]
    end else begin
      pop_23_1 <= _GEN_20395;
    end
    if (reset) begin // @[lut_35.scala 3599:47]
      pop_24_1 <= 1'h0; // @[lut_35.scala 3599:47]
    end else begin
      pop_24_1 <= _GEN_20396;
    end
    if (reset) begin // @[lut_35.scala 3600:47]
      pop_25_1 <= 1'h0; // @[lut_35.scala 3600:47]
    end else begin
      pop_25_1 <= _GEN_20397;
    end
    if (reset) begin // @[lut_35.scala 3601:47]
      pop_26_1 <= 1'h0; // @[lut_35.scala 3601:47]
    end else begin
      pop_26_1 <= _GEN_20398;
    end
    if (reset) begin // @[lut_35.scala 3602:47]
      pop_27_1 <= 1'h0; // @[lut_35.scala 3602:47]
    end else begin
      pop_27_1 <= _GEN_20399;
    end
    if (reset) begin // @[lut_35.scala 3603:47]
      pop_28_1 <= 1'h0; // @[lut_35.scala 3603:47]
    end else begin
      pop_28_1 <= _GEN_20400;
    end
    if (reset) begin // @[lut_35.scala 3604:47]
      pop_29_1 <= 1'h0; // @[lut_35.scala 3604:47]
    end else begin
      pop_29_1 <= _GEN_20401;
    end
    if (reset) begin // @[lut_35.scala 3605:47]
      pop_30_1 <= 1'h0; // @[lut_35.scala 3605:47]
    end else begin
      pop_30_1 <= _GEN_20402;
    end
    if (reset) begin // @[lut_35.scala 3606:47]
      pop_31_1 <= 1'h0; // @[lut_35.scala 3606:47]
    end else begin
      pop_31_1 <= _GEN_20403;
    end
    if (reset) begin // @[lut_35.scala 3607:47]
      pop_32_1 <= 1'h0; // @[lut_35.scala 3607:47]
    end else begin
      pop_32_1 <= _GEN_20404;
    end
    if (reset) begin // @[lut_35.scala 3608:47]
      pop_33_1 <= 1'h0; // @[lut_35.scala 3608:47]
    end else begin
      pop_33_1 <= _GEN_20405;
    end
    if (reset) begin // @[lut_35.scala 3609:47]
      pop_34_1 <= 1'h0; // @[lut_35.scala 3609:47]
    end else begin
      pop_34_1 <= _GEN_20406;
    end
    if (reset) begin // @[lut_35.scala 3611:47]
      pop_valid_2 <= 1'h0; // @[lut_35.scala 3611:47]
    end else begin
      pop_valid_2 <= _GEN_20407;
    end
    if (reset) begin // @[lut_35.scala 3613:47]
      pop_ray_id_2 <= 32'h0; // @[lut_35.scala 3613:47]
    end else if (pop_1 & pop_valid) begin // @[lut_35.scala 3687:46]
      if (read_stack0_pop == pop_ray_id & pop_valid) begin // @[lut_35.scala 3688:67]
        pop_ray_id_2 <= pop_ray_id; // @[lut_35.scala 3726:34]
      end else if (read_stack1_pop == pop_ray_id & pop_valid) begin // @[lut_35.scala 3728:77]
        pop_ray_id_2 <= pop_ray_id; // @[lut_35.scala 3766:38]
      end else begin
        pop_ray_id_2 <= _GEN_20292;
      end
    end
    if (reset) begin // @[lut_35.scala 3614:47]
      pop_hitT_2 <= 32'h0; // @[lut_35.scala 3614:47]
    end else if (pop_1 & pop_valid) begin // @[lut_35.scala 3687:46]
      if (read_stack0_pop == pop_ray_id & pop_valid) begin // @[lut_35.scala 3688:67]
        pop_hitT_2 <= pop_hitT_1; // @[lut_35.scala 3727:37]
      end else if (read_stack1_pop == pop_ray_id & pop_valid) begin // @[lut_35.scala 3728:77]
        pop_hitT_2 <= pop_hitT_1; // @[lut_35.scala 3767:41]
      end else begin
        pop_hitT_2 <= _GEN_20293;
      end
    end
    if (reset) begin // @[lut_35.scala 3616:47]
      no_match <= 1'h0; // @[lut_35.scala 3616:47]
    end else begin
      no_match <= _T_745;
    end
    if (reset) begin // @[lut_35.scala 3682:51]
      no_match_1 <= 1'h0; // @[lut_35.scala 3682:51]
    end else begin
      no_match_1 <= no_match; // @[lut_35.scala 3684:41]
    end
    if (reset) begin // @[lut_35.scala 3683:51]
      no_match_2 <= 1'h0; // @[lut_35.scala 3683:51]
    end else begin
      no_match_2 <= no_match_1; // @[lut_35.scala 3685:41]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {2{`RANDOM}};
  _RAND_2 = {2{`RANDOM}};
  _RAND_3 = {2{`RANDOM}};
  _RAND_4 = {2{`RANDOM}};
  _RAND_5 = {2{`RANDOM}};
  _RAND_6 = {2{`RANDOM}};
  _RAND_7 = {2{`RANDOM}};
  _RAND_8 = {2{`RANDOM}};
  _RAND_9 = {2{`RANDOM}};
  _RAND_10 = {2{`RANDOM}};
  _RAND_11 = {2{`RANDOM}};
  _RAND_12 = {2{`RANDOM}};
  _RAND_13 = {2{`RANDOM}};
  _RAND_14 = {2{`RANDOM}};
  _RAND_15 = {2{`RANDOM}};
  _RAND_16 = {2{`RANDOM}};
  _RAND_17 = {2{`RANDOM}};
  _RAND_18 = {2{`RANDOM}};
  _RAND_19 = {2{`RANDOM}};
  _RAND_20 = {2{`RANDOM}};
  _RAND_21 = {2{`RANDOM}};
  _RAND_22 = {2{`RANDOM}};
  _RAND_23 = {2{`RANDOM}};
  _RAND_24 = {2{`RANDOM}};
  _RAND_25 = {2{`RANDOM}};
  _RAND_26 = {2{`RANDOM}};
  _RAND_27 = {2{`RANDOM}};
  _RAND_28 = {2{`RANDOM}};
  _RAND_29 = {2{`RANDOM}};
  _RAND_30 = {2{`RANDOM}};
  _RAND_31 = {2{`RANDOM}};
  _RAND_32 = {2{`RANDOM}};
  _RAND_33 = {2{`RANDOM}};
  _RAND_34 = {2{`RANDOM}};
  _RAND_35 = {2{`RANDOM}};
  _RAND_36 = {2{`RANDOM}};
  _RAND_37 = {2{`RANDOM}};
  _RAND_38 = {2{`RANDOM}};
  _RAND_39 = {2{`RANDOM}};
  _RAND_40 = {2{`RANDOM}};
  _RAND_41 = {2{`RANDOM}};
  _RAND_42 = {2{`RANDOM}};
  _RAND_43 = {2{`RANDOM}};
  _RAND_44 = {2{`RANDOM}};
  _RAND_45 = {2{`RANDOM}};
  _RAND_46 = {2{`RANDOM}};
  _RAND_47 = {2{`RANDOM}};
  _RAND_48 = {2{`RANDOM}};
  _RAND_49 = {2{`RANDOM}};
  _RAND_50 = {2{`RANDOM}};
  _RAND_51 = {2{`RANDOM}};
  _RAND_52 = {2{`RANDOM}};
  _RAND_53 = {2{`RANDOM}};
  _RAND_54 = {2{`RANDOM}};
  _RAND_55 = {2{`RANDOM}};
  _RAND_56 = {2{`RANDOM}};
  _RAND_57 = {2{`RANDOM}};
  _RAND_58 = {2{`RANDOM}};
  _RAND_59 = {2{`RANDOM}};
  _RAND_60 = {2{`RANDOM}};
  _RAND_61 = {2{`RANDOM}};
  _RAND_62 = {2{`RANDOM}};
  _RAND_63 = {2{`RANDOM}};
  _RAND_64 = {2{`RANDOM}};
  _RAND_65 = {2{`RANDOM}};
  _RAND_66 = {2{`RANDOM}};
  _RAND_67 = {2{`RANDOM}};
  _RAND_68 = {2{`RANDOM}};
  _RAND_69 = {2{`RANDOM}};
  _RAND_70 = {2{`RANDOM}};
  _RAND_71 = {2{`RANDOM}};
  _RAND_72 = {2{`RANDOM}};
  _RAND_73 = {2{`RANDOM}};
  _RAND_74 = {2{`RANDOM}};
  _RAND_75 = {2{`RANDOM}};
  _RAND_76 = {2{`RANDOM}};
  _RAND_77 = {2{`RANDOM}};
  _RAND_78 = {2{`RANDOM}};
  _RAND_79 = {2{`RANDOM}};
  _RAND_80 = {2{`RANDOM}};
  _RAND_81 = {2{`RANDOM}};
  _RAND_82 = {2{`RANDOM}};
  _RAND_83 = {2{`RANDOM}};
  _RAND_84 = {2{`RANDOM}};
  _RAND_85 = {2{`RANDOM}};
  _RAND_86 = {2{`RANDOM}};
  _RAND_87 = {2{`RANDOM}};
  _RAND_88 = {2{`RANDOM}};
  _RAND_89 = {2{`RANDOM}};
  _RAND_90 = {2{`RANDOM}};
  _RAND_91 = {2{`RANDOM}};
  _RAND_92 = {2{`RANDOM}};
  _RAND_93 = {2{`RANDOM}};
  _RAND_94 = {2{`RANDOM}};
  _RAND_95 = {2{`RANDOM}};
  _RAND_96 = {2{`RANDOM}};
  _RAND_97 = {2{`RANDOM}};
  _RAND_98 = {2{`RANDOM}};
  _RAND_99 = {2{`RANDOM}};
  _RAND_100 = {2{`RANDOM}};
  _RAND_101 = {2{`RANDOM}};
  _RAND_102 = {2{`RANDOM}};
  _RAND_103 = {2{`RANDOM}};
  _RAND_104 = {2{`RANDOM}};
  _RAND_105 = {2{`RANDOM}};
  _RAND_106 = {2{`RANDOM}};
  _RAND_107 = {2{`RANDOM}};
  _RAND_108 = {2{`RANDOM}};
  _RAND_109 = {2{`RANDOM}};
  _RAND_110 = {2{`RANDOM}};
  _RAND_111 = {2{`RANDOM}};
  _RAND_112 = {2{`RANDOM}};
  _RAND_113 = {2{`RANDOM}};
  _RAND_114 = {2{`RANDOM}};
  _RAND_115 = {2{`RANDOM}};
  _RAND_116 = {2{`RANDOM}};
  _RAND_117 = {2{`RANDOM}};
  _RAND_118 = {2{`RANDOM}};
  _RAND_119 = {2{`RANDOM}};
  _RAND_120 = {2{`RANDOM}};
  _RAND_121 = {2{`RANDOM}};
  _RAND_122 = {2{`RANDOM}};
  _RAND_123 = {2{`RANDOM}};
  _RAND_124 = {2{`RANDOM}};
  _RAND_125 = {2{`RANDOM}};
  _RAND_126 = {2{`RANDOM}};
  _RAND_127 = {2{`RANDOM}};
  _RAND_128 = {2{`RANDOM}};
  _RAND_129 = {2{`RANDOM}};
  _RAND_130 = {2{`RANDOM}};
  _RAND_131 = {2{`RANDOM}};
  _RAND_132 = {2{`RANDOM}};
  _RAND_133 = {2{`RANDOM}};
  _RAND_134 = {2{`RANDOM}};
  _RAND_135 = {2{`RANDOM}};
  _RAND_136 = {2{`RANDOM}};
  _RAND_137 = {2{`RANDOM}};
  _RAND_138 = {2{`RANDOM}};
  _RAND_139 = {2{`RANDOM}};
  _RAND_140 = {2{`RANDOM}};
  _RAND_141 = {2{`RANDOM}};
  _RAND_142 = {2{`RANDOM}};
  _RAND_143 = {2{`RANDOM}};
  _RAND_144 = {2{`RANDOM}};
  _RAND_145 = {2{`RANDOM}};
  _RAND_146 = {2{`RANDOM}};
  _RAND_147 = {2{`RANDOM}};
  _RAND_148 = {2{`RANDOM}};
  _RAND_149 = {2{`RANDOM}};
  _RAND_150 = {2{`RANDOM}};
  _RAND_151 = {2{`RANDOM}};
  _RAND_152 = {2{`RANDOM}};
  _RAND_153 = {2{`RANDOM}};
  _RAND_154 = {2{`RANDOM}};
  _RAND_155 = {2{`RANDOM}};
  _RAND_156 = {2{`RANDOM}};
  _RAND_157 = {2{`RANDOM}};
  _RAND_158 = {2{`RANDOM}};
  _RAND_159 = {2{`RANDOM}};
  _RAND_160 = {2{`RANDOM}};
  _RAND_161 = {2{`RANDOM}};
  _RAND_162 = {2{`RANDOM}};
  _RAND_163 = {2{`RANDOM}};
  _RAND_164 = {2{`RANDOM}};
  _RAND_165 = {2{`RANDOM}};
  _RAND_166 = {2{`RANDOM}};
  _RAND_167 = {2{`RANDOM}};
  _RAND_168 = {2{`RANDOM}};
  _RAND_169 = {2{`RANDOM}};
  _RAND_170 = {2{`RANDOM}};
  _RAND_171 = {2{`RANDOM}};
  _RAND_172 = {2{`RANDOM}};
  _RAND_173 = {2{`RANDOM}};
  _RAND_174 = {2{`RANDOM}};
  _RAND_175 = {2{`RANDOM}};
  _RAND_176 = {2{`RANDOM}};
  _RAND_177 = {2{`RANDOM}};
  _RAND_178 = {2{`RANDOM}};
  _RAND_179 = {2{`RANDOM}};
  _RAND_180 = {2{`RANDOM}};
  _RAND_181 = {2{`RANDOM}};
  _RAND_182 = {2{`RANDOM}};
  _RAND_183 = {2{`RANDOM}};
  _RAND_184 = {2{`RANDOM}};
  _RAND_185 = {2{`RANDOM}};
  _RAND_186 = {2{`RANDOM}};
  _RAND_187 = {2{`RANDOM}};
  _RAND_188 = {2{`RANDOM}};
  _RAND_189 = {2{`RANDOM}};
  _RAND_190 = {2{`RANDOM}};
  _RAND_191 = {2{`RANDOM}};
  _RAND_192 = {2{`RANDOM}};
  _RAND_193 = {2{`RANDOM}};
  _RAND_194 = {2{`RANDOM}};
  _RAND_195 = {2{`RANDOM}};
  _RAND_196 = {2{`RANDOM}};
  _RAND_197 = {2{`RANDOM}};
  _RAND_198 = {2{`RANDOM}};
  _RAND_199 = {2{`RANDOM}};
  _RAND_200 = {2{`RANDOM}};
  _RAND_201 = {2{`RANDOM}};
  _RAND_202 = {2{`RANDOM}};
  _RAND_203 = {2{`RANDOM}};
  _RAND_204 = {2{`RANDOM}};
  _RAND_205 = {2{`RANDOM}};
  _RAND_206 = {2{`RANDOM}};
  _RAND_207 = {2{`RANDOM}};
  _RAND_208 = {2{`RANDOM}};
  _RAND_209 = {2{`RANDOM}};
  _RAND_210 = {2{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 35; initvar = initvar+1)
    LUT_mem[initvar] = _RAND_0[32:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  read_stack0 = _RAND_211[31:0];
  _RAND_212 = {1{`RANDOM}};
  read_stack1 = _RAND_212[31:0];
  _RAND_213 = {1{`RANDOM}};
  read_stack2 = _RAND_213[31:0];
  _RAND_214 = {1{`RANDOM}};
  read_stack3 = _RAND_214[31:0];
  _RAND_215 = {1{`RANDOM}};
  read_stack4 = _RAND_215[31:0];
  _RAND_216 = {1{`RANDOM}};
  read_stack5 = _RAND_216[31:0];
  _RAND_217 = {1{`RANDOM}};
  read_stack6 = _RAND_217[31:0];
  _RAND_218 = {1{`RANDOM}};
  read_stack7 = _RAND_218[31:0];
  _RAND_219 = {1{`RANDOM}};
  read_stack8 = _RAND_219[31:0];
  _RAND_220 = {1{`RANDOM}};
  read_stack9 = _RAND_220[31:0];
  _RAND_221 = {1{`RANDOM}};
  read_stack10 = _RAND_221[31:0];
  _RAND_222 = {1{`RANDOM}};
  read_stack11 = _RAND_222[31:0];
  _RAND_223 = {1{`RANDOM}};
  read_stack12 = _RAND_223[31:0];
  _RAND_224 = {1{`RANDOM}};
  read_stack13 = _RAND_224[31:0];
  _RAND_225 = {1{`RANDOM}};
  read_stack14 = _RAND_225[31:0];
  _RAND_226 = {1{`RANDOM}};
  read_stack15 = _RAND_226[31:0];
  _RAND_227 = {1{`RANDOM}};
  read_stack16 = _RAND_227[31:0];
  _RAND_228 = {1{`RANDOM}};
  read_stack17 = _RAND_228[31:0];
  _RAND_229 = {1{`RANDOM}};
  read_stack18 = _RAND_229[31:0];
  _RAND_230 = {1{`RANDOM}};
  read_stack19 = _RAND_230[31:0];
  _RAND_231 = {1{`RANDOM}};
  read_stack20 = _RAND_231[31:0];
  _RAND_232 = {1{`RANDOM}};
  read_stack21 = _RAND_232[31:0];
  _RAND_233 = {1{`RANDOM}};
  read_stack22 = _RAND_233[31:0];
  _RAND_234 = {1{`RANDOM}};
  read_stack23 = _RAND_234[31:0];
  _RAND_235 = {1{`RANDOM}};
  read_stack24 = _RAND_235[31:0];
  _RAND_236 = {1{`RANDOM}};
  read_stack25 = _RAND_236[31:0];
  _RAND_237 = {1{`RANDOM}};
  read_stack26 = _RAND_237[31:0];
  _RAND_238 = {1{`RANDOM}};
  read_stack27 = _RAND_238[31:0];
  _RAND_239 = {1{`RANDOM}};
  read_stack28 = _RAND_239[31:0];
  _RAND_240 = {1{`RANDOM}};
  read_stack29 = _RAND_240[31:0];
  _RAND_241 = {1{`RANDOM}};
  read_stack30 = _RAND_241[31:0];
  _RAND_242 = {1{`RANDOM}};
  read_stack31 = _RAND_242[31:0];
  _RAND_243 = {1{`RANDOM}};
  read_stack32 = _RAND_243[31:0];
  _RAND_244 = {1{`RANDOM}};
  read_stack33 = _RAND_244[31:0];
  _RAND_245 = {1{`RANDOM}};
  read_stack34 = _RAND_245[31:0];
  _RAND_246 = {1{`RANDOM}};
  push_0_1 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  push_1_1 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  push_2_1 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  push_3_1 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  push_4_1 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  push_5_1 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  push_6_1 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  push_7_1 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  push_8_1 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  push_9_1 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  push_10_1 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  push_11_1 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  push_12_1 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  push_13_1 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  push_14_1 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  push_15_1 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  push_16_1 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  push_17_1 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  push_18_1 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  push_19_1 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  push_20_1 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  push_21_1 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  push_22_1 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  push_23_1 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  push_24_1 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  push_25_1 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  push_26_1 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  push_27_1 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  push_28_1 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  push_29_1 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  push_30_1 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  push_31_1 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  push_32_1 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  push_33_1 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  push_34_1 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  push_1 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  push_valid = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  push_ray_id = _RAND_283[31:0];
  _RAND_284 = {1{`RANDOM}};
  push_valid_2 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  pop_1 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  read_stack0_pop = _RAND_286[31:0];
  _RAND_287 = {1{`RANDOM}};
  read_stack1_pop = _RAND_287[31:0];
  _RAND_288 = {1{`RANDOM}};
  read_stack2_pop = _RAND_288[31:0];
  _RAND_289 = {1{`RANDOM}};
  read_stack3_pop = _RAND_289[31:0];
  _RAND_290 = {1{`RANDOM}};
  read_stack4_pop = _RAND_290[31:0];
  _RAND_291 = {1{`RANDOM}};
  read_stack5_pop = _RAND_291[31:0];
  _RAND_292 = {1{`RANDOM}};
  read_stack6_pop = _RAND_292[31:0];
  _RAND_293 = {1{`RANDOM}};
  read_stack7_pop = _RAND_293[31:0];
  _RAND_294 = {1{`RANDOM}};
  read_stack8_pop = _RAND_294[31:0];
  _RAND_295 = {1{`RANDOM}};
  read_stack9_pop = _RAND_295[31:0];
  _RAND_296 = {1{`RANDOM}};
  read_stack10_pop = _RAND_296[31:0];
  _RAND_297 = {1{`RANDOM}};
  read_stack11_pop = _RAND_297[31:0];
  _RAND_298 = {1{`RANDOM}};
  read_stack12_pop = _RAND_298[31:0];
  _RAND_299 = {1{`RANDOM}};
  read_stack13_pop = _RAND_299[31:0];
  _RAND_300 = {1{`RANDOM}};
  read_stack14_pop = _RAND_300[31:0];
  _RAND_301 = {1{`RANDOM}};
  read_stack15_pop = _RAND_301[31:0];
  _RAND_302 = {1{`RANDOM}};
  read_stack16_pop = _RAND_302[31:0];
  _RAND_303 = {1{`RANDOM}};
  read_stack17_pop = _RAND_303[31:0];
  _RAND_304 = {1{`RANDOM}};
  read_stack18_pop = _RAND_304[31:0];
  _RAND_305 = {1{`RANDOM}};
  read_stack19_pop = _RAND_305[31:0];
  _RAND_306 = {1{`RANDOM}};
  read_stack20_pop = _RAND_306[31:0];
  _RAND_307 = {1{`RANDOM}};
  read_stack21_pop = _RAND_307[31:0];
  _RAND_308 = {1{`RANDOM}};
  read_stack22_pop = _RAND_308[31:0];
  _RAND_309 = {1{`RANDOM}};
  read_stack23_pop = _RAND_309[31:0];
  _RAND_310 = {1{`RANDOM}};
  read_stack24_pop = _RAND_310[31:0];
  _RAND_311 = {1{`RANDOM}};
  read_stack25_pop = _RAND_311[31:0];
  _RAND_312 = {1{`RANDOM}};
  read_stack26_pop = _RAND_312[31:0];
  _RAND_313 = {1{`RANDOM}};
  read_stack27_pop = _RAND_313[31:0];
  _RAND_314 = {1{`RANDOM}};
  read_stack28_pop = _RAND_314[31:0];
  _RAND_315 = {1{`RANDOM}};
  read_stack29_pop = _RAND_315[31:0];
  _RAND_316 = {1{`RANDOM}};
  read_stack30_pop = _RAND_316[31:0];
  _RAND_317 = {1{`RANDOM}};
  read_stack31_pop = _RAND_317[31:0];
  _RAND_318 = {1{`RANDOM}};
  read_stack32_pop = _RAND_318[31:0];
  _RAND_319 = {1{`RANDOM}};
  read_stack33_pop = _RAND_319[31:0];
  _RAND_320 = {1{`RANDOM}};
  read_stack34_pop = _RAND_320[31:0];
  _RAND_321 = {1{`RANDOM}};
  pop_ray_id = _RAND_321[31:0];
  _RAND_322 = {1{`RANDOM}};
  pop_hitT_1 = _RAND_322[31:0];
  _RAND_323 = {1{`RANDOM}};
  pop_valid = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  pop_0_1 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  pop_1_1 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  pop_2_1 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  pop_3_1 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  pop_4_1 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  pop_5_1 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  pop_6_1 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  pop_7_1 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  pop_8_1 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  pop_9_1 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  pop_10_1 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  pop_11_1 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  pop_12_1 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  pop_13_1 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  pop_14_1 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  pop_15_1 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  pop_16_1 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  pop_17_1 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  pop_18_1 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  pop_19_1 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  pop_20_1 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  pop_21_1 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  pop_22_1 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  pop_23_1 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  pop_24_1 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  pop_25_1 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  pop_26_1 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  pop_27_1 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  pop_28_1 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  pop_29_1 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  pop_30_1 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  pop_31_1 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  pop_32_1 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  pop_33_1 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  pop_34_1 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  pop_valid_2 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  pop_ray_id_2 = _RAND_360[31:0];
  _RAND_361 = {1{`RANDOM}};
  pop_hitT_2 = _RAND_361[31:0];
  _RAND_362 = {1{`RANDOM}};
  no_match = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  no_match_1 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  no_match_2 = _RAND_364[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Stack(
  input         clock,
  input         reset,
  input         io_push,
  input         io_pop,
  input  [31:0] io_dataIn,
  input  [31:0] io_ray_id,
  output [31:0] io_dataOut,
  output        io_empty,
  input  [31:0] io_hit_in,
  output [31:0] io_hit_out,
  output [31:0] io_ray_out,
  output        io_enable
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] stack_mem [0:31]; // @[stack.scala 26:24]
  wire [31:0] stack_mem_MPORT_1_data; // @[stack.scala 26:24]
  wire [4:0] stack_mem_MPORT_1_addr; // @[stack.scala 26:24]
  wire [31:0] stack_mem_MPORT_data; // @[stack.scala 26:24]
  wire [4:0] stack_mem_MPORT_addr; // @[stack.scala 26:24]
  wire  stack_mem_MPORT_mask; // @[stack.scala 26:24]
  wire  stack_mem_MPORT_en; // @[stack.scala 26:24]
  reg [5:0] sp; // @[stack.scala 27:21]
  reg [31:0] out; // @[stack.scala 28:22]
  reg [31:0] hit_1; // @[stack.scala 29:23]
  reg [31:0] ray_1; // @[stack.scala 30:23]
  reg  enable; // @[stack.scala 31:25]
  wire  _T = sp < 6'h20; // @[stack.scala 37:25]
  wire  _T_1 = io_push & sp < 6'h20; // @[stack.scala 37:18]
  wire [5:0] _T_4 = sp + 6'h1; // @[stack.scala 39:18]
  wire  _T_6 = io_pop & sp >= 6'h1; // @[stack.scala 42:24]
  wire [5:0] _T_8 = sp - 6'h1; // @[stack.scala 43:28]
  assign stack_mem_MPORT_1_addr = _T_8[4:0];
  assign stack_mem_MPORT_1_data = stack_mem[stack_mem_MPORT_1_addr]; // @[stack.scala 26:24]
  assign stack_mem_MPORT_data = io_dataIn;
  assign stack_mem_MPORT_addr = sp[4:0];
  assign stack_mem_MPORT_mask = 1'h1;
  assign stack_mem_MPORT_en = io_push & _T;
  assign io_dataOut = out; // @[stack.scala 61:16]
  assign io_empty = sp == 6'h0; // @[stack.scala 60:21]
  assign io_hit_out = hit_1; // @[stack.scala 62:18]
  assign io_ray_out = ray_1; // @[stack.scala 63:21]
  assign io_enable = enable; // @[stack.scala 64:18]
  always @(posedge clock) begin
    if(stack_mem_MPORT_en & stack_mem_MPORT_mask) begin
      stack_mem[stack_mem_MPORT_addr] <= stack_mem_MPORT_data; // @[stack.scala 26:24]
    end
    if (reset) begin // @[stack.scala 27:21]
      sp <= 6'h0; // @[stack.scala 27:21]
    end else if (io_push & sp < 6'h20) begin // @[stack.scala 37:42]
      sp <= _T_4; // @[stack.scala 39:12]
    end else if (io_pop & sp >= 6'h1) begin // @[stack.scala 42:39]
      sp <= _T_8; // @[stack.scala 44:12]
    end
    if (reset) begin // @[stack.scala 28:22]
      out <= 32'sh0; // @[stack.scala 28:22]
    end else if (!(io_push & sp < 6'h20)) begin // @[stack.scala 37:42]
      if (io_pop & sp >= 6'h1) begin // @[stack.scala 42:39]
        out <= stack_mem_MPORT_1_data; // @[stack.scala 43:13]
      end
    end
    if (reset) begin // @[stack.scala 29:23]
      hit_1 <= 32'h0; // @[stack.scala 29:23]
    end else if (!(io_push & sp < 6'h20)) begin // @[stack.scala 37:42]
      if (io_pop & sp >= 6'h1) begin // @[stack.scala 42:39]
        hit_1 <= io_hit_in; // @[stack.scala 45:15]
      end else begin
        hit_1 <= 32'h0; // @[stack.scala 49:16]
      end
    end
    if (reset) begin // @[stack.scala 30:23]
      ray_1 <= 32'h0; // @[stack.scala 30:23]
    end else if (!(io_push & sp < 6'h20)) begin // @[stack.scala 37:42]
      if (io_pop & sp >= 6'h1) begin // @[stack.scala 42:39]
        ray_1 <= io_ray_id; // @[stack.scala 46:15]
      end else begin
        ray_1 <= 32'h0; // @[stack.scala 50:15]
      end
    end
    if (reset) begin // @[stack.scala 31:25]
      enable <= 1'h0; // @[stack.scala 31:25]
    end else if (io_push & sp < 6'h20) begin // @[stack.scala 37:42]
      enable <= 1'h0; // @[stack.scala 40:15]
    end else begin
      enable <= _T_6;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    stack_mem[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  sp = _RAND_1[5:0];
  _RAND_2 = {1{`RANDOM}};
  out = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  hit_1 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  ray_1 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  enable = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Stackmanage(
  input         clock,
  input         reset,
  input         io_push,
  input         io_push_en,
  input         io_pop,
  input         io_pop_en,
  input  [31:0] io_ray_id_push,
  input  [31:0] io_ray_id_pop,
  input  [31:0] io_node_id_push_in,
  input  [31:0] io_hitT_in,
  output [31:0] io_hitT_out,
  output [31:0] io_node_id_out,
  output [31:0] io_ray_id_out,
  output        io_pop_valid,
  output        io_Dis_en,
  output        io_Finish
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
`endif // RANDOMIZE_REG_INIT
  wire  LUT_stack_clock; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_reset; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_push; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_push_valid; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_pop; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_pop_valid; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_empty_0; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_empty_1; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_empty_2; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_empty_3; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_empty_4; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_empty_5; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_empty_6; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_empty_7; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_empty_8; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_empty_9; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_empty_10; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_empty_11; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_empty_12; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_empty_13; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_empty_14; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_empty_15; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_empty_16; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_empty_17; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_empty_18; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_empty_19; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_empty_20; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_empty_21; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_empty_22; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_empty_23; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_empty_24; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_empty_25; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_empty_26; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_empty_27; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_empty_28; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_empty_29; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_empty_30; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_empty_31; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_empty_32; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_empty_33; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_empty_34; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_dispatch_0; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_dispatch_1; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_dispatch_2; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_dispatch_3; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_dispatch_4; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_dispatch_5; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_dispatch_6; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_dispatch_7; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_dispatch_8; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_dispatch_9; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_dispatch_10; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_dispatch_11; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_dispatch_12; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_dispatch_13; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_dispatch_14; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_dispatch_15; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_dispatch_16; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_dispatch_17; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_dispatch_18; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_dispatch_19; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_dispatch_20; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_dispatch_21; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_dispatch_22; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_dispatch_23; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_dispatch_24; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_dispatch_25; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_dispatch_26; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_dispatch_27; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_dispatch_28; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_dispatch_29; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_dispatch_30; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_dispatch_31; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_dispatch_32; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_dispatch_33; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_dispatch_34; // @[stackmanage_35.scala 33:45]
  wire [31:0] LUT_stack_io_ray_id_push; // @[stackmanage_35.scala 33:45]
  wire [31:0] LUT_stack_io_ray_id_pop; // @[stackmanage_35.scala 33:45]
  wire [31:0] LUT_stack_io_node_id_push_in; // @[stackmanage_35.scala 33:45]
  wire [31:0] LUT_stack_io_hitT_in; // @[stackmanage_35.scala 33:45]
  wire [31:0] LUT_stack_io_ray_id_pop_out; // @[stackmanage_35.scala 33:45]
  wire [31:0] LUT_stack_io_hitT_out; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_pop_0; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_pop_1; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_pop_2; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_pop_3; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_pop_4; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_pop_5; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_pop_6; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_pop_7; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_pop_8; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_pop_9; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_pop_10; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_pop_11; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_pop_12; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_pop_13; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_pop_14; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_pop_15; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_pop_16; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_pop_17; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_pop_18; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_pop_19; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_pop_20; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_pop_21; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_pop_22; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_pop_23; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_pop_24; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_pop_25; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_pop_26; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_pop_27; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_pop_28; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_pop_29; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_pop_30; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_pop_31; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_pop_32; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_pop_33; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_pop_34; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_pop_en; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_push_0; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_push_1; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_push_2; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_push_3; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_push_4; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_push_5; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_push_6; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_push_7; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_push_8; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_push_9; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_push_10; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_push_11; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_push_12; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_push_13; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_push_14; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_push_15; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_push_16; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_push_17; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_push_18; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_push_19; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_push_20; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_push_21; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_push_22; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_push_23; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_push_24; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_push_25; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_push_26; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_push_27; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_push_28; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_push_29; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_push_30; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_push_31; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_push_32; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_push_33; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_push_34; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_push_en; // @[stackmanage_35.scala 33:45]
  wire  LUT_stack_io_no_match; // @[stackmanage_35.scala 33:45]
  wire  Stack_0_clock; // @[stackmanage_35.scala 34:48]
  wire  Stack_0_reset; // @[stackmanage_35.scala 34:48]
  wire  Stack_0_io_push; // @[stackmanage_35.scala 34:48]
  wire  Stack_0_io_pop; // @[stackmanage_35.scala 34:48]
  wire [31:0] Stack_0_io_dataIn; // @[stackmanage_35.scala 34:48]
  wire [31:0] Stack_0_io_ray_id; // @[stackmanage_35.scala 34:48]
  wire [31:0] Stack_0_io_dataOut; // @[stackmanage_35.scala 34:48]
  wire  Stack_0_io_empty; // @[stackmanage_35.scala 34:48]
  wire [31:0] Stack_0_io_hit_in; // @[stackmanage_35.scala 34:48]
  wire [31:0] Stack_0_io_hit_out; // @[stackmanage_35.scala 34:48]
  wire [31:0] Stack_0_io_ray_out; // @[stackmanage_35.scala 34:48]
  wire  Stack_0_io_enable; // @[stackmanage_35.scala 34:48]
  wire  Stack_1_clock; // @[stackmanage_35.scala 35:48]
  wire  Stack_1_reset; // @[stackmanage_35.scala 35:48]
  wire  Stack_1_io_push; // @[stackmanage_35.scala 35:48]
  wire  Stack_1_io_pop; // @[stackmanage_35.scala 35:48]
  wire [31:0] Stack_1_io_dataIn; // @[stackmanage_35.scala 35:48]
  wire [31:0] Stack_1_io_ray_id; // @[stackmanage_35.scala 35:48]
  wire [31:0] Stack_1_io_dataOut; // @[stackmanage_35.scala 35:48]
  wire  Stack_1_io_empty; // @[stackmanage_35.scala 35:48]
  wire [31:0] Stack_1_io_hit_in; // @[stackmanage_35.scala 35:48]
  wire [31:0] Stack_1_io_hit_out; // @[stackmanage_35.scala 35:48]
  wire [31:0] Stack_1_io_ray_out; // @[stackmanage_35.scala 35:48]
  wire  Stack_1_io_enable; // @[stackmanage_35.scala 35:48]
  wire  Stack_2_clock; // @[stackmanage_35.scala 36:48]
  wire  Stack_2_reset; // @[stackmanage_35.scala 36:48]
  wire  Stack_2_io_push; // @[stackmanage_35.scala 36:48]
  wire  Stack_2_io_pop; // @[stackmanage_35.scala 36:48]
  wire [31:0] Stack_2_io_dataIn; // @[stackmanage_35.scala 36:48]
  wire [31:0] Stack_2_io_ray_id; // @[stackmanage_35.scala 36:48]
  wire [31:0] Stack_2_io_dataOut; // @[stackmanage_35.scala 36:48]
  wire  Stack_2_io_empty; // @[stackmanage_35.scala 36:48]
  wire [31:0] Stack_2_io_hit_in; // @[stackmanage_35.scala 36:48]
  wire [31:0] Stack_2_io_hit_out; // @[stackmanage_35.scala 36:48]
  wire [31:0] Stack_2_io_ray_out; // @[stackmanage_35.scala 36:48]
  wire  Stack_2_io_enable; // @[stackmanage_35.scala 36:48]
  wire  Stack_3_clock; // @[stackmanage_35.scala 37:48]
  wire  Stack_3_reset; // @[stackmanage_35.scala 37:48]
  wire  Stack_3_io_push; // @[stackmanage_35.scala 37:48]
  wire  Stack_3_io_pop; // @[stackmanage_35.scala 37:48]
  wire [31:0] Stack_3_io_dataIn; // @[stackmanage_35.scala 37:48]
  wire [31:0] Stack_3_io_ray_id; // @[stackmanage_35.scala 37:48]
  wire [31:0] Stack_3_io_dataOut; // @[stackmanage_35.scala 37:48]
  wire  Stack_3_io_empty; // @[stackmanage_35.scala 37:48]
  wire [31:0] Stack_3_io_hit_in; // @[stackmanage_35.scala 37:48]
  wire [31:0] Stack_3_io_hit_out; // @[stackmanage_35.scala 37:48]
  wire [31:0] Stack_3_io_ray_out; // @[stackmanage_35.scala 37:48]
  wire  Stack_3_io_enable; // @[stackmanage_35.scala 37:48]
  wire  Stack_4_clock; // @[stackmanage_35.scala 38:48]
  wire  Stack_4_reset; // @[stackmanage_35.scala 38:48]
  wire  Stack_4_io_push; // @[stackmanage_35.scala 38:48]
  wire  Stack_4_io_pop; // @[stackmanage_35.scala 38:48]
  wire [31:0] Stack_4_io_dataIn; // @[stackmanage_35.scala 38:48]
  wire [31:0] Stack_4_io_ray_id; // @[stackmanage_35.scala 38:48]
  wire [31:0] Stack_4_io_dataOut; // @[stackmanage_35.scala 38:48]
  wire  Stack_4_io_empty; // @[stackmanage_35.scala 38:48]
  wire [31:0] Stack_4_io_hit_in; // @[stackmanage_35.scala 38:48]
  wire [31:0] Stack_4_io_hit_out; // @[stackmanage_35.scala 38:48]
  wire [31:0] Stack_4_io_ray_out; // @[stackmanage_35.scala 38:48]
  wire  Stack_4_io_enable; // @[stackmanage_35.scala 38:48]
  wire  Stack_5_clock; // @[stackmanage_35.scala 39:48]
  wire  Stack_5_reset; // @[stackmanage_35.scala 39:48]
  wire  Stack_5_io_push; // @[stackmanage_35.scala 39:48]
  wire  Stack_5_io_pop; // @[stackmanage_35.scala 39:48]
  wire [31:0] Stack_5_io_dataIn; // @[stackmanage_35.scala 39:48]
  wire [31:0] Stack_5_io_ray_id; // @[stackmanage_35.scala 39:48]
  wire [31:0] Stack_5_io_dataOut; // @[stackmanage_35.scala 39:48]
  wire  Stack_5_io_empty; // @[stackmanage_35.scala 39:48]
  wire [31:0] Stack_5_io_hit_in; // @[stackmanage_35.scala 39:48]
  wire [31:0] Stack_5_io_hit_out; // @[stackmanage_35.scala 39:48]
  wire [31:0] Stack_5_io_ray_out; // @[stackmanage_35.scala 39:48]
  wire  Stack_5_io_enable; // @[stackmanage_35.scala 39:48]
  wire  Stack_6_clock; // @[stackmanage_35.scala 40:48]
  wire  Stack_6_reset; // @[stackmanage_35.scala 40:48]
  wire  Stack_6_io_push; // @[stackmanage_35.scala 40:48]
  wire  Stack_6_io_pop; // @[stackmanage_35.scala 40:48]
  wire [31:0] Stack_6_io_dataIn; // @[stackmanage_35.scala 40:48]
  wire [31:0] Stack_6_io_ray_id; // @[stackmanage_35.scala 40:48]
  wire [31:0] Stack_6_io_dataOut; // @[stackmanage_35.scala 40:48]
  wire  Stack_6_io_empty; // @[stackmanage_35.scala 40:48]
  wire [31:0] Stack_6_io_hit_in; // @[stackmanage_35.scala 40:48]
  wire [31:0] Stack_6_io_hit_out; // @[stackmanage_35.scala 40:48]
  wire [31:0] Stack_6_io_ray_out; // @[stackmanage_35.scala 40:48]
  wire  Stack_6_io_enable; // @[stackmanage_35.scala 40:48]
  wire  Stack_7_clock; // @[stackmanage_35.scala 41:48]
  wire  Stack_7_reset; // @[stackmanage_35.scala 41:48]
  wire  Stack_7_io_push; // @[stackmanage_35.scala 41:48]
  wire  Stack_7_io_pop; // @[stackmanage_35.scala 41:48]
  wire [31:0] Stack_7_io_dataIn; // @[stackmanage_35.scala 41:48]
  wire [31:0] Stack_7_io_ray_id; // @[stackmanage_35.scala 41:48]
  wire [31:0] Stack_7_io_dataOut; // @[stackmanage_35.scala 41:48]
  wire  Stack_7_io_empty; // @[stackmanage_35.scala 41:48]
  wire [31:0] Stack_7_io_hit_in; // @[stackmanage_35.scala 41:48]
  wire [31:0] Stack_7_io_hit_out; // @[stackmanage_35.scala 41:48]
  wire [31:0] Stack_7_io_ray_out; // @[stackmanage_35.scala 41:48]
  wire  Stack_7_io_enable; // @[stackmanage_35.scala 41:48]
  wire  Stack_8_clock; // @[stackmanage_35.scala 42:48]
  wire  Stack_8_reset; // @[stackmanage_35.scala 42:48]
  wire  Stack_8_io_push; // @[stackmanage_35.scala 42:48]
  wire  Stack_8_io_pop; // @[stackmanage_35.scala 42:48]
  wire [31:0] Stack_8_io_dataIn; // @[stackmanage_35.scala 42:48]
  wire [31:0] Stack_8_io_ray_id; // @[stackmanage_35.scala 42:48]
  wire [31:0] Stack_8_io_dataOut; // @[stackmanage_35.scala 42:48]
  wire  Stack_8_io_empty; // @[stackmanage_35.scala 42:48]
  wire [31:0] Stack_8_io_hit_in; // @[stackmanage_35.scala 42:48]
  wire [31:0] Stack_8_io_hit_out; // @[stackmanage_35.scala 42:48]
  wire [31:0] Stack_8_io_ray_out; // @[stackmanage_35.scala 42:48]
  wire  Stack_8_io_enable; // @[stackmanage_35.scala 42:48]
  wire  Stack_9_clock; // @[stackmanage_35.scala 43:48]
  wire  Stack_9_reset; // @[stackmanage_35.scala 43:48]
  wire  Stack_9_io_push; // @[stackmanage_35.scala 43:48]
  wire  Stack_9_io_pop; // @[stackmanage_35.scala 43:48]
  wire [31:0] Stack_9_io_dataIn; // @[stackmanage_35.scala 43:48]
  wire [31:0] Stack_9_io_ray_id; // @[stackmanage_35.scala 43:48]
  wire [31:0] Stack_9_io_dataOut; // @[stackmanage_35.scala 43:48]
  wire  Stack_9_io_empty; // @[stackmanage_35.scala 43:48]
  wire [31:0] Stack_9_io_hit_in; // @[stackmanage_35.scala 43:48]
  wire [31:0] Stack_9_io_hit_out; // @[stackmanage_35.scala 43:48]
  wire [31:0] Stack_9_io_ray_out; // @[stackmanage_35.scala 43:48]
  wire  Stack_9_io_enable; // @[stackmanage_35.scala 43:48]
  wire  Stack_10_clock; // @[stackmanage_35.scala 44:47]
  wire  Stack_10_reset; // @[stackmanage_35.scala 44:47]
  wire  Stack_10_io_push; // @[stackmanage_35.scala 44:47]
  wire  Stack_10_io_pop; // @[stackmanage_35.scala 44:47]
  wire [31:0] Stack_10_io_dataIn; // @[stackmanage_35.scala 44:47]
  wire [31:0] Stack_10_io_ray_id; // @[stackmanage_35.scala 44:47]
  wire [31:0] Stack_10_io_dataOut; // @[stackmanage_35.scala 44:47]
  wire  Stack_10_io_empty; // @[stackmanage_35.scala 44:47]
  wire [31:0] Stack_10_io_hit_in; // @[stackmanage_35.scala 44:47]
  wire [31:0] Stack_10_io_hit_out; // @[stackmanage_35.scala 44:47]
  wire [31:0] Stack_10_io_ray_out; // @[stackmanage_35.scala 44:47]
  wire  Stack_10_io_enable; // @[stackmanage_35.scala 44:47]
  wire  Stack_11_clock; // @[stackmanage_35.scala 45:47]
  wire  Stack_11_reset; // @[stackmanage_35.scala 45:47]
  wire  Stack_11_io_push; // @[stackmanage_35.scala 45:47]
  wire  Stack_11_io_pop; // @[stackmanage_35.scala 45:47]
  wire [31:0] Stack_11_io_dataIn; // @[stackmanage_35.scala 45:47]
  wire [31:0] Stack_11_io_ray_id; // @[stackmanage_35.scala 45:47]
  wire [31:0] Stack_11_io_dataOut; // @[stackmanage_35.scala 45:47]
  wire  Stack_11_io_empty; // @[stackmanage_35.scala 45:47]
  wire [31:0] Stack_11_io_hit_in; // @[stackmanage_35.scala 45:47]
  wire [31:0] Stack_11_io_hit_out; // @[stackmanage_35.scala 45:47]
  wire [31:0] Stack_11_io_ray_out; // @[stackmanage_35.scala 45:47]
  wire  Stack_11_io_enable; // @[stackmanage_35.scala 45:47]
  wire  Stack_12_clock; // @[stackmanage_35.scala 46:47]
  wire  Stack_12_reset; // @[stackmanage_35.scala 46:47]
  wire  Stack_12_io_push; // @[stackmanage_35.scala 46:47]
  wire  Stack_12_io_pop; // @[stackmanage_35.scala 46:47]
  wire [31:0] Stack_12_io_dataIn; // @[stackmanage_35.scala 46:47]
  wire [31:0] Stack_12_io_ray_id; // @[stackmanage_35.scala 46:47]
  wire [31:0] Stack_12_io_dataOut; // @[stackmanage_35.scala 46:47]
  wire  Stack_12_io_empty; // @[stackmanage_35.scala 46:47]
  wire [31:0] Stack_12_io_hit_in; // @[stackmanage_35.scala 46:47]
  wire [31:0] Stack_12_io_hit_out; // @[stackmanage_35.scala 46:47]
  wire [31:0] Stack_12_io_ray_out; // @[stackmanage_35.scala 46:47]
  wire  Stack_12_io_enable; // @[stackmanage_35.scala 46:47]
  wire  Stack_13_clock; // @[stackmanage_35.scala 47:47]
  wire  Stack_13_reset; // @[stackmanage_35.scala 47:47]
  wire  Stack_13_io_push; // @[stackmanage_35.scala 47:47]
  wire  Stack_13_io_pop; // @[stackmanage_35.scala 47:47]
  wire [31:0] Stack_13_io_dataIn; // @[stackmanage_35.scala 47:47]
  wire [31:0] Stack_13_io_ray_id; // @[stackmanage_35.scala 47:47]
  wire [31:0] Stack_13_io_dataOut; // @[stackmanage_35.scala 47:47]
  wire  Stack_13_io_empty; // @[stackmanage_35.scala 47:47]
  wire [31:0] Stack_13_io_hit_in; // @[stackmanage_35.scala 47:47]
  wire [31:0] Stack_13_io_hit_out; // @[stackmanage_35.scala 47:47]
  wire [31:0] Stack_13_io_ray_out; // @[stackmanage_35.scala 47:47]
  wire  Stack_13_io_enable; // @[stackmanage_35.scala 47:47]
  wire  Stack_14_clock; // @[stackmanage_35.scala 48:47]
  wire  Stack_14_reset; // @[stackmanage_35.scala 48:47]
  wire  Stack_14_io_push; // @[stackmanage_35.scala 48:47]
  wire  Stack_14_io_pop; // @[stackmanage_35.scala 48:47]
  wire [31:0] Stack_14_io_dataIn; // @[stackmanage_35.scala 48:47]
  wire [31:0] Stack_14_io_ray_id; // @[stackmanage_35.scala 48:47]
  wire [31:0] Stack_14_io_dataOut; // @[stackmanage_35.scala 48:47]
  wire  Stack_14_io_empty; // @[stackmanage_35.scala 48:47]
  wire [31:0] Stack_14_io_hit_in; // @[stackmanage_35.scala 48:47]
  wire [31:0] Stack_14_io_hit_out; // @[stackmanage_35.scala 48:47]
  wire [31:0] Stack_14_io_ray_out; // @[stackmanage_35.scala 48:47]
  wire  Stack_14_io_enable; // @[stackmanage_35.scala 48:47]
  wire  Stack_15_clock; // @[stackmanage_35.scala 49:47]
  wire  Stack_15_reset; // @[stackmanage_35.scala 49:47]
  wire  Stack_15_io_push; // @[stackmanage_35.scala 49:47]
  wire  Stack_15_io_pop; // @[stackmanage_35.scala 49:47]
  wire [31:0] Stack_15_io_dataIn; // @[stackmanage_35.scala 49:47]
  wire [31:0] Stack_15_io_ray_id; // @[stackmanage_35.scala 49:47]
  wire [31:0] Stack_15_io_dataOut; // @[stackmanage_35.scala 49:47]
  wire  Stack_15_io_empty; // @[stackmanage_35.scala 49:47]
  wire [31:0] Stack_15_io_hit_in; // @[stackmanage_35.scala 49:47]
  wire [31:0] Stack_15_io_hit_out; // @[stackmanage_35.scala 49:47]
  wire [31:0] Stack_15_io_ray_out; // @[stackmanage_35.scala 49:47]
  wire  Stack_15_io_enable; // @[stackmanage_35.scala 49:47]
  wire  Stack_16_clock; // @[stackmanage_35.scala 50:49]
  wire  Stack_16_reset; // @[stackmanage_35.scala 50:49]
  wire  Stack_16_io_push; // @[stackmanage_35.scala 50:49]
  wire  Stack_16_io_pop; // @[stackmanage_35.scala 50:49]
  wire [31:0] Stack_16_io_dataIn; // @[stackmanage_35.scala 50:49]
  wire [31:0] Stack_16_io_ray_id; // @[stackmanage_35.scala 50:49]
  wire [31:0] Stack_16_io_dataOut; // @[stackmanage_35.scala 50:49]
  wire  Stack_16_io_empty; // @[stackmanage_35.scala 50:49]
  wire [31:0] Stack_16_io_hit_in; // @[stackmanage_35.scala 50:49]
  wire [31:0] Stack_16_io_hit_out; // @[stackmanage_35.scala 50:49]
  wire [31:0] Stack_16_io_ray_out; // @[stackmanage_35.scala 50:49]
  wire  Stack_16_io_enable; // @[stackmanage_35.scala 50:49]
  wire  Stack_17_clock; // @[stackmanage_35.scala 51:49]
  wire  Stack_17_reset; // @[stackmanage_35.scala 51:49]
  wire  Stack_17_io_push; // @[stackmanage_35.scala 51:49]
  wire  Stack_17_io_pop; // @[stackmanage_35.scala 51:49]
  wire [31:0] Stack_17_io_dataIn; // @[stackmanage_35.scala 51:49]
  wire [31:0] Stack_17_io_ray_id; // @[stackmanage_35.scala 51:49]
  wire [31:0] Stack_17_io_dataOut; // @[stackmanage_35.scala 51:49]
  wire  Stack_17_io_empty; // @[stackmanage_35.scala 51:49]
  wire [31:0] Stack_17_io_hit_in; // @[stackmanage_35.scala 51:49]
  wire [31:0] Stack_17_io_hit_out; // @[stackmanage_35.scala 51:49]
  wire [31:0] Stack_17_io_ray_out; // @[stackmanage_35.scala 51:49]
  wire  Stack_17_io_enable; // @[stackmanage_35.scala 51:49]
  wire  Stack_18_clock; // @[stackmanage_35.scala 52:49]
  wire  Stack_18_reset; // @[stackmanage_35.scala 52:49]
  wire  Stack_18_io_push; // @[stackmanage_35.scala 52:49]
  wire  Stack_18_io_pop; // @[stackmanage_35.scala 52:49]
  wire [31:0] Stack_18_io_dataIn; // @[stackmanage_35.scala 52:49]
  wire [31:0] Stack_18_io_ray_id; // @[stackmanage_35.scala 52:49]
  wire [31:0] Stack_18_io_dataOut; // @[stackmanage_35.scala 52:49]
  wire  Stack_18_io_empty; // @[stackmanage_35.scala 52:49]
  wire [31:0] Stack_18_io_hit_in; // @[stackmanage_35.scala 52:49]
  wire [31:0] Stack_18_io_hit_out; // @[stackmanage_35.scala 52:49]
  wire [31:0] Stack_18_io_ray_out; // @[stackmanage_35.scala 52:49]
  wire  Stack_18_io_enable; // @[stackmanage_35.scala 52:49]
  wire  Stack_19_clock; // @[stackmanage_35.scala 53:49]
  wire  Stack_19_reset; // @[stackmanage_35.scala 53:49]
  wire  Stack_19_io_push; // @[stackmanage_35.scala 53:49]
  wire  Stack_19_io_pop; // @[stackmanage_35.scala 53:49]
  wire [31:0] Stack_19_io_dataIn; // @[stackmanage_35.scala 53:49]
  wire [31:0] Stack_19_io_ray_id; // @[stackmanage_35.scala 53:49]
  wire [31:0] Stack_19_io_dataOut; // @[stackmanage_35.scala 53:49]
  wire  Stack_19_io_empty; // @[stackmanage_35.scala 53:49]
  wire [31:0] Stack_19_io_hit_in; // @[stackmanage_35.scala 53:49]
  wire [31:0] Stack_19_io_hit_out; // @[stackmanage_35.scala 53:49]
  wire [31:0] Stack_19_io_ray_out; // @[stackmanage_35.scala 53:49]
  wire  Stack_19_io_enable; // @[stackmanage_35.scala 53:49]
  wire  Stack_20_clock; // @[stackmanage_35.scala 54:49]
  wire  Stack_20_reset; // @[stackmanage_35.scala 54:49]
  wire  Stack_20_io_push; // @[stackmanage_35.scala 54:49]
  wire  Stack_20_io_pop; // @[stackmanage_35.scala 54:49]
  wire [31:0] Stack_20_io_dataIn; // @[stackmanage_35.scala 54:49]
  wire [31:0] Stack_20_io_ray_id; // @[stackmanage_35.scala 54:49]
  wire [31:0] Stack_20_io_dataOut; // @[stackmanage_35.scala 54:49]
  wire  Stack_20_io_empty; // @[stackmanage_35.scala 54:49]
  wire [31:0] Stack_20_io_hit_in; // @[stackmanage_35.scala 54:49]
  wire [31:0] Stack_20_io_hit_out; // @[stackmanage_35.scala 54:49]
  wire [31:0] Stack_20_io_ray_out; // @[stackmanage_35.scala 54:49]
  wire  Stack_20_io_enable; // @[stackmanage_35.scala 54:49]
  wire  Stack_21_clock; // @[stackmanage_35.scala 55:49]
  wire  Stack_21_reset; // @[stackmanage_35.scala 55:49]
  wire  Stack_21_io_push; // @[stackmanage_35.scala 55:49]
  wire  Stack_21_io_pop; // @[stackmanage_35.scala 55:49]
  wire [31:0] Stack_21_io_dataIn; // @[stackmanage_35.scala 55:49]
  wire [31:0] Stack_21_io_ray_id; // @[stackmanage_35.scala 55:49]
  wire [31:0] Stack_21_io_dataOut; // @[stackmanage_35.scala 55:49]
  wire  Stack_21_io_empty; // @[stackmanage_35.scala 55:49]
  wire [31:0] Stack_21_io_hit_in; // @[stackmanage_35.scala 55:49]
  wire [31:0] Stack_21_io_hit_out; // @[stackmanage_35.scala 55:49]
  wire [31:0] Stack_21_io_ray_out; // @[stackmanage_35.scala 55:49]
  wire  Stack_21_io_enable; // @[stackmanage_35.scala 55:49]
  wire  Stack_22_clock; // @[stackmanage_35.scala 56:49]
  wire  Stack_22_reset; // @[stackmanage_35.scala 56:49]
  wire  Stack_22_io_push; // @[stackmanage_35.scala 56:49]
  wire  Stack_22_io_pop; // @[stackmanage_35.scala 56:49]
  wire [31:0] Stack_22_io_dataIn; // @[stackmanage_35.scala 56:49]
  wire [31:0] Stack_22_io_ray_id; // @[stackmanage_35.scala 56:49]
  wire [31:0] Stack_22_io_dataOut; // @[stackmanage_35.scala 56:49]
  wire  Stack_22_io_empty; // @[stackmanage_35.scala 56:49]
  wire [31:0] Stack_22_io_hit_in; // @[stackmanage_35.scala 56:49]
  wire [31:0] Stack_22_io_hit_out; // @[stackmanage_35.scala 56:49]
  wire [31:0] Stack_22_io_ray_out; // @[stackmanage_35.scala 56:49]
  wire  Stack_22_io_enable; // @[stackmanage_35.scala 56:49]
  wire  Stack_23_clock; // @[stackmanage_35.scala 57:48]
  wire  Stack_23_reset; // @[stackmanage_35.scala 57:48]
  wire  Stack_23_io_push; // @[stackmanage_35.scala 57:48]
  wire  Stack_23_io_pop; // @[stackmanage_35.scala 57:48]
  wire [31:0] Stack_23_io_dataIn; // @[stackmanage_35.scala 57:48]
  wire [31:0] Stack_23_io_ray_id; // @[stackmanage_35.scala 57:48]
  wire [31:0] Stack_23_io_dataOut; // @[stackmanage_35.scala 57:48]
  wire  Stack_23_io_empty; // @[stackmanage_35.scala 57:48]
  wire [31:0] Stack_23_io_hit_in; // @[stackmanage_35.scala 57:48]
  wire [31:0] Stack_23_io_hit_out; // @[stackmanage_35.scala 57:48]
  wire [31:0] Stack_23_io_ray_out; // @[stackmanage_35.scala 57:48]
  wire  Stack_23_io_enable; // @[stackmanage_35.scala 57:48]
  wire  Stack_24_clock; // @[stackmanage_35.scala 58:48]
  wire  Stack_24_reset; // @[stackmanage_35.scala 58:48]
  wire  Stack_24_io_push; // @[stackmanage_35.scala 58:48]
  wire  Stack_24_io_pop; // @[stackmanage_35.scala 58:48]
  wire [31:0] Stack_24_io_dataIn; // @[stackmanage_35.scala 58:48]
  wire [31:0] Stack_24_io_ray_id; // @[stackmanage_35.scala 58:48]
  wire [31:0] Stack_24_io_dataOut; // @[stackmanage_35.scala 58:48]
  wire  Stack_24_io_empty; // @[stackmanage_35.scala 58:48]
  wire [31:0] Stack_24_io_hit_in; // @[stackmanage_35.scala 58:48]
  wire [31:0] Stack_24_io_hit_out; // @[stackmanage_35.scala 58:48]
  wire [31:0] Stack_24_io_ray_out; // @[stackmanage_35.scala 58:48]
  wire  Stack_24_io_enable; // @[stackmanage_35.scala 58:48]
  wire  Stack_25_clock; // @[stackmanage_35.scala 59:49]
  wire  Stack_25_reset; // @[stackmanage_35.scala 59:49]
  wire  Stack_25_io_push; // @[stackmanage_35.scala 59:49]
  wire  Stack_25_io_pop; // @[stackmanage_35.scala 59:49]
  wire [31:0] Stack_25_io_dataIn; // @[stackmanage_35.scala 59:49]
  wire [31:0] Stack_25_io_ray_id; // @[stackmanage_35.scala 59:49]
  wire [31:0] Stack_25_io_dataOut; // @[stackmanage_35.scala 59:49]
  wire  Stack_25_io_empty; // @[stackmanage_35.scala 59:49]
  wire [31:0] Stack_25_io_hit_in; // @[stackmanage_35.scala 59:49]
  wire [31:0] Stack_25_io_hit_out; // @[stackmanage_35.scala 59:49]
  wire [31:0] Stack_25_io_ray_out; // @[stackmanage_35.scala 59:49]
  wire  Stack_25_io_enable; // @[stackmanage_35.scala 59:49]
  wire  Stack_26_clock; // @[stackmanage_35.scala 60:47]
  wire  Stack_26_reset; // @[stackmanage_35.scala 60:47]
  wire  Stack_26_io_push; // @[stackmanage_35.scala 60:47]
  wire  Stack_26_io_pop; // @[stackmanage_35.scala 60:47]
  wire [31:0] Stack_26_io_dataIn; // @[stackmanage_35.scala 60:47]
  wire [31:0] Stack_26_io_ray_id; // @[stackmanage_35.scala 60:47]
  wire [31:0] Stack_26_io_dataOut; // @[stackmanage_35.scala 60:47]
  wire  Stack_26_io_empty; // @[stackmanage_35.scala 60:47]
  wire [31:0] Stack_26_io_hit_in; // @[stackmanage_35.scala 60:47]
  wire [31:0] Stack_26_io_hit_out; // @[stackmanage_35.scala 60:47]
  wire [31:0] Stack_26_io_ray_out; // @[stackmanage_35.scala 60:47]
  wire  Stack_26_io_enable; // @[stackmanage_35.scala 60:47]
  wire  Stack_27_clock; // @[stackmanage_35.scala 61:47]
  wire  Stack_27_reset; // @[stackmanage_35.scala 61:47]
  wire  Stack_27_io_push; // @[stackmanage_35.scala 61:47]
  wire  Stack_27_io_pop; // @[stackmanage_35.scala 61:47]
  wire [31:0] Stack_27_io_dataIn; // @[stackmanage_35.scala 61:47]
  wire [31:0] Stack_27_io_ray_id; // @[stackmanage_35.scala 61:47]
  wire [31:0] Stack_27_io_dataOut; // @[stackmanage_35.scala 61:47]
  wire  Stack_27_io_empty; // @[stackmanage_35.scala 61:47]
  wire [31:0] Stack_27_io_hit_in; // @[stackmanage_35.scala 61:47]
  wire [31:0] Stack_27_io_hit_out; // @[stackmanage_35.scala 61:47]
  wire [31:0] Stack_27_io_ray_out; // @[stackmanage_35.scala 61:47]
  wire  Stack_27_io_enable; // @[stackmanage_35.scala 61:47]
  wire  Stack_28_clock; // @[stackmanage_35.scala 62:47]
  wire  Stack_28_reset; // @[stackmanage_35.scala 62:47]
  wire  Stack_28_io_push; // @[stackmanage_35.scala 62:47]
  wire  Stack_28_io_pop; // @[stackmanage_35.scala 62:47]
  wire [31:0] Stack_28_io_dataIn; // @[stackmanage_35.scala 62:47]
  wire [31:0] Stack_28_io_ray_id; // @[stackmanage_35.scala 62:47]
  wire [31:0] Stack_28_io_dataOut; // @[stackmanage_35.scala 62:47]
  wire  Stack_28_io_empty; // @[stackmanage_35.scala 62:47]
  wire [31:0] Stack_28_io_hit_in; // @[stackmanage_35.scala 62:47]
  wire [31:0] Stack_28_io_hit_out; // @[stackmanage_35.scala 62:47]
  wire [31:0] Stack_28_io_ray_out; // @[stackmanage_35.scala 62:47]
  wire  Stack_28_io_enable; // @[stackmanage_35.scala 62:47]
  wire  Stack_29_clock; // @[stackmanage_35.scala 63:47]
  wire  Stack_29_reset; // @[stackmanage_35.scala 63:47]
  wire  Stack_29_io_push; // @[stackmanage_35.scala 63:47]
  wire  Stack_29_io_pop; // @[stackmanage_35.scala 63:47]
  wire [31:0] Stack_29_io_dataIn; // @[stackmanage_35.scala 63:47]
  wire [31:0] Stack_29_io_ray_id; // @[stackmanage_35.scala 63:47]
  wire [31:0] Stack_29_io_dataOut; // @[stackmanage_35.scala 63:47]
  wire  Stack_29_io_empty; // @[stackmanage_35.scala 63:47]
  wire [31:0] Stack_29_io_hit_in; // @[stackmanage_35.scala 63:47]
  wire [31:0] Stack_29_io_hit_out; // @[stackmanage_35.scala 63:47]
  wire [31:0] Stack_29_io_ray_out; // @[stackmanage_35.scala 63:47]
  wire  Stack_29_io_enable; // @[stackmanage_35.scala 63:47]
  wire  Stack_30_clock; // @[stackmanage_35.scala 64:47]
  wire  Stack_30_reset; // @[stackmanage_35.scala 64:47]
  wire  Stack_30_io_push; // @[stackmanage_35.scala 64:47]
  wire  Stack_30_io_pop; // @[stackmanage_35.scala 64:47]
  wire [31:0] Stack_30_io_dataIn; // @[stackmanage_35.scala 64:47]
  wire [31:0] Stack_30_io_ray_id; // @[stackmanage_35.scala 64:47]
  wire [31:0] Stack_30_io_dataOut; // @[stackmanage_35.scala 64:47]
  wire  Stack_30_io_empty; // @[stackmanage_35.scala 64:47]
  wire [31:0] Stack_30_io_hit_in; // @[stackmanage_35.scala 64:47]
  wire [31:0] Stack_30_io_hit_out; // @[stackmanage_35.scala 64:47]
  wire [31:0] Stack_30_io_ray_out; // @[stackmanage_35.scala 64:47]
  wire  Stack_30_io_enable; // @[stackmanage_35.scala 64:47]
  wire  Stack_31_clock; // @[stackmanage_35.scala 65:47]
  wire  Stack_31_reset; // @[stackmanage_35.scala 65:47]
  wire  Stack_31_io_push; // @[stackmanage_35.scala 65:47]
  wire  Stack_31_io_pop; // @[stackmanage_35.scala 65:47]
  wire [31:0] Stack_31_io_dataIn; // @[stackmanage_35.scala 65:47]
  wire [31:0] Stack_31_io_ray_id; // @[stackmanage_35.scala 65:47]
  wire [31:0] Stack_31_io_dataOut; // @[stackmanage_35.scala 65:47]
  wire  Stack_31_io_empty; // @[stackmanage_35.scala 65:47]
  wire [31:0] Stack_31_io_hit_in; // @[stackmanage_35.scala 65:47]
  wire [31:0] Stack_31_io_hit_out; // @[stackmanage_35.scala 65:47]
  wire [31:0] Stack_31_io_ray_out; // @[stackmanage_35.scala 65:47]
  wire  Stack_31_io_enable; // @[stackmanage_35.scala 65:47]
  wire  Stack_32_clock; // @[stackmanage_35.scala 66:49]
  wire  Stack_32_reset; // @[stackmanage_35.scala 66:49]
  wire  Stack_32_io_push; // @[stackmanage_35.scala 66:49]
  wire  Stack_32_io_pop; // @[stackmanage_35.scala 66:49]
  wire [31:0] Stack_32_io_dataIn; // @[stackmanage_35.scala 66:49]
  wire [31:0] Stack_32_io_ray_id; // @[stackmanage_35.scala 66:49]
  wire [31:0] Stack_32_io_dataOut; // @[stackmanage_35.scala 66:49]
  wire  Stack_32_io_empty; // @[stackmanage_35.scala 66:49]
  wire [31:0] Stack_32_io_hit_in; // @[stackmanage_35.scala 66:49]
  wire [31:0] Stack_32_io_hit_out; // @[stackmanage_35.scala 66:49]
  wire [31:0] Stack_32_io_ray_out; // @[stackmanage_35.scala 66:49]
  wire  Stack_32_io_enable; // @[stackmanage_35.scala 66:49]
  wire  Stack_33_clock; // @[stackmanage_35.scala 67:48]
  wire  Stack_33_reset; // @[stackmanage_35.scala 67:48]
  wire  Stack_33_io_push; // @[stackmanage_35.scala 67:48]
  wire  Stack_33_io_pop; // @[stackmanage_35.scala 67:48]
  wire [31:0] Stack_33_io_dataIn; // @[stackmanage_35.scala 67:48]
  wire [31:0] Stack_33_io_ray_id; // @[stackmanage_35.scala 67:48]
  wire [31:0] Stack_33_io_dataOut; // @[stackmanage_35.scala 67:48]
  wire  Stack_33_io_empty; // @[stackmanage_35.scala 67:48]
  wire [31:0] Stack_33_io_hit_in; // @[stackmanage_35.scala 67:48]
  wire [31:0] Stack_33_io_hit_out; // @[stackmanage_35.scala 67:48]
  wire [31:0] Stack_33_io_ray_out; // @[stackmanage_35.scala 67:48]
  wire  Stack_33_io_enable; // @[stackmanage_35.scala 67:48]
  wire  Stack_34_clock; // @[stackmanage_35.scala 68:48]
  wire  Stack_34_reset; // @[stackmanage_35.scala 68:48]
  wire  Stack_34_io_push; // @[stackmanage_35.scala 68:48]
  wire  Stack_34_io_pop; // @[stackmanage_35.scala 68:48]
  wire [31:0] Stack_34_io_dataIn; // @[stackmanage_35.scala 68:48]
  wire [31:0] Stack_34_io_ray_id; // @[stackmanage_35.scala 68:48]
  wire [31:0] Stack_34_io_dataOut; // @[stackmanage_35.scala 68:48]
  wire  Stack_34_io_empty; // @[stackmanage_35.scala 68:48]
  wire [31:0] Stack_34_io_hit_in; // @[stackmanage_35.scala 68:48]
  wire [31:0] Stack_34_io_hit_out; // @[stackmanage_35.scala 68:48]
  wire [31:0] Stack_34_io_ray_out; // @[stackmanage_35.scala 68:48]
  wire  Stack_34_io_enable; // @[stackmanage_35.scala 68:48]
  reg [31:0] node_push_in_1; // @[stackmanage_35.scala 331:34]
  reg [31:0] node_push_in_2; // @[stackmanage_35.scala 332:34]
  wire  _T_1 = LUT_stack_io_push_en; // @[stackmanage_35.scala 339:57]
  wire [31:0] _GEN_0 = LUT_stack_io_push_34 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 1563:71 stackmanage_35.scala 1564:30 stackmanage_35.scala 1634:31]
  wire [31:0] _GEN_2 = LUT_stack_io_push_33 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 1527:71 stackmanage_35.scala 1528:30]
  wire [31:0] _GEN_4 = LUT_stack_io_push_33 & _T_1 ? $signed(32'sh0) : $signed(_GEN_0); // @[stackmanage_35.scala 1527:71 stackmanage_35.scala 1562:31]
  wire [31:0] _GEN_5 = LUT_stack_io_push_32 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 1491:71 stackmanage_35.scala 1492:30]
  wire [31:0] _GEN_7 = LUT_stack_io_push_32 & _T_1 ? $signed(32'sh0) : $signed(_GEN_2); // @[stackmanage_35.scala 1491:71 stackmanage_35.scala 1525:31]
  wire [31:0] _GEN_8 = LUT_stack_io_push_32 & _T_1 ? $signed(32'sh0) : $signed(_GEN_4); // @[stackmanage_35.scala 1491:71 stackmanage_35.scala 1526:31]
  wire [31:0] _GEN_9 = LUT_stack_io_push_31 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 1455:72 stackmanage_35.scala 1456:30]
  wire [31:0] _GEN_11 = LUT_stack_io_push_31 & _T_1 ? $signed(32'sh0) : $signed(_GEN_5); // @[stackmanage_35.scala 1455:72 stackmanage_35.scala 1488:31]
  wire [31:0] _GEN_12 = LUT_stack_io_push_31 & _T_1 ? $signed(32'sh0) : $signed(_GEN_7); // @[stackmanage_35.scala 1455:72 stackmanage_35.scala 1489:31]
  wire [31:0] _GEN_13 = LUT_stack_io_push_31 & _T_1 ? $signed(32'sh0) : $signed(_GEN_8); // @[stackmanage_35.scala 1455:72 stackmanage_35.scala 1490:31]
  wire [31:0] _GEN_14 = LUT_stack_io_push_30 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 1419:72 stackmanage_35.scala 1420:30]
  wire [31:0] _GEN_16 = LUT_stack_io_push_30 & _T_1 ? $signed(32'sh0) : $signed(_GEN_9); // @[stackmanage_35.scala 1419:72 stackmanage_35.scala 1451:31]
  wire [31:0] _GEN_17 = LUT_stack_io_push_30 & _T_1 ? $signed(32'sh0) : $signed(_GEN_11); // @[stackmanage_35.scala 1419:72 stackmanage_35.scala 1452:31]
  wire [31:0] _GEN_18 = LUT_stack_io_push_30 & _T_1 ? $signed(32'sh0) : $signed(_GEN_12); // @[stackmanage_35.scala 1419:72 stackmanage_35.scala 1453:31]
  wire [31:0] _GEN_19 = LUT_stack_io_push_30 & _T_1 ? $signed(32'sh0) : $signed(_GEN_13); // @[stackmanage_35.scala 1419:72 stackmanage_35.scala 1454:31]
  wire [31:0] _GEN_20 = LUT_stack_io_push_29 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 1383:72 stackmanage_35.scala 1384:30]
  wire [31:0] _GEN_22 = LUT_stack_io_push_29 & _T_1 ? $signed(32'sh0) : $signed(_GEN_14); // @[stackmanage_35.scala 1383:72 stackmanage_35.scala 1414:31]
  wire [31:0] _GEN_23 = LUT_stack_io_push_29 & _T_1 ? $signed(32'sh0) : $signed(_GEN_16); // @[stackmanage_35.scala 1383:72 stackmanage_35.scala 1415:31]
  wire [31:0] _GEN_24 = LUT_stack_io_push_29 & _T_1 ? $signed(32'sh0) : $signed(_GEN_17); // @[stackmanage_35.scala 1383:72 stackmanage_35.scala 1416:31]
  wire [31:0] _GEN_25 = LUT_stack_io_push_29 & _T_1 ? $signed(32'sh0) : $signed(_GEN_18); // @[stackmanage_35.scala 1383:72 stackmanage_35.scala 1417:31]
  wire [31:0] _GEN_26 = LUT_stack_io_push_29 & _T_1 ? $signed(32'sh0) : $signed(_GEN_19); // @[stackmanage_35.scala 1383:72 stackmanage_35.scala 1418:31]
  wire [31:0] _GEN_27 = LUT_stack_io_push_28 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 1347:72 stackmanage_35.scala 1348:30]
  wire [31:0] _GEN_29 = LUT_stack_io_push_28 & _T_1 ? $signed(32'sh0) : $signed(_GEN_20); // @[stackmanage_35.scala 1347:72 stackmanage_35.scala 1377:31]
  wire [31:0] _GEN_30 = LUT_stack_io_push_28 & _T_1 ? $signed(32'sh0) : $signed(_GEN_22); // @[stackmanage_35.scala 1347:72 stackmanage_35.scala 1378:31]
  wire [31:0] _GEN_31 = LUT_stack_io_push_28 & _T_1 ? $signed(32'sh0) : $signed(_GEN_23); // @[stackmanage_35.scala 1347:72 stackmanage_35.scala 1379:31]
  wire [31:0] _GEN_32 = LUT_stack_io_push_28 & _T_1 ? $signed(32'sh0) : $signed(_GEN_24); // @[stackmanage_35.scala 1347:72 stackmanage_35.scala 1380:31]
  wire [31:0] _GEN_33 = LUT_stack_io_push_28 & _T_1 ? $signed(32'sh0) : $signed(_GEN_25); // @[stackmanage_35.scala 1347:72 stackmanage_35.scala 1381:31]
  wire [31:0] _GEN_34 = LUT_stack_io_push_28 & _T_1 ? $signed(32'sh0) : $signed(_GEN_26); // @[stackmanage_35.scala 1347:72 stackmanage_35.scala 1382:31]
  wire [31:0] _GEN_35 = LUT_stack_io_push_27 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 1311:72 stackmanage_35.scala 1312:30]
  wire [31:0] _GEN_37 = LUT_stack_io_push_27 & _T_1 ? $signed(32'sh0) : $signed(_GEN_27); // @[stackmanage_35.scala 1311:72 stackmanage_35.scala 1340:31]
  wire [31:0] _GEN_38 = LUT_stack_io_push_27 & _T_1 ? $signed(32'sh0) : $signed(_GEN_29); // @[stackmanage_35.scala 1311:72 stackmanage_35.scala 1341:31]
  wire [31:0] _GEN_39 = LUT_stack_io_push_27 & _T_1 ? $signed(32'sh0) : $signed(_GEN_30); // @[stackmanage_35.scala 1311:72 stackmanage_35.scala 1342:31]
  wire [31:0] _GEN_40 = LUT_stack_io_push_27 & _T_1 ? $signed(32'sh0) : $signed(_GEN_31); // @[stackmanage_35.scala 1311:72 stackmanage_35.scala 1343:31]
  wire [31:0] _GEN_41 = LUT_stack_io_push_27 & _T_1 ? $signed(32'sh0) : $signed(_GEN_32); // @[stackmanage_35.scala 1311:72 stackmanage_35.scala 1344:31]
  wire [31:0] _GEN_42 = LUT_stack_io_push_27 & _T_1 ? $signed(32'sh0) : $signed(_GEN_33); // @[stackmanage_35.scala 1311:72 stackmanage_35.scala 1345:31]
  wire [31:0] _GEN_43 = LUT_stack_io_push_27 & _T_1 ? $signed(32'sh0) : $signed(_GEN_34); // @[stackmanage_35.scala 1311:72 stackmanage_35.scala 1346:31]
  wire [31:0] _GEN_44 = LUT_stack_io_push_26 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 1275:71 stackmanage_35.scala 1276:30]
  wire [31:0] _GEN_46 = LUT_stack_io_push_26 & _T_1 ? $signed(32'sh0) : $signed(_GEN_35); // @[stackmanage_35.scala 1275:71 stackmanage_35.scala 1303:31]
  wire [31:0] _GEN_47 = LUT_stack_io_push_26 & _T_1 ? $signed(32'sh0) : $signed(_GEN_37); // @[stackmanage_35.scala 1275:71 stackmanage_35.scala 1304:31]
  wire [31:0] _GEN_48 = LUT_stack_io_push_26 & _T_1 ? $signed(32'sh0) : $signed(_GEN_38); // @[stackmanage_35.scala 1275:71 stackmanage_35.scala 1305:31]
  wire [31:0] _GEN_49 = LUT_stack_io_push_26 & _T_1 ? $signed(32'sh0) : $signed(_GEN_39); // @[stackmanage_35.scala 1275:71 stackmanage_35.scala 1306:31]
  wire [31:0] _GEN_50 = LUT_stack_io_push_26 & _T_1 ? $signed(32'sh0) : $signed(_GEN_40); // @[stackmanage_35.scala 1275:71 stackmanage_35.scala 1307:31]
  wire [31:0] _GEN_51 = LUT_stack_io_push_26 & _T_1 ? $signed(32'sh0) : $signed(_GEN_41); // @[stackmanage_35.scala 1275:71 stackmanage_35.scala 1308:31]
  wire [31:0] _GEN_52 = LUT_stack_io_push_26 & _T_1 ? $signed(32'sh0) : $signed(_GEN_42); // @[stackmanage_35.scala 1275:71 stackmanage_35.scala 1309:31]
  wire [31:0] _GEN_53 = LUT_stack_io_push_26 & _T_1 ? $signed(32'sh0) : $signed(_GEN_43); // @[stackmanage_35.scala 1275:71 stackmanage_35.scala 1310:31]
  wire [31:0] _GEN_54 = LUT_stack_io_push_25 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 1239:71 stackmanage_35.scala 1240:30]
  wire [31:0] _GEN_56 = LUT_stack_io_push_25 & _T_1 ? $signed(32'sh0) : $signed(_GEN_44); // @[stackmanage_35.scala 1239:71 stackmanage_35.scala 1266:31]
  wire [31:0] _GEN_57 = LUT_stack_io_push_25 & _T_1 ? $signed(32'sh0) : $signed(_GEN_46); // @[stackmanage_35.scala 1239:71 stackmanage_35.scala 1267:31]
  wire [31:0] _GEN_58 = LUT_stack_io_push_25 & _T_1 ? $signed(32'sh0) : $signed(_GEN_47); // @[stackmanage_35.scala 1239:71 stackmanage_35.scala 1268:31]
  wire [31:0] _GEN_59 = LUT_stack_io_push_25 & _T_1 ? $signed(32'sh0) : $signed(_GEN_48); // @[stackmanage_35.scala 1239:71 stackmanage_35.scala 1269:31]
  wire [31:0] _GEN_60 = LUT_stack_io_push_25 & _T_1 ? $signed(32'sh0) : $signed(_GEN_49); // @[stackmanage_35.scala 1239:71 stackmanage_35.scala 1270:31]
  wire [31:0] _GEN_61 = LUT_stack_io_push_25 & _T_1 ? $signed(32'sh0) : $signed(_GEN_50); // @[stackmanage_35.scala 1239:71 stackmanage_35.scala 1271:31]
  wire [31:0] _GEN_62 = LUT_stack_io_push_25 & _T_1 ? $signed(32'sh0) : $signed(_GEN_51); // @[stackmanage_35.scala 1239:71 stackmanage_35.scala 1272:31]
  wire [31:0] _GEN_63 = LUT_stack_io_push_25 & _T_1 ? $signed(32'sh0) : $signed(_GEN_52); // @[stackmanage_35.scala 1239:71 stackmanage_35.scala 1273:31]
  wire [31:0] _GEN_64 = LUT_stack_io_push_25 & _T_1 ? $signed(32'sh0) : $signed(_GEN_53); // @[stackmanage_35.scala 1239:71 stackmanage_35.scala 1274:31]
  wire [31:0] _GEN_65 = LUT_stack_io_push_24 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 1203:71 stackmanage_35.scala 1204:30]
  wire [31:0] _GEN_67 = LUT_stack_io_push_24 & _T_1 ? $signed(32'sh0) : $signed(_GEN_54); // @[stackmanage_35.scala 1203:71 stackmanage_35.scala 1229:31]
  wire [31:0] _GEN_68 = LUT_stack_io_push_24 & _T_1 ? $signed(32'sh0) : $signed(_GEN_56); // @[stackmanage_35.scala 1203:71 stackmanage_35.scala 1230:31]
  wire [31:0] _GEN_69 = LUT_stack_io_push_24 & _T_1 ? $signed(32'sh0) : $signed(_GEN_57); // @[stackmanage_35.scala 1203:71 stackmanage_35.scala 1231:31]
  wire [31:0] _GEN_70 = LUT_stack_io_push_24 & _T_1 ? $signed(32'sh0) : $signed(_GEN_58); // @[stackmanage_35.scala 1203:71 stackmanage_35.scala 1232:31]
  wire [31:0] _GEN_71 = LUT_stack_io_push_24 & _T_1 ? $signed(32'sh0) : $signed(_GEN_59); // @[stackmanage_35.scala 1203:71 stackmanage_35.scala 1233:31]
  wire [31:0] _GEN_72 = LUT_stack_io_push_24 & _T_1 ? $signed(32'sh0) : $signed(_GEN_60); // @[stackmanage_35.scala 1203:71 stackmanage_35.scala 1234:31]
  wire [31:0] _GEN_73 = LUT_stack_io_push_24 & _T_1 ? $signed(32'sh0) : $signed(_GEN_61); // @[stackmanage_35.scala 1203:71 stackmanage_35.scala 1235:31]
  wire [31:0] _GEN_74 = LUT_stack_io_push_24 & _T_1 ? $signed(32'sh0) : $signed(_GEN_62); // @[stackmanage_35.scala 1203:71 stackmanage_35.scala 1236:31]
  wire [31:0] _GEN_75 = LUT_stack_io_push_24 & _T_1 ? $signed(32'sh0) : $signed(_GEN_63); // @[stackmanage_35.scala 1203:71 stackmanage_35.scala 1237:31]
  wire [31:0] _GEN_76 = LUT_stack_io_push_24 & _T_1 ? $signed(32'sh0) : $signed(_GEN_64); // @[stackmanage_35.scala 1203:71 stackmanage_35.scala 1238:31]
  wire [31:0] _GEN_77 = LUT_stack_io_push_23 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 1167:71 stackmanage_35.scala 1168:30]
  wire [31:0] _GEN_79 = LUT_stack_io_push_23 & _T_1 ? $signed(32'sh0) : $signed(_GEN_65); // @[stackmanage_35.scala 1167:71 stackmanage_35.scala 1192:31]
  wire [31:0] _GEN_80 = LUT_stack_io_push_23 & _T_1 ? $signed(32'sh0) : $signed(_GEN_67); // @[stackmanage_35.scala 1167:71 stackmanage_35.scala 1193:31]
  wire [31:0] _GEN_81 = LUT_stack_io_push_23 & _T_1 ? $signed(32'sh0) : $signed(_GEN_68); // @[stackmanage_35.scala 1167:71 stackmanage_35.scala 1194:31]
  wire [31:0] _GEN_82 = LUT_stack_io_push_23 & _T_1 ? $signed(32'sh0) : $signed(_GEN_69); // @[stackmanage_35.scala 1167:71 stackmanage_35.scala 1195:31]
  wire [31:0] _GEN_83 = LUT_stack_io_push_23 & _T_1 ? $signed(32'sh0) : $signed(_GEN_70); // @[stackmanage_35.scala 1167:71 stackmanage_35.scala 1196:31]
  wire [31:0] _GEN_84 = LUT_stack_io_push_23 & _T_1 ? $signed(32'sh0) : $signed(_GEN_71); // @[stackmanage_35.scala 1167:71 stackmanage_35.scala 1197:31]
  wire [31:0] _GEN_85 = LUT_stack_io_push_23 & _T_1 ? $signed(32'sh0) : $signed(_GEN_72); // @[stackmanage_35.scala 1167:71 stackmanage_35.scala 1198:31]
  wire [31:0] _GEN_86 = LUT_stack_io_push_23 & _T_1 ? $signed(32'sh0) : $signed(_GEN_73); // @[stackmanage_35.scala 1167:71 stackmanage_35.scala 1199:31]
  wire [31:0] _GEN_87 = LUT_stack_io_push_23 & _T_1 ? $signed(32'sh0) : $signed(_GEN_74); // @[stackmanage_35.scala 1167:71 stackmanage_35.scala 1200:31]
  wire [31:0] _GEN_88 = LUT_stack_io_push_23 & _T_1 ? $signed(32'sh0) : $signed(_GEN_75); // @[stackmanage_35.scala 1167:71 stackmanage_35.scala 1201:31]
  wire [31:0] _GEN_89 = LUT_stack_io_push_23 & _T_1 ? $signed(32'sh0) : $signed(_GEN_76); // @[stackmanage_35.scala 1167:71 stackmanage_35.scala 1202:31]
  wire [31:0] _GEN_90 = LUT_stack_io_push_22 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 1131:71 stackmanage_35.scala 1132:30]
  wire [31:0] _GEN_92 = LUT_stack_io_push_22 & _T_1 ? $signed(32'sh0) : $signed(_GEN_77); // @[stackmanage_35.scala 1131:71 stackmanage_35.scala 1155:31]
  wire [31:0] _GEN_93 = LUT_stack_io_push_22 & _T_1 ? $signed(32'sh0) : $signed(_GEN_79); // @[stackmanage_35.scala 1131:71 stackmanage_35.scala 1156:31]
  wire [31:0] _GEN_94 = LUT_stack_io_push_22 & _T_1 ? $signed(32'sh0) : $signed(_GEN_80); // @[stackmanage_35.scala 1131:71 stackmanage_35.scala 1157:31]
  wire [31:0] _GEN_95 = LUT_stack_io_push_22 & _T_1 ? $signed(32'sh0) : $signed(_GEN_81); // @[stackmanage_35.scala 1131:71 stackmanage_35.scala 1158:31]
  wire [31:0] _GEN_96 = LUT_stack_io_push_22 & _T_1 ? $signed(32'sh0) : $signed(_GEN_82); // @[stackmanage_35.scala 1131:71 stackmanage_35.scala 1159:31]
  wire [31:0] _GEN_97 = LUT_stack_io_push_22 & _T_1 ? $signed(32'sh0) : $signed(_GEN_83); // @[stackmanage_35.scala 1131:71 stackmanage_35.scala 1160:31]
  wire [31:0] _GEN_98 = LUT_stack_io_push_22 & _T_1 ? $signed(32'sh0) : $signed(_GEN_84); // @[stackmanage_35.scala 1131:71 stackmanage_35.scala 1161:31]
  wire [31:0] _GEN_99 = LUT_stack_io_push_22 & _T_1 ? $signed(32'sh0) : $signed(_GEN_85); // @[stackmanage_35.scala 1131:71 stackmanage_35.scala 1162:31]
  wire [31:0] _GEN_100 = LUT_stack_io_push_22 & _T_1 ? $signed(32'sh0) : $signed(_GEN_86); // @[stackmanage_35.scala 1131:71 stackmanage_35.scala 1163:31]
  wire [31:0] _GEN_101 = LUT_stack_io_push_22 & _T_1 ? $signed(32'sh0) : $signed(_GEN_87); // @[stackmanage_35.scala 1131:71 stackmanage_35.scala 1164:31]
  wire [31:0] _GEN_102 = LUT_stack_io_push_22 & _T_1 ? $signed(32'sh0) : $signed(_GEN_88); // @[stackmanage_35.scala 1131:71 stackmanage_35.scala 1165:31]
  wire [31:0] _GEN_103 = LUT_stack_io_push_22 & _T_1 ? $signed(32'sh0) : $signed(_GEN_89); // @[stackmanage_35.scala 1131:71 stackmanage_35.scala 1166:31]
  wire [31:0] _GEN_104 = LUT_stack_io_push_21 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 1095:71 stackmanage_35.scala 1096:30]
  wire [31:0] _GEN_106 = LUT_stack_io_push_21 & _T_1 ? $signed(32'sh0) : $signed(_GEN_90); // @[stackmanage_35.scala 1095:71 stackmanage_35.scala 1118:31]
  wire [31:0] _GEN_107 = LUT_stack_io_push_21 & _T_1 ? $signed(32'sh0) : $signed(_GEN_92); // @[stackmanage_35.scala 1095:71 stackmanage_35.scala 1119:31]
  wire [31:0] _GEN_108 = LUT_stack_io_push_21 & _T_1 ? $signed(32'sh0) : $signed(_GEN_93); // @[stackmanage_35.scala 1095:71 stackmanage_35.scala 1120:31]
  wire [31:0] _GEN_109 = LUT_stack_io_push_21 & _T_1 ? $signed(32'sh0) : $signed(_GEN_94); // @[stackmanage_35.scala 1095:71 stackmanage_35.scala 1121:31]
  wire [31:0] _GEN_110 = LUT_stack_io_push_21 & _T_1 ? $signed(32'sh0) : $signed(_GEN_95); // @[stackmanage_35.scala 1095:71 stackmanage_35.scala 1122:31]
  wire [31:0] _GEN_111 = LUT_stack_io_push_21 & _T_1 ? $signed(32'sh0) : $signed(_GEN_96); // @[stackmanage_35.scala 1095:71 stackmanage_35.scala 1123:31]
  wire [31:0] _GEN_112 = LUT_stack_io_push_21 & _T_1 ? $signed(32'sh0) : $signed(_GEN_97); // @[stackmanage_35.scala 1095:71 stackmanage_35.scala 1124:31]
  wire [31:0] _GEN_113 = LUT_stack_io_push_21 & _T_1 ? $signed(32'sh0) : $signed(_GEN_98); // @[stackmanage_35.scala 1095:71 stackmanage_35.scala 1125:31]
  wire [31:0] _GEN_114 = LUT_stack_io_push_21 & _T_1 ? $signed(32'sh0) : $signed(_GEN_99); // @[stackmanage_35.scala 1095:71 stackmanage_35.scala 1126:31]
  wire [31:0] _GEN_115 = LUT_stack_io_push_21 & _T_1 ? $signed(32'sh0) : $signed(_GEN_100); // @[stackmanage_35.scala 1095:71 stackmanage_35.scala 1127:31]
  wire [31:0] _GEN_116 = LUT_stack_io_push_21 & _T_1 ? $signed(32'sh0) : $signed(_GEN_101); // @[stackmanage_35.scala 1095:71 stackmanage_35.scala 1128:31]
  wire [31:0] _GEN_117 = LUT_stack_io_push_21 & _T_1 ? $signed(32'sh0) : $signed(_GEN_102); // @[stackmanage_35.scala 1095:71 stackmanage_35.scala 1129:31]
  wire [31:0] _GEN_118 = LUT_stack_io_push_21 & _T_1 ? $signed(32'sh0) : $signed(_GEN_103); // @[stackmanage_35.scala 1095:71 stackmanage_35.scala 1130:31]
  wire [31:0] _GEN_119 = LUT_stack_io_push_20 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 1059:71 stackmanage_35.scala 1060:30]
  wire [31:0] _GEN_121 = LUT_stack_io_push_20 & _T_1 ? $signed(32'sh0) : $signed(_GEN_104); // @[stackmanage_35.scala 1059:71 stackmanage_35.scala 1081:31]
  wire [31:0] _GEN_122 = LUT_stack_io_push_20 & _T_1 ? $signed(32'sh0) : $signed(_GEN_106); // @[stackmanage_35.scala 1059:71 stackmanage_35.scala 1082:31]
  wire [31:0] _GEN_123 = LUT_stack_io_push_20 & _T_1 ? $signed(32'sh0) : $signed(_GEN_107); // @[stackmanage_35.scala 1059:71 stackmanage_35.scala 1083:31]
  wire [31:0] _GEN_124 = LUT_stack_io_push_20 & _T_1 ? $signed(32'sh0) : $signed(_GEN_108); // @[stackmanage_35.scala 1059:71 stackmanage_35.scala 1084:31]
  wire [31:0] _GEN_125 = LUT_stack_io_push_20 & _T_1 ? $signed(32'sh0) : $signed(_GEN_109); // @[stackmanage_35.scala 1059:71 stackmanage_35.scala 1085:31]
  wire [31:0] _GEN_126 = LUT_stack_io_push_20 & _T_1 ? $signed(32'sh0) : $signed(_GEN_110); // @[stackmanage_35.scala 1059:71 stackmanage_35.scala 1086:31]
  wire [31:0] _GEN_127 = LUT_stack_io_push_20 & _T_1 ? $signed(32'sh0) : $signed(_GEN_111); // @[stackmanage_35.scala 1059:71 stackmanage_35.scala 1087:31]
  wire [31:0] _GEN_128 = LUT_stack_io_push_20 & _T_1 ? $signed(32'sh0) : $signed(_GEN_112); // @[stackmanage_35.scala 1059:71 stackmanage_35.scala 1088:31]
  wire [31:0] _GEN_129 = LUT_stack_io_push_20 & _T_1 ? $signed(32'sh0) : $signed(_GEN_113); // @[stackmanage_35.scala 1059:71 stackmanage_35.scala 1089:31]
  wire [31:0] _GEN_130 = LUT_stack_io_push_20 & _T_1 ? $signed(32'sh0) : $signed(_GEN_114); // @[stackmanage_35.scala 1059:71 stackmanage_35.scala 1090:31]
  wire [31:0] _GEN_131 = LUT_stack_io_push_20 & _T_1 ? $signed(32'sh0) : $signed(_GEN_115); // @[stackmanage_35.scala 1059:71 stackmanage_35.scala 1091:31]
  wire [31:0] _GEN_132 = LUT_stack_io_push_20 & _T_1 ? $signed(32'sh0) : $signed(_GEN_116); // @[stackmanage_35.scala 1059:71 stackmanage_35.scala 1092:31]
  wire [31:0] _GEN_133 = LUT_stack_io_push_20 & _T_1 ? $signed(32'sh0) : $signed(_GEN_117); // @[stackmanage_35.scala 1059:71 stackmanage_35.scala 1093:31]
  wire [31:0] _GEN_134 = LUT_stack_io_push_20 & _T_1 ? $signed(32'sh0) : $signed(_GEN_118); // @[stackmanage_35.scala 1059:71 stackmanage_35.scala 1094:31]
  wire [31:0] _GEN_135 = LUT_stack_io_push_19 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 1023:71 stackmanage_35.scala 1024:30]
  wire [31:0] _GEN_137 = LUT_stack_io_push_19 & _T_1 ? $signed(32'sh0) : $signed(_GEN_119); // @[stackmanage_35.scala 1023:71 stackmanage_35.scala 1044:31]
  wire [31:0] _GEN_138 = LUT_stack_io_push_19 & _T_1 ? $signed(32'sh0) : $signed(_GEN_121); // @[stackmanage_35.scala 1023:71 stackmanage_35.scala 1045:31]
  wire [31:0] _GEN_139 = LUT_stack_io_push_19 & _T_1 ? $signed(32'sh0) : $signed(_GEN_122); // @[stackmanage_35.scala 1023:71 stackmanage_35.scala 1046:31]
  wire [31:0] _GEN_140 = LUT_stack_io_push_19 & _T_1 ? $signed(32'sh0) : $signed(_GEN_123); // @[stackmanage_35.scala 1023:71 stackmanage_35.scala 1047:31]
  wire [31:0] _GEN_141 = LUT_stack_io_push_19 & _T_1 ? $signed(32'sh0) : $signed(_GEN_124); // @[stackmanage_35.scala 1023:71 stackmanage_35.scala 1048:31]
  wire [31:0] _GEN_142 = LUT_stack_io_push_19 & _T_1 ? $signed(32'sh0) : $signed(_GEN_125); // @[stackmanage_35.scala 1023:71 stackmanage_35.scala 1049:31]
  wire [31:0] _GEN_143 = LUT_stack_io_push_19 & _T_1 ? $signed(32'sh0) : $signed(_GEN_126); // @[stackmanage_35.scala 1023:71 stackmanage_35.scala 1050:31]
  wire [31:0] _GEN_144 = LUT_stack_io_push_19 & _T_1 ? $signed(32'sh0) : $signed(_GEN_127); // @[stackmanage_35.scala 1023:71 stackmanage_35.scala 1051:31]
  wire [31:0] _GEN_145 = LUT_stack_io_push_19 & _T_1 ? $signed(32'sh0) : $signed(_GEN_128); // @[stackmanage_35.scala 1023:71 stackmanage_35.scala 1052:31]
  wire [31:0] _GEN_146 = LUT_stack_io_push_19 & _T_1 ? $signed(32'sh0) : $signed(_GEN_129); // @[stackmanage_35.scala 1023:71 stackmanage_35.scala 1053:31]
  wire [31:0] _GEN_147 = LUT_stack_io_push_19 & _T_1 ? $signed(32'sh0) : $signed(_GEN_130); // @[stackmanage_35.scala 1023:71 stackmanage_35.scala 1054:31]
  wire [31:0] _GEN_148 = LUT_stack_io_push_19 & _T_1 ? $signed(32'sh0) : $signed(_GEN_131); // @[stackmanage_35.scala 1023:71 stackmanage_35.scala 1055:31]
  wire [31:0] _GEN_149 = LUT_stack_io_push_19 & _T_1 ? $signed(32'sh0) : $signed(_GEN_132); // @[stackmanage_35.scala 1023:71 stackmanage_35.scala 1056:31]
  wire [31:0] _GEN_150 = LUT_stack_io_push_19 & _T_1 ? $signed(32'sh0) : $signed(_GEN_133); // @[stackmanage_35.scala 1023:71 stackmanage_35.scala 1057:31]
  wire [31:0] _GEN_151 = LUT_stack_io_push_19 & _T_1 ? $signed(32'sh0) : $signed(_GEN_134); // @[stackmanage_35.scala 1023:71 stackmanage_35.scala 1058:31]
  wire [31:0] _GEN_152 = LUT_stack_io_push_18 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 987:71 stackmanage_35.scala 988:30]
  wire [31:0] _GEN_154 = LUT_stack_io_push_18 & _T_1 ? $signed(32'sh0) : $signed(_GEN_135); // @[stackmanage_35.scala 987:71 stackmanage_35.scala 1007:31]
  wire [31:0] _GEN_155 = LUT_stack_io_push_18 & _T_1 ? $signed(32'sh0) : $signed(_GEN_137); // @[stackmanage_35.scala 987:71 stackmanage_35.scala 1008:31]
  wire [31:0] _GEN_156 = LUT_stack_io_push_18 & _T_1 ? $signed(32'sh0) : $signed(_GEN_138); // @[stackmanage_35.scala 987:71 stackmanage_35.scala 1009:31]
  wire [31:0] _GEN_157 = LUT_stack_io_push_18 & _T_1 ? $signed(32'sh0) : $signed(_GEN_139); // @[stackmanage_35.scala 987:71 stackmanage_35.scala 1010:31]
  wire [31:0] _GEN_158 = LUT_stack_io_push_18 & _T_1 ? $signed(32'sh0) : $signed(_GEN_140); // @[stackmanage_35.scala 987:71 stackmanage_35.scala 1011:31]
  wire [31:0] _GEN_159 = LUT_stack_io_push_18 & _T_1 ? $signed(32'sh0) : $signed(_GEN_141); // @[stackmanage_35.scala 987:71 stackmanage_35.scala 1012:31]
  wire [31:0] _GEN_160 = LUT_stack_io_push_18 & _T_1 ? $signed(32'sh0) : $signed(_GEN_142); // @[stackmanage_35.scala 987:71 stackmanage_35.scala 1013:31]
  wire [31:0] _GEN_161 = LUT_stack_io_push_18 & _T_1 ? $signed(32'sh0) : $signed(_GEN_143); // @[stackmanage_35.scala 987:71 stackmanage_35.scala 1014:31]
  wire [31:0] _GEN_162 = LUT_stack_io_push_18 & _T_1 ? $signed(32'sh0) : $signed(_GEN_144); // @[stackmanage_35.scala 987:71 stackmanage_35.scala 1015:31]
  wire [31:0] _GEN_163 = LUT_stack_io_push_18 & _T_1 ? $signed(32'sh0) : $signed(_GEN_145); // @[stackmanage_35.scala 987:71 stackmanage_35.scala 1016:31]
  wire [31:0] _GEN_164 = LUT_stack_io_push_18 & _T_1 ? $signed(32'sh0) : $signed(_GEN_146); // @[stackmanage_35.scala 987:71 stackmanage_35.scala 1017:31]
  wire [31:0] _GEN_165 = LUT_stack_io_push_18 & _T_1 ? $signed(32'sh0) : $signed(_GEN_147); // @[stackmanage_35.scala 987:71 stackmanage_35.scala 1018:31]
  wire [31:0] _GEN_166 = LUT_stack_io_push_18 & _T_1 ? $signed(32'sh0) : $signed(_GEN_148); // @[stackmanage_35.scala 987:71 stackmanage_35.scala 1019:31]
  wire [31:0] _GEN_167 = LUT_stack_io_push_18 & _T_1 ? $signed(32'sh0) : $signed(_GEN_149); // @[stackmanage_35.scala 987:71 stackmanage_35.scala 1020:31]
  wire [31:0] _GEN_168 = LUT_stack_io_push_18 & _T_1 ? $signed(32'sh0) : $signed(_GEN_150); // @[stackmanage_35.scala 987:71 stackmanage_35.scala 1021:31]
  wire [31:0] _GEN_169 = LUT_stack_io_push_18 & _T_1 ? $signed(32'sh0) : $signed(_GEN_151); // @[stackmanage_35.scala 987:71 stackmanage_35.scala 1022:31]
  wire [31:0] _GEN_170 = LUT_stack_io_push_17 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 951:71 stackmanage_35.scala 952:30]
  wire [31:0] _GEN_172 = LUT_stack_io_push_17 & _T_1 ? $signed(32'sh0) : $signed(_GEN_152); // @[stackmanage_35.scala 951:71 stackmanage_35.scala 970:31]
  wire [31:0] _GEN_173 = LUT_stack_io_push_17 & _T_1 ? $signed(32'sh0) : $signed(_GEN_154); // @[stackmanage_35.scala 951:71 stackmanage_35.scala 971:31]
  wire [31:0] _GEN_174 = LUT_stack_io_push_17 & _T_1 ? $signed(32'sh0) : $signed(_GEN_155); // @[stackmanage_35.scala 951:71 stackmanage_35.scala 972:31]
  wire [31:0] _GEN_175 = LUT_stack_io_push_17 & _T_1 ? $signed(32'sh0) : $signed(_GEN_156); // @[stackmanage_35.scala 951:71 stackmanage_35.scala 973:31]
  wire [31:0] _GEN_176 = LUT_stack_io_push_17 & _T_1 ? $signed(32'sh0) : $signed(_GEN_157); // @[stackmanage_35.scala 951:71 stackmanage_35.scala 974:31]
  wire [31:0] _GEN_177 = LUT_stack_io_push_17 & _T_1 ? $signed(32'sh0) : $signed(_GEN_158); // @[stackmanage_35.scala 951:71 stackmanage_35.scala 975:31]
  wire [31:0] _GEN_178 = LUT_stack_io_push_17 & _T_1 ? $signed(32'sh0) : $signed(_GEN_159); // @[stackmanage_35.scala 951:71 stackmanage_35.scala 976:31]
  wire [31:0] _GEN_179 = LUT_stack_io_push_17 & _T_1 ? $signed(32'sh0) : $signed(_GEN_160); // @[stackmanage_35.scala 951:71 stackmanage_35.scala 977:31]
  wire [31:0] _GEN_180 = LUT_stack_io_push_17 & _T_1 ? $signed(32'sh0) : $signed(_GEN_161); // @[stackmanage_35.scala 951:71 stackmanage_35.scala 978:31]
  wire [31:0] _GEN_181 = LUT_stack_io_push_17 & _T_1 ? $signed(32'sh0) : $signed(_GEN_162); // @[stackmanage_35.scala 951:71 stackmanage_35.scala 979:31]
  wire [31:0] _GEN_182 = LUT_stack_io_push_17 & _T_1 ? $signed(32'sh0) : $signed(_GEN_163); // @[stackmanage_35.scala 951:71 stackmanage_35.scala 980:31]
  wire [31:0] _GEN_183 = LUT_stack_io_push_17 & _T_1 ? $signed(32'sh0) : $signed(_GEN_164); // @[stackmanage_35.scala 951:71 stackmanage_35.scala 981:31]
  wire [31:0] _GEN_184 = LUT_stack_io_push_17 & _T_1 ? $signed(32'sh0) : $signed(_GEN_165); // @[stackmanage_35.scala 951:71 stackmanage_35.scala 982:31]
  wire [31:0] _GEN_185 = LUT_stack_io_push_17 & _T_1 ? $signed(32'sh0) : $signed(_GEN_166); // @[stackmanage_35.scala 951:71 stackmanage_35.scala 983:31]
  wire [31:0] _GEN_186 = LUT_stack_io_push_17 & _T_1 ? $signed(32'sh0) : $signed(_GEN_167); // @[stackmanage_35.scala 951:71 stackmanage_35.scala 984:31]
  wire [31:0] _GEN_187 = LUT_stack_io_push_17 & _T_1 ? $signed(32'sh0) : $signed(_GEN_168); // @[stackmanage_35.scala 951:71 stackmanage_35.scala 985:31]
  wire [31:0] _GEN_188 = LUT_stack_io_push_17 & _T_1 ? $signed(32'sh0) : $signed(_GEN_169); // @[stackmanage_35.scala 951:71 stackmanage_35.scala 986:31]
  wire [31:0] _GEN_189 = LUT_stack_io_push_16 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 915:71 stackmanage_35.scala 916:30]
  wire [31:0] _GEN_191 = LUT_stack_io_push_16 & _T_1 ? $signed(32'sh0) : $signed(_GEN_170); // @[stackmanage_35.scala 915:71 stackmanage_35.scala 933:31]
  wire [31:0] _GEN_192 = LUT_stack_io_push_16 & _T_1 ? $signed(32'sh0) : $signed(_GEN_172); // @[stackmanage_35.scala 915:71 stackmanage_35.scala 934:31]
  wire [31:0] _GEN_193 = LUT_stack_io_push_16 & _T_1 ? $signed(32'sh0) : $signed(_GEN_173); // @[stackmanage_35.scala 915:71 stackmanage_35.scala 935:31]
  wire [31:0] _GEN_194 = LUT_stack_io_push_16 & _T_1 ? $signed(32'sh0) : $signed(_GEN_174); // @[stackmanage_35.scala 915:71 stackmanage_35.scala 936:31]
  wire [31:0] _GEN_195 = LUT_stack_io_push_16 & _T_1 ? $signed(32'sh0) : $signed(_GEN_175); // @[stackmanage_35.scala 915:71 stackmanage_35.scala 937:31]
  wire [31:0] _GEN_196 = LUT_stack_io_push_16 & _T_1 ? $signed(32'sh0) : $signed(_GEN_176); // @[stackmanage_35.scala 915:71 stackmanage_35.scala 938:31]
  wire [31:0] _GEN_197 = LUT_stack_io_push_16 & _T_1 ? $signed(32'sh0) : $signed(_GEN_177); // @[stackmanage_35.scala 915:71 stackmanage_35.scala 939:31]
  wire [31:0] _GEN_198 = LUT_stack_io_push_16 & _T_1 ? $signed(32'sh0) : $signed(_GEN_178); // @[stackmanage_35.scala 915:71 stackmanage_35.scala 940:31]
  wire [31:0] _GEN_199 = LUT_stack_io_push_16 & _T_1 ? $signed(32'sh0) : $signed(_GEN_179); // @[stackmanage_35.scala 915:71 stackmanage_35.scala 941:31]
  wire [31:0] _GEN_200 = LUT_stack_io_push_16 & _T_1 ? $signed(32'sh0) : $signed(_GEN_180); // @[stackmanage_35.scala 915:71 stackmanage_35.scala 942:31]
  wire [31:0] _GEN_201 = LUT_stack_io_push_16 & _T_1 ? $signed(32'sh0) : $signed(_GEN_181); // @[stackmanage_35.scala 915:71 stackmanage_35.scala 943:31]
  wire [31:0] _GEN_202 = LUT_stack_io_push_16 & _T_1 ? $signed(32'sh0) : $signed(_GEN_182); // @[stackmanage_35.scala 915:71 stackmanage_35.scala 944:31]
  wire [31:0] _GEN_203 = LUT_stack_io_push_16 & _T_1 ? $signed(32'sh0) : $signed(_GEN_183); // @[stackmanage_35.scala 915:71 stackmanage_35.scala 945:31]
  wire [31:0] _GEN_204 = LUT_stack_io_push_16 & _T_1 ? $signed(32'sh0) : $signed(_GEN_184); // @[stackmanage_35.scala 915:71 stackmanage_35.scala 946:31]
  wire [31:0] _GEN_205 = LUT_stack_io_push_16 & _T_1 ? $signed(32'sh0) : $signed(_GEN_185); // @[stackmanage_35.scala 915:71 stackmanage_35.scala 947:31]
  wire [31:0] _GEN_206 = LUT_stack_io_push_16 & _T_1 ? $signed(32'sh0) : $signed(_GEN_186); // @[stackmanage_35.scala 915:71 stackmanage_35.scala 948:31]
  wire [31:0] _GEN_207 = LUT_stack_io_push_16 & _T_1 ? $signed(32'sh0) : $signed(_GEN_187); // @[stackmanage_35.scala 915:71 stackmanage_35.scala 949:31]
  wire [31:0] _GEN_208 = LUT_stack_io_push_16 & _T_1 ? $signed(32'sh0) : $signed(_GEN_188); // @[stackmanage_35.scala 915:71 stackmanage_35.scala 950:31]
  wire [31:0] _GEN_209 = LUT_stack_io_push_15 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 879:71 stackmanage_35.scala 880:30]
  wire [31:0] _GEN_211 = LUT_stack_io_push_15 & _T_1 ? $signed(32'sh0) : $signed(_GEN_189); // @[stackmanage_35.scala 879:71 stackmanage_35.scala 896:31]
  wire [31:0] _GEN_212 = LUT_stack_io_push_15 & _T_1 ? $signed(32'sh0) : $signed(_GEN_191); // @[stackmanage_35.scala 879:71 stackmanage_35.scala 897:31]
  wire [31:0] _GEN_213 = LUT_stack_io_push_15 & _T_1 ? $signed(32'sh0) : $signed(_GEN_192); // @[stackmanage_35.scala 879:71 stackmanage_35.scala 898:31]
  wire [31:0] _GEN_214 = LUT_stack_io_push_15 & _T_1 ? $signed(32'sh0) : $signed(_GEN_193); // @[stackmanage_35.scala 879:71 stackmanage_35.scala 899:31]
  wire [31:0] _GEN_215 = LUT_stack_io_push_15 & _T_1 ? $signed(32'sh0) : $signed(_GEN_194); // @[stackmanage_35.scala 879:71 stackmanage_35.scala 900:31]
  wire [31:0] _GEN_216 = LUT_stack_io_push_15 & _T_1 ? $signed(32'sh0) : $signed(_GEN_195); // @[stackmanage_35.scala 879:71 stackmanage_35.scala 901:31]
  wire [31:0] _GEN_217 = LUT_stack_io_push_15 & _T_1 ? $signed(32'sh0) : $signed(_GEN_196); // @[stackmanage_35.scala 879:71 stackmanage_35.scala 902:31]
  wire [31:0] _GEN_218 = LUT_stack_io_push_15 & _T_1 ? $signed(32'sh0) : $signed(_GEN_197); // @[stackmanage_35.scala 879:71 stackmanage_35.scala 903:31]
  wire [31:0] _GEN_219 = LUT_stack_io_push_15 & _T_1 ? $signed(32'sh0) : $signed(_GEN_198); // @[stackmanage_35.scala 879:71 stackmanage_35.scala 904:31]
  wire [31:0] _GEN_220 = LUT_stack_io_push_15 & _T_1 ? $signed(32'sh0) : $signed(_GEN_199); // @[stackmanage_35.scala 879:71 stackmanage_35.scala 905:31]
  wire [31:0] _GEN_221 = LUT_stack_io_push_15 & _T_1 ? $signed(32'sh0) : $signed(_GEN_200); // @[stackmanage_35.scala 879:71 stackmanage_35.scala 906:31]
  wire [31:0] _GEN_222 = LUT_stack_io_push_15 & _T_1 ? $signed(32'sh0) : $signed(_GEN_201); // @[stackmanage_35.scala 879:71 stackmanage_35.scala 907:31]
  wire [31:0] _GEN_223 = LUT_stack_io_push_15 & _T_1 ? $signed(32'sh0) : $signed(_GEN_202); // @[stackmanage_35.scala 879:71 stackmanage_35.scala 908:31]
  wire [31:0] _GEN_224 = LUT_stack_io_push_15 & _T_1 ? $signed(32'sh0) : $signed(_GEN_203); // @[stackmanage_35.scala 879:71 stackmanage_35.scala 909:31]
  wire [31:0] _GEN_225 = LUT_stack_io_push_15 & _T_1 ? $signed(32'sh0) : $signed(_GEN_204); // @[stackmanage_35.scala 879:71 stackmanage_35.scala 910:31]
  wire [31:0] _GEN_226 = LUT_stack_io_push_15 & _T_1 ? $signed(32'sh0) : $signed(_GEN_205); // @[stackmanage_35.scala 879:71 stackmanage_35.scala 911:31]
  wire [31:0] _GEN_227 = LUT_stack_io_push_15 & _T_1 ? $signed(32'sh0) : $signed(_GEN_206); // @[stackmanage_35.scala 879:71 stackmanage_35.scala 912:31]
  wire [31:0] _GEN_228 = LUT_stack_io_push_15 & _T_1 ? $signed(32'sh0) : $signed(_GEN_207); // @[stackmanage_35.scala 879:71 stackmanage_35.scala 913:31]
  wire [31:0] _GEN_229 = LUT_stack_io_push_15 & _T_1 ? $signed(32'sh0) : $signed(_GEN_208); // @[stackmanage_35.scala 879:71 stackmanage_35.scala 914:31]
  wire [31:0] _GEN_230 = LUT_stack_io_push_14 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 843:71 stackmanage_35.scala 844:30]
  wire [31:0] _GEN_232 = LUT_stack_io_push_14 & _T_1 ? $signed(32'sh0) : $signed(_GEN_209); // @[stackmanage_35.scala 843:71 stackmanage_35.scala 859:31]
  wire [31:0] _GEN_233 = LUT_stack_io_push_14 & _T_1 ? $signed(32'sh0) : $signed(_GEN_211); // @[stackmanage_35.scala 843:71 stackmanage_35.scala 860:31]
  wire [31:0] _GEN_234 = LUT_stack_io_push_14 & _T_1 ? $signed(32'sh0) : $signed(_GEN_212); // @[stackmanage_35.scala 843:71 stackmanage_35.scala 861:31]
  wire [31:0] _GEN_235 = LUT_stack_io_push_14 & _T_1 ? $signed(32'sh0) : $signed(_GEN_213); // @[stackmanage_35.scala 843:71 stackmanage_35.scala 862:31]
  wire [31:0] _GEN_236 = LUT_stack_io_push_14 & _T_1 ? $signed(32'sh0) : $signed(_GEN_214); // @[stackmanage_35.scala 843:71 stackmanage_35.scala 863:31]
  wire [31:0] _GEN_237 = LUT_stack_io_push_14 & _T_1 ? $signed(32'sh0) : $signed(_GEN_215); // @[stackmanage_35.scala 843:71 stackmanage_35.scala 864:31]
  wire [31:0] _GEN_238 = LUT_stack_io_push_14 & _T_1 ? $signed(32'sh0) : $signed(_GEN_216); // @[stackmanage_35.scala 843:71 stackmanage_35.scala 865:31]
  wire [31:0] _GEN_239 = LUT_stack_io_push_14 & _T_1 ? $signed(32'sh0) : $signed(_GEN_217); // @[stackmanage_35.scala 843:71 stackmanage_35.scala 866:31]
  wire [31:0] _GEN_240 = LUT_stack_io_push_14 & _T_1 ? $signed(32'sh0) : $signed(_GEN_218); // @[stackmanage_35.scala 843:71 stackmanage_35.scala 867:31]
  wire [31:0] _GEN_241 = LUT_stack_io_push_14 & _T_1 ? $signed(32'sh0) : $signed(_GEN_219); // @[stackmanage_35.scala 843:71 stackmanage_35.scala 868:31]
  wire [31:0] _GEN_242 = LUT_stack_io_push_14 & _T_1 ? $signed(32'sh0) : $signed(_GEN_220); // @[stackmanage_35.scala 843:71 stackmanage_35.scala 869:31]
  wire [31:0] _GEN_243 = LUT_stack_io_push_14 & _T_1 ? $signed(32'sh0) : $signed(_GEN_221); // @[stackmanage_35.scala 843:71 stackmanage_35.scala 870:31]
  wire [31:0] _GEN_244 = LUT_stack_io_push_14 & _T_1 ? $signed(32'sh0) : $signed(_GEN_222); // @[stackmanage_35.scala 843:71 stackmanage_35.scala 871:31]
  wire [31:0] _GEN_245 = LUT_stack_io_push_14 & _T_1 ? $signed(32'sh0) : $signed(_GEN_223); // @[stackmanage_35.scala 843:71 stackmanage_35.scala 872:31]
  wire [31:0] _GEN_246 = LUT_stack_io_push_14 & _T_1 ? $signed(32'sh0) : $signed(_GEN_224); // @[stackmanage_35.scala 843:71 stackmanage_35.scala 873:31]
  wire [31:0] _GEN_247 = LUT_stack_io_push_14 & _T_1 ? $signed(32'sh0) : $signed(_GEN_225); // @[stackmanage_35.scala 843:71 stackmanage_35.scala 874:31]
  wire [31:0] _GEN_248 = LUT_stack_io_push_14 & _T_1 ? $signed(32'sh0) : $signed(_GEN_226); // @[stackmanage_35.scala 843:71 stackmanage_35.scala 875:31]
  wire [31:0] _GEN_249 = LUT_stack_io_push_14 & _T_1 ? $signed(32'sh0) : $signed(_GEN_227); // @[stackmanage_35.scala 843:71 stackmanage_35.scala 876:31]
  wire [31:0] _GEN_250 = LUT_stack_io_push_14 & _T_1 ? $signed(32'sh0) : $signed(_GEN_228); // @[stackmanage_35.scala 843:71 stackmanage_35.scala 877:31]
  wire [31:0] _GEN_251 = LUT_stack_io_push_14 & _T_1 ? $signed(32'sh0) : $signed(_GEN_229); // @[stackmanage_35.scala 843:71 stackmanage_35.scala 878:31]
  wire [31:0] _GEN_252 = LUT_stack_io_push_13 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 807:71 stackmanage_35.scala 808:30]
  wire [31:0] _GEN_254 = LUT_stack_io_push_13 & _T_1 ? $signed(32'sh0) : $signed(_GEN_230); // @[stackmanage_35.scala 807:71 stackmanage_35.scala 822:31]
  wire [31:0] _GEN_255 = LUT_stack_io_push_13 & _T_1 ? $signed(32'sh0) : $signed(_GEN_232); // @[stackmanage_35.scala 807:71 stackmanage_35.scala 823:31]
  wire [31:0] _GEN_256 = LUT_stack_io_push_13 & _T_1 ? $signed(32'sh0) : $signed(_GEN_233); // @[stackmanage_35.scala 807:71 stackmanage_35.scala 824:31]
  wire [31:0] _GEN_257 = LUT_stack_io_push_13 & _T_1 ? $signed(32'sh0) : $signed(_GEN_234); // @[stackmanage_35.scala 807:71 stackmanage_35.scala 825:31]
  wire [31:0] _GEN_258 = LUT_stack_io_push_13 & _T_1 ? $signed(32'sh0) : $signed(_GEN_235); // @[stackmanage_35.scala 807:71 stackmanage_35.scala 826:31]
  wire [31:0] _GEN_259 = LUT_stack_io_push_13 & _T_1 ? $signed(32'sh0) : $signed(_GEN_236); // @[stackmanage_35.scala 807:71 stackmanage_35.scala 827:31]
  wire [31:0] _GEN_260 = LUT_stack_io_push_13 & _T_1 ? $signed(32'sh0) : $signed(_GEN_237); // @[stackmanage_35.scala 807:71 stackmanage_35.scala 828:31]
  wire [31:0] _GEN_261 = LUT_stack_io_push_13 & _T_1 ? $signed(32'sh0) : $signed(_GEN_238); // @[stackmanage_35.scala 807:71 stackmanage_35.scala 829:31]
  wire [31:0] _GEN_262 = LUT_stack_io_push_13 & _T_1 ? $signed(32'sh0) : $signed(_GEN_239); // @[stackmanage_35.scala 807:71 stackmanage_35.scala 830:31]
  wire [31:0] _GEN_263 = LUT_stack_io_push_13 & _T_1 ? $signed(32'sh0) : $signed(_GEN_240); // @[stackmanage_35.scala 807:71 stackmanage_35.scala 831:31]
  wire [31:0] _GEN_264 = LUT_stack_io_push_13 & _T_1 ? $signed(32'sh0) : $signed(_GEN_241); // @[stackmanage_35.scala 807:71 stackmanage_35.scala 832:31]
  wire [31:0] _GEN_265 = LUT_stack_io_push_13 & _T_1 ? $signed(32'sh0) : $signed(_GEN_242); // @[stackmanage_35.scala 807:71 stackmanage_35.scala 833:31]
  wire [31:0] _GEN_266 = LUT_stack_io_push_13 & _T_1 ? $signed(32'sh0) : $signed(_GEN_243); // @[stackmanage_35.scala 807:71 stackmanage_35.scala 834:31]
  wire [31:0] _GEN_267 = LUT_stack_io_push_13 & _T_1 ? $signed(32'sh0) : $signed(_GEN_244); // @[stackmanage_35.scala 807:71 stackmanage_35.scala 835:31]
  wire [31:0] _GEN_268 = LUT_stack_io_push_13 & _T_1 ? $signed(32'sh0) : $signed(_GEN_245); // @[stackmanage_35.scala 807:71 stackmanage_35.scala 836:31]
  wire [31:0] _GEN_269 = LUT_stack_io_push_13 & _T_1 ? $signed(32'sh0) : $signed(_GEN_246); // @[stackmanage_35.scala 807:71 stackmanage_35.scala 837:31]
  wire [31:0] _GEN_270 = LUT_stack_io_push_13 & _T_1 ? $signed(32'sh0) : $signed(_GEN_247); // @[stackmanage_35.scala 807:71 stackmanage_35.scala 838:31]
  wire [31:0] _GEN_271 = LUT_stack_io_push_13 & _T_1 ? $signed(32'sh0) : $signed(_GEN_248); // @[stackmanage_35.scala 807:71 stackmanage_35.scala 839:31]
  wire [31:0] _GEN_272 = LUT_stack_io_push_13 & _T_1 ? $signed(32'sh0) : $signed(_GEN_249); // @[stackmanage_35.scala 807:71 stackmanage_35.scala 840:31]
  wire [31:0] _GEN_273 = LUT_stack_io_push_13 & _T_1 ? $signed(32'sh0) : $signed(_GEN_250); // @[stackmanage_35.scala 807:71 stackmanage_35.scala 841:31]
  wire [31:0] _GEN_274 = LUT_stack_io_push_13 & _T_1 ? $signed(32'sh0) : $signed(_GEN_251); // @[stackmanage_35.scala 807:71 stackmanage_35.scala 842:31]
  wire [31:0] _GEN_275 = LUT_stack_io_push_12 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 771:71 stackmanage_35.scala 772:30]
  wire [31:0] _GEN_277 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_252); // @[stackmanage_35.scala 771:71 stackmanage_35.scala 785:31]
  wire [31:0] _GEN_278 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_254); // @[stackmanage_35.scala 771:71 stackmanage_35.scala 786:31]
  wire [31:0] _GEN_279 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_255); // @[stackmanage_35.scala 771:71 stackmanage_35.scala 787:31]
  wire [31:0] _GEN_280 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_256); // @[stackmanage_35.scala 771:71 stackmanage_35.scala 788:31]
  wire [31:0] _GEN_281 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_257); // @[stackmanage_35.scala 771:71 stackmanage_35.scala 789:31]
  wire [31:0] _GEN_282 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_258); // @[stackmanage_35.scala 771:71 stackmanage_35.scala 790:31]
  wire [31:0] _GEN_283 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_259); // @[stackmanage_35.scala 771:71 stackmanage_35.scala 791:31]
  wire [31:0] _GEN_284 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_260); // @[stackmanage_35.scala 771:71 stackmanage_35.scala 792:31]
  wire [31:0] _GEN_285 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_261); // @[stackmanage_35.scala 771:71 stackmanage_35.scala 793:31]
  wire [31:0] _GEN_286 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_262); // @[stackmanage_35.scala 771:71 stackmanage_35.scala 794:31]
  wire [31:0] _GEN_287 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_263); // @[stackmanage_35.scala 771:71 stackmanage_35.scala 795:31]
  wire [31:0] _GEN_288 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_264); // @[stackmanage_35.scala 771:71 stackmanage_35.scala 796:31]
  wire [31:0] _GEN_289 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_265); // @[stackmanage_35.scala 771:71 stackmanage_35.scala 797:31]
  wire [31:0] _GEN_290 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_266); // @[stackmanage_35.scala 771:71 stackmanage_35.scala 798:31]
  wire [31:0] _GEN_291 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_267); // @[stackmanage_35.scala 771:71 stackmanage_35.scala 799:31]
  wire [31:0] _GEN_292 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_268); // @[stackmanage_35.scala 771:71 stackmanage_35.scala 800:31]
  wire [31:0] _GEN_293 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_269); // @[stackmanage_35.scala 771:71 stackmanage_35.scala 801:31]
  wire [31:0] _GEN_294 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_270); // @[stackmanage_35.scala 771:71 stackmanage_35.scala 802:31]
  wire [31:0] _GEN_295 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_271); // @[stackmanage_35.scala 771:71 stackmanage_35.scala 803:31]
  wire [31:0] _GEN_296 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_272); // @[stackmanage_35.scala 771:71 stackmanage_35.scala 804:31]
  wire [31:0] _GEN_297 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_273); // @[stackmanage_35.scala 771:71 stackmanage_35.scala 805:31]
  wire [31:0] _GEN_298 = LUT_stack_io_push_12 & _T_1 ? $signed(32'sh0) : $signed(_GEN_274); // @[stackmanage_35.scala 771:71 stackmanage_35.scala 806:31]
  wire [31:0] _GEN_299 = LUT_stack_io_push_11 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 735:71 stackmanage_35.scala 736:30]
  wire [31:0] _GEN_301 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_275); // @[stackmanage_35.scala 735:71 stackmanage_35.scala 748:31]
  wire [31:0] _GEN_302 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_277); // @[stackmanage_35.scala 735:71 stackmanage_35.scala 749:31]
  wire [31:0] _GEN_303 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_278); // @[stackmanage_35.scala 735:71 stackmanage_35.scala 750:31]
  wire [31:0] _GEN_304 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_279); // @[stackmanage_35.scala 735:71 stackmanage_35.scala 751:31]
  wire [31:0] _GEN_305 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_280); // @[stackmanage_35.scala 735:71 stackmanage_35.scala 752:31]
  wire [31:0] _GEN_306 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_281); // @[stackmanage_35.scala 735:71 stackmanage_35.scala 753:31]
  wire [31:0] _GEN_307 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_282); // @[stackmanage_35.scala 735:71 stackmanage_35.scala 754:31]
  wire [31:0] _GEN_308 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_283); // @[stackmanage_35.scala 735:71 stackmanage_35.scala 755:31]
  wire [31:0] _GEN_309 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_284); // @[stackmanage_35.scala 735:71 stackmanage_35.scala 756:31]
  wire [31:0] _GEN_310 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_285); // @[stackmanage_35.scala 735:71 stackmanage_35.scala 757:31]
  wire [31:0] _GEN_311 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_286); // @[stackmanage_35.scala 735:71 stackmanage_35.scala 758:31]
  wire [31:0] _GEN_312 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_287); // @[stackmanage_35.scala 735:71 stackmanage_35.scala 759:31]
  wire [31:0] _GEN_313 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_288); // @[stackmanage_35.scala 735:71 stackmanage_35.scala 760:31]
  wire [31:0] _GEN_314 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_289); // @[stackmanage_35.scala 735:71 stackmanage_35.scala 761:31]
  wire [31:0] _GEN_315 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_290); // @[stackmanage_35.scala 735:71 stackmanage_35.scala 762:31]
  wire [31:0] _GEN_316 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_291); // @[stackmanage_35.scala 735:71 stackmanage_35.scala 763:31]
  wire [31:0] _GEN_317 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_292); // @[stackmanage_35.scala 735:71 stackmanage_35.scala 764:31]
  wire [31:0] _GEN_318 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_293); // @[stackmanage_35.scala 735:71 stackmanage_35.scala 765:31]
  wire [31:0] _GEN_319 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_294); // @[stackmanage_35.scala 735:71 stackmanage_35.scala 766:31]
  wire [31:0] _GEN_320 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_295); // @[stackmanage_35.scala 735:71 stackmanage_35.scala 767:31]
  wire [31:0] _GEN_321 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_296); // @[stackmanage_35.scala 735:71 stackmanage_35.scala 768:31]
  wire [31:0] _GEN_322 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_297); // @[stackmanage_35.scala 735:71 stackmanage_35.scala 769:31]
  wire [31:0] _GEN_323 = LUT_stack_io_push_11 & _T_1 ? $signed(32'sh0) : $signed(_GEN_298); // @[stackmanage_35.scala 735:71 stackmanage_35.scala 770:31]
  wire [31:0] _GEN_324 = LUT_stack_io_push_10 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 699:71 stackmanage_35.scala 700:30]
  wire [31:0] _GEN_326 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_299); // @[stackmanage_35.scala 699:71 stackmanage_35.scala 711:31]
  wire [31:0] _GEN_327 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_301); // @[stackmanage_35.scala 699:71 stackmanage_35.scala 712:31]
  wire [31:0] _GEN_328 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_302); // @[stackmanage_35.scala 699:71 stackmanage_35.scala 713:31]
  wire [31:0] _GEN_329 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_303); // @[stackmanage_35.scala 699:71 stackmanage_35.scala 714:31]
  wire [31:0] _GEN_330 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_304); // @[stackmanage_35.scala 699:71 stackmanage_35.scala 715:31]
  wire [31:0] _GEN_331 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_305); // @[stackmanage_35.scala 699:71 stackmanage_35.scala 716:31]
  wire [31:0] _GEN_332 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_306); // @[stackmanage_35.scala 699:71 stackmanage_35.scala 717:31]
  wire [31:0] _GEN_333 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_307); // @[stackmanage_35.scala 699:71 stackmanage_35.scala 718:31]
  wire [31:0] _GEN_334 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_308); // @[stackmanage_35.scala 699:71 stackmanage_35.scala 719:31]
  wire [31:0] _GEN_335 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_309); // @[stackmanage_35.scala 699:71 stackmanage_35.scala 720:31]
  wire [31:0] _GEN_336 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_310); // @[stackmanage_35.scala 699:71 stackmanage_35.scala 721:31]
  wire [31:0] _GEN_337 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_311); // @[stackmanage_35.scala 699:71 stackmanage_35.scala 722:31]
  wire [31:0] _GEN_338 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_312); // @[stackmanage_35.scala 699:71 stackmanage_35.scala 723:31]
  wire [31:0] _GEN_339 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_313); // @[stackmanage_35.scala 699:71 stackmanage_35.scala 724:31]
  wire [31:0] _GEN_340 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_314); // @[stackmanage_35.scala 699:71 stackmanage_35.scala 725:31]
  wire [31:0] _GEN_341 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_315); // @[stackmanage_35.scala 699:71 stackmanage_35.scala 726:31]
  wire [31:0] _GEN_342 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_316); // @[stackmanage_35.scala 699:71 stackmanage_35.scala 727:31]
  wire [31:0] _GEN_343 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_317); // @[stackmanage_35.scala 699:71 stackmanage_35.scala 728:31]
  wire [31:0] _GEN_344 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_318); // @[stackmanage_35.scala 699:71 stackmanage_35.scala 729:31]
  wire [31:0] _GEN_345 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_319); // @[stackmanage_35.scala 699:71 stackmanage_35.scala 730:31]
  wire [31:0] _GEN_346 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_320); // @[stackmanage_35.scala 699:71 stackmanage_35.scala 731:31]
  wire [31:0] _GEN_347 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_321); // @[stackmanage_35.scala 699:71 stackmanage_35.scala 732:31]
  wire [31:0] _GEN_348 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_322); // @[stackmanage_35.scala 699:71 stackmanage_35.scala 733:31]
  wire [31:0] _GEN_349 = LUT_stack_io_push_10 & _T_1 ? $signed(32'sh0) : $signed(_GEN_323); // @[stackmanage_35.scala 699:71 stackmanage_35.scala 734:31]
  wire [31:0] _GEN_350 = LUT_stack_io_push_9 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 663:70 stackmanage_35.scala 664:29]
  wire [31:0] _GEN_352 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_324); // @[stackmanage_35.scala 663:70 stackmanage_35.scala 674:31]
  wire [31:0] _GEN_353 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_326); // @[stackmanage_35.scala 663:70 stackmanage_35.scala 675:31]
  wire [31:0] _GEN_354 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_327); // @[stackmanage_35.scala 663:70 stackmanage_35.scala 676:31]
  wire [31:0] _GEN_355 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_328); // @[stackmanage_35.scala 663:70 stackmanage_35.scala 677:31]
  wire [31:0] _GEN_356 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_329); // @[stackmanage_35.scala 663:70 stackmanage_35.scala 678:31]
  wire [31:0] _GEN_357 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_330); // @[stackmanage_35.scala 663:70 stackmanage_35.scala 679:31]
  wire [31:0] _GEN_358 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_331); // @[stackmanage_35.scala 663:70 stackmanage_35.scala 680:31]
  wire [31:0] _GEN_359 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_332); // @[stackmanage_35.scala 663:70 stackmanage_35.scala 681:31]
  wire [31:0] _GEN_360 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_333); // @[stackmanage_35.scala 663:70 stackmanage_35.scala 682:31]
  wire [31:0] _GEN_361 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_334); // @[stackmanage_35.scala 663:70 stackmanage_35.scala 683:31]
  wire [31:0] _GEN_362 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_335); // @[stackmanage_35.scala 663:70 stackmanage_35.scala 684:31]
  wire [31:0] _GEN_363 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_336); // @[stackmanage_35.scala 663:70 stackmanage_35.scala 685:31]
  wire [31:0] _GEN_364 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_337); // @[stackmanage_35.scala 663:70 stackmanage_35.scala 686:31]
  wire [31:0] _GEN_365 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_338); // @[stackmanage_35.scala 663:70 stackmanage_35.scala 687:31]
  wire [31:0] _GEN_366 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_339); // @[stackmanage_35.scala 663:70 stackmanage_35.scala 688:31]
  wire [31:0] _GEN_367 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_340); // @[stackmanage_35.scala 663:70 stackmanage_35.scala 689:31]
  wire [31:0] _GEN_368 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_341); // @[stackmanage_35.scala 663:70 stackmanage_35.scala 690:31]
  wire [31:0] _GEN_369 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_342); // @[stackmanage_35.scala 663:70 stackmanage_35.scala 691:31]
  wire [31:0] _GEN_370 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_343); // @[stackmanage_35.scala 663:70 stackmanage_35.scala 692:31]
  wire [31:0] _GEN_371 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_344); // @[stackmanage_35.scala 663:70 stackmanage_35.scala 693:31]
  wire [31:0] _GEN_372 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_345); // @[stackmanage_35.scala 663:70 stackmanage_35.scala 694:31]
  wire [31:0] _GEN_373 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_346); // @[stackmanage_35.scala 663:70 stackmanage_35.scala 695:31]
  wire [31:0] _GEN_374 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_347); // @[stackmanage_35.scala 663:70 stackmanage_35.scala 696:31]
  wire [31:0] _GEN_375 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_348); // @[stackmanage_35.scala 663:70 stackmanage_35.scala 697:31]
  wire [31:0] _GEN_376 = LUT_stack_io_push_9 & _T_1 ? $signed(32'sh0) : $signed(_GEN_349); // @[stackmanage_35.scala 663:70 stackmanage_35.scala 698:31]
  wire [31:0] _GEN_377 = LUT_stack_io_push_8 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 627:70 stackmanage_35.scala 628:29]
  wire [31:0] _GEN_379 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_350); // @[stackmanage_35.scala 627:70 stackmanage_35.scala 637:30]
  wire [31:0] _GEN_380 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_352); // @[stackmanage_35.scala 627:70 stackmanage_35.scala 638:31]
  wire [31:0] _GEN_381 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_353); // @[stackmanage_35.scala 627:70 stackmanage_35.scala 639:31]
  wire [31:0] _GEN_382 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_354); // @[stackmanage_35.scala 627:70 stackmanage_35.scala 640:31]
  wire [31:0] _GEN_383 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_355); // @[stackmanage_35.scala 627:70 stackmanage_35.scala 641:31]
  wire [31:0] _GEN_384 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_356); // @[stackmanage_35.scala 627:70 stackmanage_35.scala 642:31]
  wire [31:0] _GEN_385 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_357); // @[stackmanage_35.scala 627:70 stackmanage_35.scala 643:31]
  wire [31:0] _GEN_386 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_358); // @[stackmanage_35.scala 627:70 stackmanage_35.scala 644:31]
  wire [31:0] _GEN_387 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_359); // @[stackmanage_35.scala 627:70 stackmanage_35.scala 645:31]
  wire [31:0] _GEN_388 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_360); // @[stackmanage_35.scala 627:70 stackmanage_35.scala 646:31]
  wire [31:0] _GEN_389 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_361); // @[stackmanage_35.scala 627:70 stackmanage_35.scala 647:31]
  wire [31:0] _GEN_390 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_362); // @[stackmanage_35.scala 627:70 stackmanage_35.scala 648:31]
  wire [31:0] _GEN_391 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_363); // @[stackmanage_35.scala 627:70 stackmanage_35.scala 649:31]
  wire [31:0] _GEN_392 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_364); // @[stackmanage_35.scala 627:70 stackmanage_35.scala 650:31]
  wire [31:0] _GEN_393 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_365); // @[stackmanage_35.scala 627:70 stackmanage_35.scala 651:31]
  wire [31:0] _GEN_394 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_366); // @[stackmanage_35.scala 627:70 stackmanage_35.scala 652:31]
  wire [31:0] _GEN_395 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_367); // @[stackmanage_35.scala 627:70 stackmanage_35.scala 653:31]
  wire [31:0] _GEN_396 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_368); // @[stackmanage_35.scala 627:70 stackmanage_35.scala 654:31]
  wire [31:0] _GEN_397 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_369); // @[stackmanage_35.scala 627:70 stackmanage_35.scala 655:31]
  wire [31:0] _GEN_398 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_370); // @[stackmanage_35.scala 627:70 stackmanage_35.scala 656:31]
  wire [31:0] _GEN_399 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_371); // @[stackmanage_35.scala 627:70 stackmanage_35.scala 657:31]
  wire [31:0] _GEN_400 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_372); // @[stackmanage_35.scala 627:70 stackmanage_35.scala 658:31]
  wire [31:0] _GEN_401 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_373); // @[stackmanage_35.scala 627:70 stackmanage_35.scala 659:31]
  wire [31:0] _GEN_402 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_374); // @[stackmanage_35.scala 627:70 stackmanage_35.scala 660:31]
  wire [31:0] _GEN_403 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_375); // @[stackmanage_35.scala 627:70 stackmanage_35.scala 661:31]
  wire [31:0] _GEN_404 = LUT_stack_io_push_8 & _T_1 ? $signed(32'sh0) : $signed(_GEN_376); // @[stackmanage_35.scala 627:70 stackmanage_35.scala 662:31]
  wire [31:0] _GEN_405 = LUT_stack_io_push_7 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 591:70 stackmanage_35.scala 592:29]
  wire [31:0] _GEN_407 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_377); // @[stackmanage_35.scala 591:70 stackmanage_35.scala 600:30]
  wire [31:0] _GEN_408 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_379); // @[stackmanage_35.scala 591:70 stackmanage_35.scala 601:30]
  wire [31:0] _GEN_409 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_380); // @[stackmanage_35.scala 591:70 stackmanage_35.scala 602:31]
  wire [31:0] _GEN_410 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_381); // @[stackmanage_35.scala 591:70 stackmanage_35.scala 603:31]
  wire [31:0] _GEN_411 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_382); // @[stackmanage_35.scala 591:70 stackmanage_35.scala 604:31]
  wire [31:0] _GEN_412 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_383); // @[stackmanage_35.scala 591:70 stackmanage_35.scala 605:31]
  wire [31:0] _GEN_413 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_384); // @[stackmanage_35.scala 591:70 stackmanage_35.scala 606:31]
  wire [31:0] _GEN_414 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_385); // @[stackmanage_35.scala 591:70 stackmanage_35.scala 607:31]
  wire [31:0] _GEN_415 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_386); // @[stackmanage_35.scala 591:70 stackmanage_35.scala 608:31]
  wire [31:0] _GEN_416 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_387); // @[stackmanage_35.scala 591:70 stackmanage_35.scala 609:31]
  wire [31:0] _GEN_417 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_388); // @[stackmanage_35.scala 591:70 stackmanage_35.scala 610:31]
  wire [31:0] _GEN_418 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_389); // @[stackmanage_35.scala 591:70 stackmanage_35.scala 611:31]
  wire [31:0] _GEN_419 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_390); // @[stackmanage_35.scala 591:70 stackmanage_35.scala 612:31]
  wire [31:0] _GEN_420 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_391); // @[stackmanage_35.scala 591:70 stackmanage_35.scala 613:31]
  wire [31:0] _GEN_421 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_392); // @[stackmanage_35.scala 591:70 stackmanage_35.scala 614:31]
  wire [31:0] _GEN_422 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_393); // @[stackmanage_35.scala 591:70 stackmanage_35.scala 615:31]
  wire [31:0] _GEN_423 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_394); // @[stackmanage_35.scala 591:70 stackmanage_35.scala 616:31]
  wire [31:0] _GEN_424 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_395); // @[stackmanage_35.scala 591:70 stackmanage_35.scala 617:31]
  wire [31:0] _GEN_425 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_396); // @[stackmanage_35.scala 591:70 stackmanage_35.scala 618:31]
  wire [31:0] _GEN_426 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_397); // @[stackmanage_35.scala 591:70 stackmanage_35.scala 619:31]
  wire [31:0] _GEN_427 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_398); // @[stackmanage_35.scala 591:70 stackmanage_35.scala 620:31]
  wire [31:0] _GEN_428 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_399); // @[stackmanage_35.scala 591:70 stackmanage_35.scala 621:31]
  wire [31:0] _GEN_429 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_400); // @[stackmanage_35.scala 591:70 stackmanage_35.scala 622:31]
  wire [31:0] _GEN_430 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_401); // @[stackmanage_35.scala 591:70 stackmanage_35.scala 623:31]
  wire [31:0] _GEN_431 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_402); // @[stackmanage_35.scala 591:70 stackmanage_35.scala 624:31]
  wire [31:0] _GEN_432 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_403); // @[stackmanage_35.scala 591:70 stackmanage_35.scala 625:31]
  wire [31:0] _GEN_433 = LUT_stack_io_push_7 & _T_1 ? $signed(32'sh0) : $signed(_GEN_404); // @[stackmanage_35.scala 591:70 stackmanage_35.scala 626:31]
  wire [31:0] _GEN_434 = LUT_stack_io_push_6 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 555:70 stackmanage_35.scala 556:29]
  wire [31:0] _GEN_436 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_405); // @[stackmanage_35.scala 555:70 stackmanage_35.scala 563:30]
  wire [31:0] _GEN_437 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_407); // @[stackmanage_35.scala 555:70 stackmanage_35.scala 564:30]
  wire [31:0] _GEN_438 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_408); // @[stackmanage_35.scala 555:70 stackmanage_35.scala 565:30]
  wire [31:0] _GEN_439 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_409); // @[stackmanage_35.scala 555:70 stackmanage_35.scala 566:31]
  wire [31:0] _GEN_440 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_410); // @[stackmanage_35.scala 555:70 stackmanage_35.scala 567:31]
  wire [31:0] _GEN_441 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_411); // @[stackmanage_35.scala 555:70 stackmanage_35.scala 568:31]
  wire [31:0] _GEN_442 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_412); // @[stackmanage_35.scala 555:70 stackmanage_35.scala 569:31]
  wire [31:0] _GEN_443 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_413); // @[stackmanage_35.scala 555:70 stackmanage_35.scala 570:31]
  wire [31:0] _GEN_444 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_414); // @[stackmanage_35.scala 555:70 stackmanage_35.scala 571:31]
  wire [31:0] _GEN_445 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_415); // @[stackmanage_35.scala 555:70 stackmanage_35.scala 572:31]
  wire [31:0] _GEN_446 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_416); // @[stackmanage_35.scala 555:70 stackmanage_35.scala 573:31]
  wire [31:0] _GEN_447 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_417); // @[stackmanage_35.scala 555:70 stackmanage_35.scala 574:31]
  wire [31:0] _GEN_448 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_418); // @[stackmanage_35.scala 555:70 stackmanage_35.scala 575:31]
  wire [31:0] _GEN_449 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_419); // @[stackmanage_35.scala 555:70 stackmanage_35.scala 576:31]
  wire [31:0] _GEN_450 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_420); // @[stackmanage_35.scala 555:70 stackmanage_35.scala 577:31]
  wire [31:0] _GEN_451 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_421); // @[stackmanage_35.scala 555:70 stackmanage_35.scala 578:31]
  wire [31:0] _GEN_452 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_422); // @[stackmanage_35.scala 555:70 stackmanage_35.scala 579:31]
  wire [31:0] _GEN_453 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_423); // @[stackmanage_35.scala 555:70 stackmanage_35.scala 580:31]
  wire [31:0] _GEN_454 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_424); // @[stackmanage_35.scala 555:70 stackmanage_35.scala 581:31]
  wire [31:0] _GEN_455 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_425); // @[stackmanage_35.scala 555:70 stackmanage_35.scala 582:31]
  wire [31:0] _GEN_456 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_426); // @[stackmanage_35.scala 555:70 stackmanage_35.scala 583:31]
  wire [31:0] _GEN_457 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_427); // @[stackmanage_35.scala 555:70 stackmanage_35.scala 584:31]
  wire [31:0] _GEN_458 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_428); // @[stackmanage_35.scala 555:70 stackmanage_35.scala 585:31]
  wire [31:0] _GEN_459 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_429); // @[stackmanage_35.scala 555:70 stackmanage_35.scala 586:31]
  wire [31:0] _GEN_460 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_430); // @[stackmanage_35.scala 555:70 stackmanage_35.scala 587:31]
  wire [31:0] _GEN_461 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_431); // @[stackmanage_35.scala 555:70 stackmanage_35.scala 588:31]
  wire [31:0] _GEN_462 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_432); // @[stackmanage_35.scala 555:70 stackmanage_35.scala 589:31]
  wire [31:0] _GEN_463 = LUT_stack_io_push_6 & _T_1 ? $signed(32'sh0) : $signed(_GEN_433); // @[stackmanage_35.scala 555:70 stackmanage_35.scala 590:31]
  wire [31:0] _GEN_464 = LUT_stack_io_push_5 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 519:70 stackmanage_35.scala 520:29]
  wire [31:0] _GEN_466 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_434); // @[stackmanage_35.scala 519:70 stackmanage_35.scala 526:30]
  wire [31:0] _GEN_467 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_436); // @[stackmanage_35.scala 519:70 stackmanage_35.scala 527:30]
  wire [31:0] _GEN_468 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_437); // @[stackmanage_35.scala 519:70 stackmanage_35.scala 528:30]
  wire [31:0] _GEN_469 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_438); // @[stackmanage_35.scala 519:70 stackmanage_35.scala 529:30]
  wire [31:0] _GEN_470 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_439); // @[stackmanage_35.scala 519:70 stackmanage_35.scala 530:31]
  wire [31:0] _GEN_471 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_440); // @[stackmanage_35.scala 519:70 stackmanage_35.scala 531:31]
  wire [31:0] _GEN_472 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_441); // @[stackmanage_35.scala 519:70 stackmanage_35.scala 532:31]
  wire [31:0] _GEN_473 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_442); // @[stackmanage_35.scala 519:70 stackmanage_35.scala 533:31]
  wire [31:0] _GEN_474 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_443); // @[stackmanage_35.scala 519:70 stackmanage_35.scala 534:31]
  wire [31:0] _GEN_475 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_444); // @[stackmanage_35.scala 519:70 stackmanage_35.scala 535:31]
  wire [31:0] _GEN_476 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_445); // @[stackmanage_35.scala 519:70 stackmanage_35.scala 536:31]
  wire [31:0] _GEN_477 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_446); // @[stackmanage_35.scala 519:70 stackmanage_35.scala 537:31]
  wire [31:0] _GEN_478 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_447); // @[stackmanage_35.scala 519:70 stackmanage_35.scala 538:31]
  wire [31:0] _GEN_479 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_448); // @[stackmanage_35.scala 519:70 stackmanage_35.scala 539:31]
  wire [31:0] _GEN_480 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_449); // @[stackmanage_35.scala 519:70 stackmanage_35.scala 540:31]
  wire [31:0] _GEN_481 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_450); // @[stackmanage_35.scala 519:70 stackmanage_35.scala 541:31]
  wire [31:0] _GEN_482 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_451); // @[stackmanage_35.scala 519:70 stackmanage_35.scala 542:31]
  wire [31:0] _GEN_483 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_452); // @[stackmanage_35.scala 519:70 stackmanage_35.scala 543:31]
  wire [31:0] _GEN_484 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_453); // @[stackmanage_35.scala 519:70 stackmanage_35.scala 544:31]
  wire [31:0] _GEN_485 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_454); // @[stackmanage_35.scala 519:70 stackmanage_35.scala 545:31]
  wire [31:0] _GEN_486 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_455); // @[stackmanage_35.scala 519:70 stackmanage_35.scala 546:31]
  wire [31:0] _GEN_487 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_456); // @[stackmanage_35.scala 519:70 stackmanage_35.scala 547:31]
  wire [31:0] _GEN_488 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_457); // @[stackmanage_35.scala 519:70 stackmanage_35.scala 548:31]
  wire [31:0] _GEN_489 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_458); // @[stackmanage_35.scala 519:70 stackmanage_35.scala 549:31]
  wire [31:0] _GEN_490 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_459); // @[stackmanage_35.scala 519:70 stackmanage_35.scala 550:31]
  wire [31:0] _GEN_491 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_460); // @[stackmanage_35.scala 519:70 stackmanage_35.scala 551:31]
  wire [31:0] _GEN_492 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_461); // @[stackmanage_35.scala 519:70 stackmanage_35.scala 552:31]
  wire [31:0] _GEN_493 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_462); // @[stackmanage_35.scala 519:70 stackmanage_35.scala 553:31]
  wire [31:0] _GEN_494 = LUT_stack_io_push_5 & _T_1 ? $signed(32'sh0) : $signed(_GEN_463); // @[stackmanage_35.scala 519:70 stackmanage_35.scala 554:31]
  wire [31:0] _GEN_495 = LUT_stack_io_push_4 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 483:70 stackmanage_35.scala 484:29]
  wire [31:0] _GEN_497 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_464); // @[stackmanage_35.scala 483:70 stackmanage_35.scala 489:30]
  wire [31:0] _GEN_498 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_466); // @[stackmanage_35.scala 483:70 stackmanage_35.scala 490:30]
  wire [31:0] _GEN_499 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_467); // @[stackmanage_35.scala 483:70 stackmanage_35.scala 491:30]
  wire [31:0] _GEN_500 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_468); // @[stackmanage_35.scala 483:70 stackmanage_35.scala 492:30]
  wire [31:0] _GEN_501 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_469); // @[stackmanage_35.scala 483:70 stackmanage_35.scala 493:30]
  wire [31:0] _GEN_502 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_470); // @[stackmanage_35.scala 483:70 stackmanage_35.scala 494:31]
  wire [31:0] _GEN_503 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_471); // @[stackmanage_35.scala 483:70 stackmanage_35.scala 495:31]
  wire [31:0] _GEN_504 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_472); // @[stackmanage_35.scala 483:70 stackmanage_35.scala 496:31]
  wire [31:0] _GEN_505 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_473); // @[stackmanage_35.scala 483:70 stackmanage_35.scala 497:31]
  wire [31:0] _GEN_506 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_474); // @[stackmanage_35.scala 483:70 stackmanage_35.scala 498:31]
  wire [31:0] _GEN_507 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_475); // @[stackmanage_35.scala 483:70 stackmanage_35.scala 499:31]
  wire [31:0] _GEN_508 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_476); // @[stackmanage_35.scala 483:70 stackmanage_35.scala 500:31]
  wire [31:0] _GEN_509 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_477); // @[stackmanage_35.scala 483:70 stackmanage_35.scala 501:31]
  wire [31:0] _GEN_510 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_478); // @[stackmanage_35.scala 483:70 stackmanage_35.scala 502:31]
  wire [31:0] _GEN_511 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_479); // @[stackmanage_35.scala 483:70 stackmanage_35.scala 503:31]
  wire [31:0] _GEN_512 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_480); // @[stackmanage_35.scala 483:70 stackmanage_35.scala 504:31]
  wire [31:0] _GEN_513 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_481); // @[stackmanage_35.scala 483:70 stackmanage_35.scala 505:31]
  wire [31:0] _GEN_514 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_482); // @[stackmanage_35.scala 483:70 stackmanage_35.scala 506:31]
  wire [31:0] _GEN_515 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_483); // @[stackmanage_35.scala 483:70 stackmanage_35.scala 507:31]
  wire [31:0] _GEN_516 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_484); // @[stackmanage_35.scala 483:70 stackmanage_35.scala 508:31]
  wire [31:0] _GEN_517 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_485); // @[stackmanage_35.scala 483:70 stackmanage_35.scala 509:31]
  wire [31:0] _GEN_518 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_486); // @[stackmanage_35.scala 483:70 stackmanage_35.scala 510:31]
  wire [31:0] _GEN_519 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_487); // @[stackmanage_35.scala 483:70 stackmanage_35.scala 511:31]
  wire [31:0] _GEN_520 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_488); // @[stackmanage_35.scala 483:70 stackmanage_35.scala 512:31]
  wire [31:0] _GEN_521 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_489); // @[stackmanage_35.scala 483:70 stackmanage_35.scala 513:31]
  wire [31:0] _GEN_522 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_490); // @[stackmanage_35.scala 483:70 stackmanage_35.scala 514:31]
  wire [31:0] _GEN_523 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_491); // @[stackmanage_35.scala 483:70 stackmanage_35.scala 515:31]
  wire [31:0] _GEN_524 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_492); // @[stackmanage_35.scala 483:70 stackmanage_35.scala 516:31]
  wire [31:0] _GEN_525 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_493); // @[stackmanage_35.scala 483:70 stackmanage_35.scala 517:31]
  wire [31:0] _GEN_526 = LUT_stack_io_push_4 & _T_1 ? $signed(32'sh0) : $signed(_GEN_494); // @[stackmanage_35.scala 483:70 stackmanage_35.scala 518:31]
  wire [31:0] _GEN_527 = LUT_stack_io_push_3 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 447:70 stackmanage_35.scala 448:29]
  wire [31:0] _GEN_529 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_495); // @[stackmanage_35.scala 447:70 stackmanage_35.scala 452:30]
  wire [31:0] _GEN_530 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_497); // @[stackmanage_35.scala 447:70 stackmanage_35.scala 453:30]
  wire [31:0] _GEN_531 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_498); // @[stackmanage_35.scala 447:70 stackmanage_35.scala 454:30]
  wire [31:0] _GEN_532 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_499); // @[stackmanage_35.scala 447:70 stackmanage_35.scala 455:30]
  wire [31:0] _GEN_533 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_500); // @[stackmanage_35.scala 447:70 stackmanage_35.scala 456:30]
  wire [31:0] _GEN_534 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_501); // @[stackmanage_35.scala 447:70 stackmanage_35.scala 457:30]
  wire [31:0] _GEN_535 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_502); // @[stackmanage_35.scala 447:70 stackmanage_35.scala 458:31]
  wire [31:0] _GEN_536 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_503); // @[stackmanage_35.scala 447:70 stackmanage_35.scala 459:31]
  wire [31:0] _GEN_537 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_504); // @[stackmanage_35.scala 447:70 stackmanage_35.scala 460:31]
  wire [31:0] _GEN_538 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_505); // @[stackmanage_35.scala 447:70 stackmanage_35.scala 461:31]
  wire [31:0] _GEN_539 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_506); // @[stackmanage_35.scala 447:70 stackmanage_35.scala 462:31]
  wire [31:0] _GEN_540 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_507); // @[stackmanage_35.scala 447:70 stackmanage_35.scala 463:31]
  wire [31:0] _GEN_541 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_508); // @[stackmanage_35.scala 447:70 stackmanage_35.scala 464:31]
  wire [31:0] _GEN_542 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_509); // @[stackmanage_35.scala 447:70 stackmanage_35.scala 465:31]
  wire [31:0] _GEN_543 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_510); // @[stackmanage_35.scala 447:70 stackmanage_35.scala 466:31]
  wire [31:0] _GEN_544 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_511); // @[stackmanage_35.scala 447:70 stackmanage_35.scala 467:31]
  wire [31:0] _GEN_545 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_512); // @[stackmanage_35.scala 447:70 stackmanage_35.scala 468:31]
  wire [31:0] _GEN_546 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_513); // @[stackmanage_35.scala 447:70 stackmanage_35.scala 469:31]
  wire [31:0] _GEN_547 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_514); // @[stackmanage_35.scala 447:70 stackmanage_35.scala 470:31]
  wire [31:0] _GEN_548 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_515); // @[stackmanage_35.scala 447:70 stackmanage_35.scala 471:31]
  wire [31:0] _GEN_549 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_516); // @[stackmanage_35.scala 447:70 stackmanage_35.scala 472:31]
  wire [31:0] _GEN_550 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_517); // @[stackmanage_35.scala 447:70 stackmanage_35.scala 473:31]
  wire [31:0] _GEN_551 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_518); // @[stackmanage_35.scala 447:70 stackmanage_35.scala 474:31]
  wire [31:0] _GEN_552 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_519); // @[stackmanage_35.scala 447:70 stackmanage_35.scala 475:31]
  wire [31:0] _GEN_553 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_520); // @[stackmanage_35.scala 447:70 stackmanage_35.scala 476:31]
  wire [31:0] _GEN_554 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_521); // @[stackmanage_35.scala 447:70 stackmanage_35.scala 477:31]
  wire [31:0] _GEN_555 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_522); // @[stackmanage_35.scala 447:70 stackmanage_35.scala 478:31]
  wire [31:0] _GEN_556 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_523); // @[stackmanage_35.scala 447:70 stackmanage_35.scala 479:31]
  wire [31:0] _GEN_557 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_524); // @[stackmanage_35.scala 447:70 stackmanage_35.scala 480:31]
  wire [31:0] _GEN_558 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_525); // @[stackmanage_35.scala 447:70 stackmanage_35.scala 481:31]
  wire [31:0] _GEN_559 = LUT_stack_io_push_3 & _T_1 ? $signed(32'sh0) : $signed(_GEN_526); // @[stackmanage_35.scala 447:70 stackmanage_35.scala 482:31]
  wire [31:0] _GEN_560 = LUT_stack_io_push_2 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 411:70 stackmanage_35.scala 412:29]
  wire [31:0] _GEN_562 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_527); // @[stackmanage_35.scala 411:70 stackmanage_35.scala 415:30]
  wire [31:0] _GEN_563 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_529); // @[stackmanage_35.scala 411:70 stackmanage_35.scala 416:30]
  wire [31:0] _GEN_564 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_530); // @[stackmanage_35.scala 411:70 stackmanage_35.scala 417:30]
  wire [31:0] _GEN_565 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_531); // @[stackmanage_35.scala 411:70 stackmanage_35.scala 418:30]
  wire [31:0] _GEN_566 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_532); // @[stackmanage_35.scala 411:70 stackmanage_35.scala 419:30]
  wire [31:0] _GEN_567 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_533); // @[stackmanage_35.scala 411:70 stackmanage_35.scala 420:30]
  wire [31:0] _GEN_568 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_534); // @[stackmanage_35.scala 411:70 stackmanage_35.scala 421:30]
  wire [31:0] _GEN_569 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_535); // @[stackmanage_35.scala 411:70 stackmanage_35.scala 422:31]
  wire [31:0] _GEN_570 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_536); // @[stackmanage_35.scala 411:70 stackmanage_35.scala 423:31]
  wire [31:0] _GEN_571 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_537); // @[stackmanage_35.scala 411:70 stackmanage_35.scala 424:31]
  wire [31:0] _GEN_572 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_538); // @[stackmanage_35.scala 411:70 stackmanage_35.scala 425:31]
  wire [31:0] _GEN_573 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_539); // @[stackmanage_35.scala 411:70 stackmanage_35.scala 426:31]
  wire [31:0] _GEN_574 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_540); // @[stackmanage_35.scala 411:70 stackmanage_35.scala 427:31]
  wire [31:0] _GEN_575 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_541); // @[stackmanage_35.scala 411:70 stackmanage_35.scala 428:31]
  wire [31:0] _GEN_576 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_542); // @[stackmanage_35.scala 411:70 stackmanage_35.scala 429:31]
  wire [31:0] _GEN_577 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_543); // @[stackmanage_35.scala 411:70 stackmanage_35.scala 430:31]
  wire [31:0] _GEN_578 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_544); // @[stackmanage_35.scala 411:70 stackmanage_35.scala 431:31]
  wire [31:0] _GEN_579 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_545); // @[stackmanage_35.scala 411:70 stackmanage_35.scala 432:31]
  wire [31:0] _GEN_580 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_546); // @[stackmanage_35.scala 411:70 stackmanage_35.scala 433:31]
  wire [31:0] _GEN_581 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_547); // @[stackmanage_35.scala 411:70 stackmanage_35.scala 434:31]
  wire [31:0] _GEN_582 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_548); // @[stackmanage_35.scala 411:70 stackmanage_35.scala 435:31]
  wire [31:0] _GEN_583 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_549); // @[stackmanage_35.scala 411:70 stackmanage_35.scala 436:31]
  wire [31:0] _GEN_584 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_550); // @[stackmanage_35.scala 411:70 stackmanage_35.scala 437:31]
  wire [31:0] _GEN_585 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_551); // @[stackmanage_35.scala 411:70 stackmanage_35.scala 438:31]
  wire [31:0] _GEN_586 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_552); // @[stackmanage_35.scala 411:70 stackmanage_35.scala 439:31]
  wire [31:0] _GEN_587 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_553); // @[stackmanage_35.scala 411:70 stackmanage_35.scala 440:31]
  wire [31:0] _GEN_588 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_554); // @[stackmanage_35.scala 411:70 stackmanage_35.scala 441:31]
  wire [31:0] _GEN_589 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_555); // @[stackmanage_35.scala 411:70 stackmanage_35.scala 442:31]
  wire [31:0] _GEN_590 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_556); // @[stackmanage_35.scala 411:70 stackmanage_35.scala 443:31]
  wire [31:0] _GEN_591 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_557); // @[stackmanage_35.scala 411:70 stackmanage_35.scala 444:31]
  wire [31:0] _GEN_592 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_558); // @[stackmanage_35.scala 411:70 stackmanage_35.scala 445:31]
  wire [31:0] _GEN_593 = LUT_stack_io_push_2 & _T_1 ? $signed(32'sh0) : $signed(_GEN_559); // @[stackmanage_35.scala 411:70 stackmanage_35.scala 446:31]
  wire [31:0] _GEN_594 = LUT_stack_io_push_1 & _T_1 ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 375:70 stackmanage_35.scala 376:29]
  wire [31:0] _GEN_596 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_560); // @[stackmanage_35.scala 375:70 stackmanage_35.scala 378:30]
  wire [31:0] _GEN_597 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_562); // @[stackmanage_35.scala 375:70 stackmanage_35.scala 379:30]
  wire [31:0] _GEN_598 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_563); // @[stackmanage_35.scala 375:70 stackmanage_35.scala 380:30]
  wire [31:0] _GEN_599 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_564); // @[stackmanage_35.scala 375:70 stackmanage_35.scala 381:30]
  wire [31:0] _GEN_600 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_565); // @[stackmanage_35.scala 375:70 stackmanage_35.scala 382:30]
  wire [31:0] _GEN_601 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_566); // @[stackmanage_35.scala 375:70 stackmanage_35.scala 383:30]
  wire [31:0] _GEN_602 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_567); // @[stackmanage_35.scala 375:70 stackmanage_35.scala 384:30]
  wire [31:0] _GEN_603 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_568); // @[stackmanage_35.scala 375:70 stackmanage_35.scala 385:30]
  wire [31:0] _GEN_604 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_569); // @[stackmanage_35.scala 375:70 stackmanage_35.scala 386:31]
  wire [31:0] _GEN_605 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_570); // @[stackmanage_35.scala 375:70 stackmanage_35.scala 387:31]
  wire [31:0] _GEN_606 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_571); // @[stackmanage_35.scala 375:70 stackmanage_35.scala 388:31]
  wire [31:0] _GEN_607 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_572); // @[stackmanage_35.scala 375:70 stackmanage_35.scala 389:31]
  wire [31:0] _GEN_608 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_573); // @[stackmanage_35.scala 375:70 stackmanage_35.scala 390:31]
  wire [31:0] _GEN_609 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_574); // @[stackmanage_35.scala 375:70 stackmanage_35.scala 391:31]
  wire [31:0] _GEN_610 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_575); // @[stackmanage_35.scala 375:70 stackmanage_35.scala 392:31]
  wire [31:0] _GEN_611 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_576); // @[stackmanage_35.scala 375:70 stackmanage_35.scala 393:31]
  wire [31:0] _GEN_612 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_577); // @[stackmanage_35.scala 375:70 stackmanage_35.scala 394:31]
  wire [31:0] _GEN_613 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_578); // @[stackmanage_35.scala 375:70 stackmanage_35.scala 395:31]
  wire [31:0] _GEN_614 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_579); // @[stackmanage_35.scala 375:70 stackmanage_35.scala 396:31]
  wire [31:0] _GEN_615 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_580); // @[stackmanage_35.scala 375:70 stackmanage_35.scala 397:31]
  wire [31:0] _GEN_616 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_581); // @[stackmanage_35.scala 375:70 stackmanage_35.scala 398:31]
  wire [31:0] _GEN_617 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_582); // @[stackmanage_35.scala 375:70 stackmanage_35.scala 399:31]
  wire [31:0] _GEN_618 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_583); // @[stackmanage_35.scala 375:70 stackmanage_35.scala 400:31]
  wire [31:0] _GEN_619 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_584); // @[stackmanage_35.scala 375:70 stackmanage_35.scala 401:31]
  wire [31:0] _GEN_620 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_585); // @[stackmanage_35.scala 375:70 stackmanage_35.scala 402:31]
  wire [31:0] _GEN_621 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_586); // @[stackmanage_35.scala 375:70 stackmanage_35.scala 403:31]
  wire [31:0] _GEN_622 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_587); // @[stackmanage_35.scala 375:70 stackmanage_35.scala 404:31]
  wire [31:0] _GEN_623 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_588); // @[stackmanage_35.scala 375:70 stackmanage_35.scala 405:31]
  wire [31:0] _GEN_624 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_589); // @[stackmanage_35.scala 375:70 stackmanage_35.scala 406:31]
  wire [31:0] _GEN_625 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_590); // @[stackmanage_35.scala 375:70 stackmanage_35.scala 407:31]
  wire [31:0] _GEN_626 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_591); // @[stackmanage_35.scala 375:70 stackmanage_35.scala 408:31]
  wire [31:0] _GEN_627 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_592); // @[stackmanage_35.scala 375:70 stackmanage_35.scala 409:31]
  wire [31:0] _GEN_628 = LUT_stack_io_push_1 & _T_1 ? $signed(32'sh0) : $signed(_GEN_593); // @[stackmanage_35.scala 375:70 stackmanage_35.scala 410:31]
  reg [31:0] hitT_out_temp; // @[stackmanage_35.scala 1638:34]
  reg [31:0] ray_out_temp; // @[stackmanage_35.scala 1639:35]
  reg [31:0] node_out_temp; // @[stackmanage_35.scala 1640:32]
  reg  pop_valid_1; // @[stackmanage_35.scala 1641:38]
  wire  _T_105 = LUT_stack_io_pop_en; // @[stackmanage_35.scala 1642:29]
  wire [31:0] _GEN_664 = _T_105 & LUT_stack_io_pop_34 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 4056:69 stackmanage_35.scala 4057:29 stackmanage_35.scala 4196:29]
  wire [31:0] _GEN_665 = _T_105 & LUT_stack_io_pop_34 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 4056:69 stackmanage_35.scala 4058:28 stackmanage_35.scala 4197:28]
  wire [31:0] _GEN_667 = _T_105 & LUT_stack_io_pop_33 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 3985:69 stackmanage_35.scala 3986:29]
  wire [31:0] _GEN_668 = _T_105 & LUT_stack_io_pop_33 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 3985:69 stackmanage_35.scala 3987:28]
  wire [31:0] _GEN_670 = _T_105 & LUT_stack_io_pop_33 ? 32'h0 : _GEN_664; // @[stackmanage_35.scala 3985:69 stackmanage_35.scala 4054:29]
  wire [31:0] _GEN_671 = _T_105 & LUT_stack_io_pop_33 ? 32'h0 : _GEN_665; // @[stackmanage_35.scala 3985:69 stackmanage_35.scala 4055:28]
  wire [31:0] _GEN_672 = _T_105 & LUT_stack_io_pop_32 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 3914:69 stackmanage_35.scala 3915:29]
  wire [31:0] _GEN_673 = _T_105 & LUT_stack_io_pop_32 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 3914:69 stackmanage_35.scala 3916:28]
  wire [31:0] _GEN_675 = _T_105 & LUT_stack_io_pop_32 ? 32'h0 : _GEN_667; // @[stackmanage_35.scala 3914:69 stackmanage_35.scala 3981:29]
  wire [31:0] _GEN_676 = _T_105 & LUT_stack_io_pop_32 ? 32'h0 : _GEN_668; // @[stackmanage_35.scala 3914:69 stackmanage_35.scala 3982:28]
  wire [31:0] _GEN_677 = _T_105 & LUT_stack_io_pop_32 ? 32'h0 : _GEN_670; // @[stackmanage_35.scala 3914:69 stackmanage_35.scala 3983:29]
  wire [31:0] _GEN_678 = _T_105 & LUT_stack_io_pop_32 ? 32'h0 : _GEN_671; // @[stackmanage_35.scala 3914:69 stackmanage_35.scala 3984:28]
  wire [31:0] _GEN_679 = _T_105 & LUT_stack_io_pop_31 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 3843:69 stackmanage_35.scala 3844:29]
  wire [31:0] _GEN_680 = _T_105 & LUT_stack_io_pop_31 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 3843:69 stackmanage_35.scala 3845:28]
  wire [31:0] _GEN_682 = _T_105 & LUT_stack_io_pop_31 ? 32'h0 : _GEN_672; // @[stackmanage_35.scala 3843:69 stackmanage_35.scala 3908:29]
  wire [31:0] _GEN_683 = _T_105 & LUT_stack_io_pop_31 ? 32'h0 : _GEN_673; // @[stackmanage_35.scala 3843:69 stackmanage_35.scala 3909:28]
  wire [31:0] _GEN_684 = _T_105 & LUT_stack_io_pop_31 ? 32'h0 : _GEN_675; // @[stackmanage_35.scala 3843:69 stackmanage_35.scala 3910:29]
  wire [31:0] _GEN_685 = _T_105 & LUT_stack_io_pop_31 ? 32'h0 : _GEN_676; // @[stackmanage_35.scala 3843:69 stackmanage_35.scala 3911:28]
  wire [31:0] _GEN_686 = _T_105 & LUT_stack_io_pop_31 ? 32'h0 : _GEN_677; // @[stackmanage_35.scala 3843:69 stackmanage_35.scala 3912:29]
  wire [31:0] _GEN_687 = _T_105 & LUT_stack_io_pop_31 ? 32'h0 : _GEN_678; // @[stackmanage_35.scala 3843:69 stackmanage_35.scala 3913:28]
  wire [31:0] _GEN_688 = _T_105 & LUT_stack_io_pop_30 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 3772:69 stackmanage_35.scala 3773:29]
  wire [31:0] _GEN_689 = _T_105 & LUT_stack_io_pop_30 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 3772:69 stackmanage_35.scala 3774:28]
  wire [31:0] _GEN_691 = _T_105 & LUT_stack_io_pop_30 ? 32'h0 : _GEN_679; // @[stackmanage_35.scala 3772:69 stackmanage_35.scala 3835:29]
  wire [31:0] _GEN_692 = _T_105 & LUT_stack_io_pop_30 ? 32'h0 : _GEN_680; // @[stackmanage_35.scala 3772:69 stackmanage_35.scala 3836:28]
  wire [31:0] _GEN_693 = _T_105 & LUT_stack_io_pop_30 ? 32'h0 : _GEN_682; // @[stackmanage_35.scala 3772:69 stackmanage_35.scala 3837:29]
  wire [31:0] _GEN_694 = _T_105 & LUT_stack_io_pop_30 ? 32'h0 : _GEN_683; // @[stackmanage_35.scala 3772:69 stackmanage_35.scala 3838:28]
  wire [31:0] _GEN_695 = _T_105 & LUT_stack_io_pop_30 ? 32'h0 : _GEN_684; // @[stackmanage_35.scala 3772:69 stackmanage_35.scala 3839:29]
  wire [31:0] _GEN_696 = _T_105 & LUT_stack_io_pop_30 ? 32'h0 : _GEN_685; // @[stackmanage_35.scala 3772:69 stackmanage_35.scala 3840:28]
  wire [31:0] _GEN_697 = _T_105 & LUT_stack_io_pop_30 ? 32'h0 : _GEN_686; // @[stackmanage_35.scala 3772:69 stackmanage_35.scala 3841:29]
  wire [31:0] _GEN_698 = _T_105 & LUT_stack_io_pop_30 ? 32'h0 : _GEN_687; // @[stackmanage_35.scala 3772:69 stackmanage_35.scala 3842:28]
  wire [31:0] _GEN_699 = _T_105 & LUT_stack_io_pop_29 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 3701:69 stackmanage_35.scala 3702:29]
  wire [31:0] _GEN_700 = _T_105 & LUT_stack_io_pop_29 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 3701:69 stackmanage_35.scala 3703:28]
  wire [31:0] _GEN_702 = _T_105 & LUT_stack_io_pop_29 ? 32'h0 : _GEN_688; // @[stackmanage_35.scala 3701:69 stackmanage_35.scala 3762:29]
  wire [31:0] _GEN_703 = _T_105 & LUT_stack_io_pop_29 ? 32'h0 : _GEN_689; // @[stackmanage_35.scala 3701:69 stackmanage_35.scala 3763:29]
  wire [31:0] _GEN_704 = _T_105 & LUT_stack_io_pop_29 ? 32'h0 : _GEN_691; // @[stackmanage_35.scala 3701:69 stackmanage_35.scala 3764:29]
  wire [31:0] _GEN_705 = _T_105 & LUT_stack_io_pop_29 ? 32'h0 : _GEN_692; // @[stackmanage_35.scala 3701:69 stackmanage_35.scala 3765:28]
  wire [31:0] _GEN_706 = _T_105 & LUT_stack_io_pop_29 ? 32'h0 : _GEN_693; // @[stackmanage_35.scala 3701:69 stackmanage_35.scala 3766:29]
  wire [31:0] _GEN_707 = _T_105 & LUT_stack_io_pop_29 ? 32'h0 : _GEN_694; // @[stackmanage_35.scala 3701:69 stackmanage_35.scala 3767:28]
  wire [31:0] _GEN_708 = _T_105 & LUT_stack_io_pop_29 ? 32'h0 : _GEN_695; // @[stackmanage_35.scala 3701:69 stackmanage_35.scala 3768:29]
  wire [31:0] _GEN_709 = _T_105 & LUT_stack_io_pop_29 ? 32'h0 : _GEN_696; // @[stackmanage_35.scala 3701:69 stackmanage_35.scala 3769:28]
  wire [31:0] _GEN_710 = _T_105 & LUT_stack_io_pop_29 ? 32'h0 : _GEN_697; // @[stackmanage_35.scala 3701:69 stackmanage_35.scala 3770:29]
  wire [31:0] _GEN_711 = _T_105 & LUT_stack_io_pop_29 ? 32'h0 : _GEN_698; // @[stackmanage_35.scala 3701:69 stackmanage_35.scala 3771:28]
  wire [31:0] _GEN_712 = _T_105 & LUT_stack_io_pop_28 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 3630:70 stackmanage_35.scala 3631:29]
  wire [31:0] _GEN_713 = _T_105 & LUT_stack_io_pop_28 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 3630:70 stackmanage_35.scala 3632:28]
  wire [31:0] _GEN_715 = _T_105 & LUT_stack_io_pop_28 ? 32'h0 : _GEN_699; // @[stackmanage_35.scala 3630:70 stackmanage_35.scala 3689:29]
  wire [31:0] _GEN_716 = _T_105 & LUT_stack_io_pop_28 ? 32'h0 : _GEN_700; // @[stackmanage_35.scala 3630:70 stackmanage_35.scala 3690:28]
  wire [31:0] _GEN_717 = _T_105 & LUT_stack_io_pop_28 ? 32'h0 : _GEN_702; // @[stackmanage_35.scala 3630:70 stackmanage_35.scala 3691:29]
  wire [31:0] _GEN_718 = _T_105 & LUT_stack_io_pop_28 ? 32'h0 : _GEN_703; // @[stackmanage_35.scala 3630:70 stackmanage_35.scala 3692:29]
  wire [31:0] _GEN_719 = _T_105 & LUT_stack_io_pop_28 ? 32'h0 : _GEN_704; // @[stackmanage_35.scala 3630:70 stackmanage_35.scala 3693:29]
  wire [31:0] _GEN_720 = _T_105 & LUT_stack_io_pop_28 ? 32'h0 : _GEN_705; // @[stackmanage_35.scala 3630:70 stackmanage_35.scala 3694:28]
  wire [31:0] _GEN_721 = _T_105 & LUT_stack_io_pop_28 ? 32'h0 : _GEN_706; // @[stackmanage_35.scala 3630:70 stackmanage_35.scala 3695:29]
  wire [31:0] _GEN_722 = _T_105 & LUT_stack_io_pop_28 ? 32'h0 : _GEN_707; // @[stackmanage_35.scala 3630:70 stackmanage_35.scala 3696:28]
  wire [31:0] _GEN_723 = _T_105 & LUT_stack_io_pop_28 ? 32'h0 : _GEN_708; // @[stackmanage_35.scala 3630:70 stackmanage_35.scala 3697:29]
  wire [31:0] _GEN_724 = _T_105 & LUT_stack_io_pop_28 ? 32'h0 : _GEN_709; // @[stackmanage_35.scala 3630:70 stackmanage_35.scala 3698:28]
  wire [31:0] _GEN_725 = _T_105 & LUT_stack_io_pop_28 ? 32'h0 : _GEN_710; // @[stackmanage_35.scala 3630:70 stackmanage_35.scala 3699:29]
  wire [31:0] _GEN_726 = _T_105 & LUT_stack_io_pop_28 ? 32'h0 : _GEN_711; // @[stackmanage_35.scala 3630:70 stackmanage_35.scala 3700:28]
  wire [31:0] _GEN_727 = _T_105 & LUT_stack_io_pop_27 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 3559:69 stackmanage_35.scala 3560:29]
  wire [31:0] _GEN_728 = _T_105 & LUT_stack_io_pop_27 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 3559:69 stackmanage_35.scala 3561:28]
  wire [31:0] _GEN_730 = _T_105 & LUT_stack_io_pop_27 ? 32'h0 : _GEN_712; // @[stackmanage_35.scala 3559:69 stackmanage_35.scala 3616:29]
  wire [31:0] _GEN_731 = _T_105 & LUT_stack_io_pop_27 ? 32'h0 : _GEN_713; // @[stackmanage_35.scala 3559:69 stackmanage_35.scala 3617:28]
  wire [31:0] _GEN_732 = _T_105 & LUT_stack_io_pop_27 ? 32'h0 : _GEN_715; // @[stackmanage_35.scala 3559:69 stackmanage_35.scala 3618:29]
  wire [31:0] _GEN_733 = _T_105 & LUT_stack_io_pop_27 ? 32'h0 : _GEN_716; // @[stackmanage_35.scala 3559:69 stackmanage_35.scala 3619:28]
  wire [31:0] _GEN_734 = _T_105 & LUT_stack_io_pop_27 ? 32'h0 : _GEN_717; // @[stackmanage_35.scala 3559:69 stackmanage_35.scala 3620:29]
  wire [31:0] _GEN_735 = _T_105 & LUT_stack_io_pop_27 ? 32'h0 : _GEN_718; // @[stackmanage_35.scala 3559:69 stackmanage_35.scala 3621:29]
  wire [31:0] _GEN_736 = _T_105 & LUT_stack_io_pop_27 ? 32'h0 : _GEN_719; // @[stackmanage_35.scala 3559:69 stackmanage_35.scala 3622:29]
  wire [31:0] _GEN_737 = _T_105 & LUT_stack_io_pop_27 ? 32'h0 : _GEN_720; // @[stackmanage_35.scala 3559:69 stackmanage_35.scala 3623:28]
  wire [31:0] _GEN_738 = _T_105 & LUT_stack_io_pop_27 ? 32'h0 : _GEN_721; // @[stackmanage_35.scala 3559:69 stackmanage_35.scala 3624:29]
  wire [31:0] _GEN_739 = _T_105 & LUT_stack_io_pop_27 ? 32'h0 : _GEN_722; // @[stackmanage_35.scala 3559:69 stackmanage_35.scala 3625:28]
  wire [31:0] _GEN_740 = _T_105 & LUT_stack_io_pop_27 ? 32'h0 : _GEN_723; // @[stackmanage_35.scala 3559:69 stackmanage_35.scala 3626:29]
  wire [31:0] _GEN_741 = _T_105 & LUT_stack_io_pop_27 ? 32'h0 : _GEN_724; // @[stackmanage_35.scala 3559:69 stackmanage_35.scala 3627:28]
  wire [31:0] _GEN_742 = _T_105 & LUT_stack_io_pop_27 ? 32'h0 : _GEN_725; // @[stackmanage_35.scala 3559:69 stackmanage_35.scala 3628:29]
  wire [31:0] _GEN_743 = _T_105 & LUT_stack_io_pop_27 ? 32'h0 : _GEN_726; // @[stackmanage_35.scala 3559:69 stackmanage_35.scala 3629:28]
  wire [31:0] _GEN_744 = _T_105 & LUT_stack_io_pop_26 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 3488:70 stackmanage_35.scala 3489:29]
  wire [31:0] _GEN_745 = _T_105 & LUT_stack_io_pop_26 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 3488:70 stackmanage_35.scala 3490:28]
  wire [31:0] _GEN_747 = _T_105 & LUT_stack_io_pop_26 ? 32'h0 : _GEN_727; // @[stackmanage_35.scala 3488:70 stackmanage_35.scala 3543:29]
  wire [31:0] _GEN_748 = _T_105 & LUT_stack_io_pop_26 ? 32'h0 : _GEN_728; // @[stackmanage_35.scala 3488:70 stackmanage_35.scala 3544:28]
  wire [31:0] _GEN_749 = _T_105 & LUT_stack_io_pop_26 ? 32'h0 : _GEN_730; // @[stackmanage_35.scala 3488:70 stackmanage_35.scala 3545:29]
  wire [31:0] _GEN_750 = _T_105 & LUT_stack_io_pop_26 ? 32'h0 : _GEN_731; // @[stackmanage_35.scala 3488:70 stackmanage_35.scala 3546:28]
  wire [31:0] _GEN_751 = _T_105 & LUT_stack_io_pop_26 ? 32'h0 : _GEN_732; // @[stackmanage_35.scala 3488:70 stackmanage_35.scala 3547:29]
  wire [31:0] _GEN_752 = _T_105 & LUT_stack_io_pop_26 ? 32'h0 : _GEN_733; // @[stackmanage_35.scala 3488:70 stackmanage_35.scala 3548:28]
  wire [31:0] _GEN_753 = _T_105 & LUT_stack_io_pop_26 ? 32'h0 : _GEN_734; // @[stackmanage_35.scala 3488:70 stackmanage_35.scala 3549:29]
  wire [31:0] _GEN_754 = _T_105 & LUT_stack_io_pop_26 ? 32'h0 : _GEN_735; // @[stackmanage_35.scala 3488:70 stackmanage_35.scala 3550:29]
  wire [31:0] _GEN_755 = _T_105 & LUT_stack_io_pop_26 ? 32'h0 : _GEN_736; // @[stackmanage_35.scala 3488:70 stackmanage_35.scala 3551:29]
  wire [31:0] _GEN_756 = _T_105 & LUT_stack_io_pop_26 ? 32'h0 : _GEN_737; // @[stackmanage_35.scala 3488:70 stackmanage_35.scala 3552:28]
  wire [31:0] _GEN_757 = _T_105 & LUT_stack_io_pop_26 ? 32'h0 : _GEN_738; // @[stackmanage_35.scala 3488:70 stackmanage_35.scala 3553:29]
  wire [31:0] _GEN_758 = _T_105 & LUT_stack_io_pop_26 ? 32'h0 : _GEN_739; // @[stackmanage_35.scala 3488:70 stackmanage_35.scala 3554:28]
  wire [31:0] _GEN_759 = _T_105 & LUT_stack_io_pop_26 ? 32'h0 : _GEN_740; // @[stackmanage_35.scala 3488:70 stackmanage_35.scala 3555:29]
  wire [31:0] _GEN_760 = _T_105 & LUT_stack_io_pop_26 ? 32'h0 : _GEN_741; // @[stackmanage_35.scala 3488:70 stackmanage_35.scala 3556:28]
  wire [31:0] _GEN_761 = _T_105 & LUT_stack_io_pop_26 ? 32'h0 : _GEN_742; // @[stackmanage_35.scala 3488:70 stackmanage_35.scala 3557:29]
  wire [31:0] _GEN_762 = _T_105 & LUT_stack_io_pop_26 ? 32'h0 : _GEN_743; // @[stackmanage_35.scala 3488:70 stackmanage_35.scala 3558:28]
  wire [31:0] _GEN_763 = _T_105 & LUT_stack_io_pop_25 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 3417:69 stackmanage_35.scala 3418:29]
  wire [31:0] _GEN_764 = _T_105 & LUT_stack_io_pop_25 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 3417:69 stackmanage_35.scala 3419:28]
  wire [31:0] _GEN_766 = _T_105 & LUT_stack_io_pop_25 ? 32'h0 : _GEN_744; // @[stackmanage_35.scala 3417:69 stackmanage_35.scala 3470:29]
  wire [31:0] _GEN_767 = _T_105 & LUT_stack_io_pop_25 ? 32'h0 : _GEN_745; // @[stackmanage_35.scala 3417:69 stackmanage_35.scala 3471:28]
  wire [31:0] _GEN_768 = _T_105 & LUT_stack_io_pop_25 ? 32'h0 : _GEN_747; // @[stackmanage_35.scala 3417:69 stackmanage_35.scala 3472:29]
  wire [31:0] _GEN_769 = _T_105 & LUT_stack_io_pop_25 ? 32'h0 : _GEN_748; // @[stackmanage_35.scala 3417:69 stackmanage_35.scala 3473:28]
  wire [31:0] _GEN_770 = _T_105 & LUT_stack_io_pop_25 ? 32'h0 : _GEN_749; // @[stackmanage_35.scala 3417:69 stackmanage_35.scala 3474:29]
  wire [31:0] _GEN_771 = _T_105 & LUT_stack_io_pop_25 ? 32'h0 : _GEN_750; // @[stackmanage_35.scala 3417:69 stackmanage_35.scala 3475:28]
  wire [31:0] _GEN_772 = _T_105 & LUT_stack_io_pop_25 ? 32'h0 : _GEN_751; // @[stackmanage_35.scala 3417:69 stackmanage_35.scala 3476:29]
  wire [31:0] _GEN_773 = _T_105 & LUT_stack_io_pop_25 ? 32'h0 : _GEN_752; // @[stackmanage_35.scala 3417:69 stackmanage_35.scala 3477:28]
  wire [31:0] _GEN_774 = _T_105 & LUT_stack_io_pop_25 ? 32'h0 : _GEN_753; // @[stackmanage_35.scala 3417:69 stackmanage_35.scala 3478:29]
  wire [31:0] _GEN_775 = _T_105 & LUT_stack_io_pop_25 ? 32'h0 : _GEN_754; // @[stackmanage_35.scala 3417:69 stackmanage_35.scala 3479:29]
  wire [31:0] _GEN_776 = _T_105 & LUT_stack_io_pop_25 ? 32'h0 : _GEN_755; // @[stackmanage_35.scala 3417:69 stackmanage_35.scala 3480:29]
  wire [31:0] _GEN_777 = _T_105 & LUT_stack_io_pop_25 ? 32'h0 : _GEN_756; // @[stackmanage_35.scala 3417:69 stackmanage_35.scala 3481:28]
  wire [31:0] _GEN_778 = _T_105 & LUT_stack_io_pop_25 ? 32'h0 : _GEN_757; // @[stackmanage_35.scala 3417:69 stackmanage_35.scala 3482:29]
  wire [31:0] _GEN_779 = _T_105 & LUT_stack_io_pop_25 ? 32'h0 : _GEN_758; // @[stackmanage_35.scala 3417:69 stackmanage_35.scala 3483:28]
  wire [31:0] _GEN_780 = _T_105 & LUT_stack_io_pop_25 ? 32'h0 : _GEN_759; // @[stackmanage_35.scala 3417:69 stackmanage_35.scala 3484:29]
  wire [31:0] _GEN_781 = _T_105 & LUT_stack_io_pop_25 ? 32'h0 : _GEN_760; // @[stackmanage_35.scala 3417:69 stackmanage_35.scala 3485:28]
  wire [31:0] _GEN_782 = _T_105 & LUT_stack_io_pop_25 ? 32'h0 : _GEN_761; // @[stackmanage_35.scala 3417:69 stackmanage_35.scala 3486:29]
  wire [31:0] _GEN_783 = _T_105 & LUT_stack_io_pop_25 ? 32'h0 : _GEN_762; // @[stackmanage_35.scala 3417:69 stackmanage_35.scala 3487:28]
  wire [31:0] _GEN_784 = _T_105 & LUT_stack_io_pop_24 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 3346:69 stackmanage_35.scala 3347:29]
  wire [31:0] _GEN_785 = _T_105 & LUT_stack_io_pop_24 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 3346:69 stackmanage_35.scala 3348:28]
  wire [31:0] _GEN_787 = _T_105 & LUT_stack_io_pop_24 ? 32'h0 : _GEN_763; // @[stackmanage_35.scala 3346:69 stackmanage_35.scala 3397:29]
  wire [31:0] _GEN_788 = _T_105 & LUT_stack_io_pop_24 ? 32'h0 : _GEN_764; // @[stackmanage_35.scala 3346:69 stackmanage_35.scala 3398:28]
  wire [31:0] _GEN_789 = _T_105 & LUT_stack_io_pop_24 ? 32'h0 : _GEN_766; // @[stackmanage_35.scala 3346:69 stackmanage_35.scala 3399:29]
  wire [31:0] _GEN_790 = _T_105 & LUT_stack_io_pop_24 ? 32'h0 : _GEN_767; // @[stackmanage_35.scala 3346:69 stackmanage_35.scala 3400:28]
  wire [31:0] _GEN_791 = _T_105 & LUT_stack_io_pop_24 ? 32'h0 : _GEN_768; // @[stackmanage_35.scala 3346:69 stackmanage_35.scala 3401:29]
  wire [31:0] _GEN_792 = _T_105 & LUT_stack_io_pop_24 ? 32'h0 : _GEN_769; // @[stackmanage_35.scala 3346:69 stackmanage_35.scala 3402:28]
  wire [31:0] _GEN_793 = _T_105 & LUT_stack_io_pop_24 ? 32'h0 : _GEN_770; // @[stackmanage_35.scala 3346:69 stackmanage_35.scala 3403:29]
  wire [31:0] _GEN_794 = _T_105 & LUT_stack_io_pop_24 ? 32'h0 : _GEN_771; // @[stackmanage_35.scala 3346:69 stackmanage_35.scala 3404:28]
  wire [31:0] _GEN_795 = _T_105 & LUT_stack_io_pop_24 ? 32'h0 : _GEN_772; // @[stackmanage_35.scala 3346:69 stackmanage_35.scala 3405:29]
  wire [31:0] _GEN_796 = _T_105 & LUT_stack_io_pop_24 ? 32'h0 : _GEN_773; // @[stackmanage_35.scala 3346:69 stackmanage_35.scala 3406:28]
  wire [31:0] _GEN_797 = _T_105 & LUT_stack_io_pop_24 ? 32'h0 : _GEN_774; // @[stackmanage_35.scala 3346:69 stackmanage_35.scala 3407:29]
  wire [31:0] _GEN_798 = _T_105 & LUT_stack_io_pop_24 ? 32'h0 : _GEN_775; // @[stackmanage_35.scala 3346:69 stackmanage_35.scala 3408:29]
  wire [31:0] _GEN_799 = _T_105 & LUT_stack_io_pop_24 ? 32'h0 : _GEN_776; // @[stackmanage_35.scala 3346:69 stackmanage_35.scala 3409:29]
  wire [31:0] _GEN_800 = _T_105 & LUT_stack_io_pop_24 ? 32'h0 : _GEN_777; // @[stackmanage_35.scala 3346:69 stackmanage_35.scala 3410:28]
  wire [31:0] _GEN_801 = _T_105 & LUT_stack_io_pop_24 ? 32'h0 : _GEN_778; // @[stackmanage_35.scala 3346:69 stackmanage_35.scala 3411:29]
  wire [31:0] _GEN_802 = _T_105 & LUT_stack_io_pop_24 ? 32'h0 : _GEN_779; // @[stackmanage_35.scala 3346:69 stackmanage_35.scala 3412:28]
  wire [31:0] _GEN_803 = _T_105 & LUT_stack_io_pop_24 ? 32'h0 : _GEN_780; // @[stackmanage_35.scala 3346:69 stackmanage_35.scala 3413:29]
  wire [31:0] _GEN_804 = _T_105 & LUT_stack_io_pop_24 ? 32'h0 : _GEN_781; // @[stackmanage_35.scala 3346:69 stackmanage_35.scala 3414:28]
  wire [31:0] _GEN_805 = _T_105 & LUT_stack_io_pop_24 ? 32'h0 : _GEN_782; // @[stackmanage_35.scala 3346:69 stackmanage_35.scala 3415:29]
  wire [31:0] _GEN_806 = _T_105 & LUT_stack_io_pop_24 ? 32'h0 : _GEN_783; // @[stackmanage_35.scala 3346:69 stackmanage_35.scala 3416:28]
  wire [31:0] _GEN_807 = _T_105 & LUT_stack_io_pop_23 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 3275:69 stackmanage_35.scala 3276:29]
  wire [31:0] _GEN_808 = _T_105 & LUT_stack_io_pop_23 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 3275:69 stackmanage_35.scala 3277:28]
  wire [31:0] _GEN_810 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_784; // @[stackmanage_35.scala 3275:69 stackmanage_35.scala 3324:29]
  wire [31:0] _GEN_811 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_785; // @[stackmanage_35.scala 3275:69 stackmanage_35.scala 3325:28]
  wire [31:0] _GEN_812 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_787; // @[stackmanage_35.scala 3275:69 stackmanage_35.scala 3326:29]
  wire [31:0] _GEN_813 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_788; // @[stackmanage_35.scala 3275:69 stackmanage_35.scala 3327:28]
  wire [31:0] _GEN_814 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_789; // @[stackmanage_35.scala 3275:69 stackmanage_35.scala 3328:29]
  wire [31:0] _GEN_815 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_790; // @[stackmanage_35.scala 3275:69 stackmanage_35.scala 3329:28]
  wire [31:0] _GEN_816 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_791; // @[stackmanage_35.scala 3275:69 stackmanage_35.scala 3330:29]
  wire [31:0] _GEN_817 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_792; // @[stackmanage_35.scala 3275:69 stackmanage_35.scala 3331:28]
  wire [31:0] _GEN_818 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_793; // @[stackmanage_35.scala 3275:69 stackmanage_35.scala 3332:29]
  wire [31:0] _GEN_819 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_794; // @[stackmanage_35.scala 3275:69 stackmanage_35.scala 3333:28]
  wire [31:0] _GEN_820 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_795; // @[stackmanage_35.scala 3275:69 stackmanage_35.scala 3334:29]
  wire [31:0] _GEN_821 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_796; // @[stackmanage_35.scala 3275:69 stackmanage_35.scala 3335:28]
  wire [31:0] _GEN_822 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_797; // @[stackmanage_35.scala 3275:69 stackmanage_35.scala 3336:29]
  wire [31:0] _GEN_823 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_798; // @[stackmanage_35.scala 3275:69 stackmanage_35.scala 3337:29]
  wire [31:0] _GEN_824 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_799; // @[stackmanage_35.scala 3275:69 stackmanage_35.scala 3338:29]
  wire [31:0] _GEN_825 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_800; // @[stackmanage_35.scala 3275:69 stackmanage_35.scala 3339:28]
  wire [31:0] _GEN_826 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_801; // @[stackmanage_35.scala 3275:69 stackmanage_35.scala 3340:29]
  wire [31:0] _GEN_827 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_802; // @[stackmanage_35.scala 3275:69 stackmanage_35.scala 3341:28]
  wire [31:0] _GEN_828 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_803; // @[stackmanage_35.scala 3275:69 stackmanage_35.scala 3342:29]
  wire [31:0] _GEN_829 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_804; // @[stackmanage_35.scala 3275:69 stackmanage_35.scala 3343:28]
  wire [31:0] _GEN_830 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_805; // @[stackmanage_35.scala 3275:69 stackmanage_35.scala 3344:29]
  wire [31:0] _GEN_831 = _T_105 & LUT_stack_io_pop_23 ? 32'h0 : _GEN_806; // @[stackmanage_35.scala 3275:69 stackmanage_35.scala 3345:28]
  wire [31:0] _GEN_832 = _T_105 & LUT_stack_io_pop_22 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 3204:69 stackmanage_35.scala 3205:29]
  wire [31:0] _GEN_833 = _T_105 & LUT_stack_io_pop_22 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 3204:69 stackmanage_35.scala 3206:28]
  wire [31:0] _GEN_835 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_807; // @[stackmanage_35.scala 3204:69 stackmanage_35.scala 3251:29]
  wire [31:0] _GEN_836 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_808; // @[stackmanage_35.scala 3204:69 stackmanage_35.scala 3252:28]
  wire [31:0] _GEN_837 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_810; // @[stackmanage_35.scala 3204:69 stackmanage_35.scala 3253:29]
  wire [31:0] _GEN_838 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_811; // @[stackmanage_35.scala 3204:69 stackmanage_35.scala 3254:28]
  wire [31:0] _GEN_839 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_812; // @[stackmanage_35.scala 3204:69 stackmanage_35.scala 3255:29]
  wire [31:0] _GEN_840 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_813; // @[stackmanage_35.scala 3204:69 stackmanage_35.scala 3256:28]
  wire [31:0] _GEN_841 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_814; // @[stackmanage_35.scala 3204:69 stackmanage_35.scala 3257:29]
  wire [31:0] _GEN_842 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_815; // @[stackmanage_35.scala 3204:69 stackmanage_35.scala 3258:28]
  wire [31:0] _GEN_843 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_816; // @[stackmanage_35.scala 3204:69 stackmanage_35.scala 3259:29]
  wire [31:0] _GEN_844 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_817; // @[stackmanage_35.scala 3204:69 stackmanage_35.scala 3260:28]
  wire [31:0] _GEN_845 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_818; // @[stackmanage_35.scala 3204:69 stackmanage_35.scala 3261:29]
  wire [31:0] _GEN_846 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_819; // @[stackmanage_35.scala 3204:69 stackmanage_35.scala 3262:28]
  wire [31:0] _GEN_847 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_820; // @[stackmanage_35.scala 3204:69 stackmanage_35.scala 3263:29]
  wire [31:0] _GEN_848 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_821; // @[stackmanage_35.scala 3204:69 stackmanage_35.scala 3264:28]
  wire [31:0] _GEN_849 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_822; // @[stackmanage_35.scala 3204:69 stackmanage_35.scala 3265:29]
  wire [31:0] _GEN_850 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_823; // @[stackmanage_35.scala 3204:69 stackmanage_35.scala 3266:29]
  wire [31:0] _GEN_851 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_824; // @[stackmanage_35.scala 3204:69 stackmanage_35.scala 3267:29]
  wire [31:0] _GEN_852 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_825; // @[stackmanage_35.scala 3204:69 stackmanage_35.scala 3268:28]
  wire [31:0] _GEN_853 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_826; // @[stackmanage_35.scala 3204:69 stackmanage_35.scala 3269:29]
  wire [31:0] _GEN_854 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_827; // @[stackmanage_35.scala 3204:69 stackmanage_35.scala 3270:28]
  wire [31:0] _GEN_855 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_828; // @[stackmanage_35.scala 3204:69 stackmanage_35.scala 3271:29]
  wire [31:0] _GEN_856 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_829; // @[stackmanage_35.scala 3204:69 stackmanage_35.scala 3272:28]
  wire [31:0] _GEN_857 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_830; // @[stackmanage_35.scala 3204:69 stackmanage_35.scala 3273:29]
  wire [31:0] _GEN_858 = _T_105 & LUT_stack_io_pop_22 ? 32'h0 : _GEN_831; // @[stackmanage_35.scala 3204:69 stackmanage_35.scala 3274:28]
  wire [31:0] _GEN_859 = _T_105 & LUT_stack_io_pop_21 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 3133:69 stackmanage_35.scala 3134:29]
  wire [31:0] _GEN_860 = _T_105 & LUT_stack_io_pop_21 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 3133:69 stackmanage_35.scala 3135:28]
  wire [31:0] _GEN_862 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_832; // @[stackmanage_35.scala 3133:69 stackmanage_35.scala 3178:29]
  wire [31:0] _GEN_863 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_833; // @[stackmanage_35.scala 3133:69 stackmanage_35.scala 3179:28]
  wire [31:0] _GEN_864 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_835; // @[stackmanage_35.scala 3133:69 stackmanage_35.scala 3180:29]
  wire [31:0] _GEN_865 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_836; // @[stackmanage_35.scala 3133:69 stackmanage_35.scala 3181:28]
  wire [31:0] _GEN_866 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_837; // @[stackmanage_35.scala 3133:69 stackmanage_35.scala 3182:29]
  wire [31:0] _GEN_867 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_838; // @[stackmanage_35.scala 3133:69 stackmanage_35.scala 3183:28]
  wire [31:0] _GEN_868 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_839; // @[stackmanage_35.scala 3133:69 stackmanage_35.scala 3184:29]
  wire [31:0] _GEN_869 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_840; // @[stackmanage_35.scala 3133:69 stackmanage_35.scala 3185:28]
  wire [31:0] _GEN_870 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_841; // @[stackmanage_35.scala 3133:69 stackmanage_35.scala 3186:29]
  wire [31:0] _GEN_871 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_842; // @[stackmanage_35.scala 3133:69 stackmanage_35.scala 3187:28]
  wire [31:0] _GEN_872 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_843; // @[stackmanage_35.scala 3133:69 stackmanage_35.scala 3188:29]
  wire [31:0] _GEN_873 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_844; // @[stackmanage_35.scala 3133:69 stackmanage_35.scala 3189:28]
  wire [31:0] _GEN_874 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_845; // @[stackmanage_35.scala 3133:69 stackmanage_35.scala 3190:29]
  wire [31:0] _GEN_875 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_846; // @[stackmanage_35.scala 3133:69 stackmanage_35.scala 3191:28]
  wire [31:0] _GEN_876 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_847; // @[stackmanage_35.scala 3133:69 stackmanage_35.scala 3192:29]
  wire [31:0] _GEN_877 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_848; // @[stackmanage_35.scala 3133:69 stackmanage_35.scala 3193:28]
  wire [31:0] _GEN_878 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_849; // @[stackmanage_35.scala 3133:69 stackmanage_35.scala 3194:29]
  wire [31:0] _GEN_879 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_850; // @[stackmanage_35.scala 3133:69 stackmanage_35.scala 3195:29]
  wire [31:0] _GEN_880 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_851; // @[stackmanage_35.scala 3133:69 stackmanage_35.scala 3196:29]
  wire [31:0] _GEN_881 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_852; // @[stackmanage_35.scala 3133:69 stackmanage_35.scala 3197:28]
  wire [31:0] _GEN_882 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_853; // @[stackmanage_35.scala 3133:69 stackmanage_35.scala 3198:29]
  wire [31:0] _GEN_883 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_854; // @[stackmanage_35.scala 3133:69 stackmanage_35.scala 3199:28]
  wire [31:0] _GEN_884 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_855; // @[stackmanage_35.scala 3133:69 stackmanage_35.scala 3200:29]
  wire [31:0] _GEN_885 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_856; // @[stackmanage_35.scala 3133:69 stackmanage_35.scala 3201:28]
  wire [31:0] _GEN_886 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_857; // @[stackmanage_35.scala 3133:69 stackmanage_35.scala 3202:29]
  wire [31:0] _GEN_887 = _T_105 & LUT_stack_io_pop_21 ? 32'h0 : _GEN_858; // @[stackmanage_35.scala 3133:69 stackmanage_35.scala 3203:28]
  wire [31:0] _GEN_888 = _T_105 & LUT_stack_io_pop_20 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 3062:69 stackmanage_35.scala 3063:29]
  wire [31:0] _GEN_889 = _T_105 & LUT_stack_io_pop_20 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 3062:69 stackmanage_35.scala 3064:28]
  wire [31:0] _GEN_891 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_859; // @[stackmanage_35.scala 3062:69 stackmanage_35.scala 3105:29]
  wire [31:0] _GEN_892 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_860; // @[stackmanage_35.scala 3062:69 stackmanage_35.scala 3106:28]
  wire [31:0] _GEN_893 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_862; // @[stackmanage_35.scala 3062:69 stackmanage_35.scala 3107:29]
  wire [31:0] _GEN_894 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_863; // @[stackmanage_35.scala 3062:69 stackmanage_35.scala 3108:28]
  wire [31:0] _GEN_895 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_864; // @[stackmanage_35.scala 3062:69 stackmanage_35.scala 3109:29]
  wire [31:0] _GEN_896 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_865; // @[stackmanage_35.scala 3062:69 stackmanage_35.scala 3110:28]
  wire [31:0] _GEN_897 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_866; // @[stackmanage_35.scala 3062:69 stackmanage_35.scala 3111:29]
  wire [31:0] _GEN_898 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_867; // @[stackmanage_35.scala 3062:69 stackmanage_35.scala 3112:28]
  wire [31:0] _GEN_899 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_868; // @[stackmanage_35.scala 3062:69 stackmanage_35.scala 3113:29]
  wire [31:0] _GEN_900 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_869; // @[stackmanage_35.scala 3062:69 stackmanage_35.scala 3114:28]
  wire [31:0] _GEN_901 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_870; // @[stackmanage_35.scala 3062:69 stackmanage_35.scala 3115:29]
  wire [31:0] _GEN_902 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_871; // @[stackmanage_35.scala 3062:69 stackmanage_35.scala 3116:28]
  wire [31:0] _GEN_903 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_872; // @[stackmanage_35.scala 3062:69 stackmanage_35.scala 3117:29]
  wire [31:0] _GEN_904 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_873; // @[stackmanage_35.scala 3062:69 stackmanage_35.scala 3118:28]
  wire [31:0] _GEN_905 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_874; // @[stackmanage_35.scala 3062:69 stackmanage_35.scala 3119:29]
  wire [31:0] _GEN_906 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_875; // @[stackmanage_35.scala 3062:69 stackmanage_35.scala 3120:28]
  wire [31:0] _GEN_907 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_876; // @[stackmanage_35.scala 3062:69 stackmanage_35.scala 3121:29]
  wire [31:0] _GEN_908 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_877; // @[stackmanage_35.scala 3062:69 stackmanage_35.scala 3122:28]
  wire [31:0] _GEN_909 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_878; // @[stackmanage_35.scala 3062:69 stackmanage_35.scala 3123:29]
  wire [31:0] _GEN_910 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_879; // @[stackmanage_35.scala 3062:69 stackmanage_35.scala 3124:29]
  wire [31:0] _GEN_911 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_880; // @[stackmanage_35.scala 3062:69 stackmanage_35.scala 3125:29]
  wire [31:0] _GEN_912 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_881; // @[stackmanage_35.scala 3062:69 stackmanage_35.scala 3126:28]
  wire [31:0] _GEN_913 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_882; // @[stackmanage_35.scala 3062:69 stackmanage_35.scala 3127:29]
  wire [31:0] _GEN_914 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_883; // @[stackmanage_35.scala 3062:69 stackmanage_35.scala 3128:28]
  wire [31:0] _GEN_915 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_884; // @[stackmanage_35.scala 3062:69 stackmanage_35.scala 3129:29]
  wire [31:0] _GEN_916 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_885; // @[stackmanage_35.scala 3062:69 stackmanage_35.scala 3130:28]
  wire [31:0] _GEN_917 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_886; // @[stackmanage_35.scala 3062:69 stackmanage_35.scala 3131:29]
  wire [31:0] _GEN_918 = _T_105 & LUT_stack_io_pop_20 ? 32'h0 : _GEN_887; // @[stackmanage_35.scala 3062:69 stackmanage_35.scala 3132:28]
  wire [31:0] _GEN_919 = _T_105 & LUT_stack_io_pop_19 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 2991:69 stackmanage_35.scala 2992:29]
  wire [31:0] _GEN_920 = _T_105 & LUT_stack_io_pop_19 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 2991:69 stackmanage_35.scala 2993:28]
  wire [31:0] _GEN_922 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_888; // @[stackmanage_35.scala 2991:69 stackmanage_35.scala 3032:29]
  wire [31:0] _GEN_923 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_889; // @[stackmanage_35.scala 2991:69 stackmanage_35.scala 3033:29]
  wire [31:0] _GEN_924 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_891; // @[stackmanage_35.scala 2991:69 stackmanage_35.scala 3034:29]
  wire [31:0] _GEN_925 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_892; // @[stackmanage_35.scala 2991:69 stackmanage_35.scala 3035:28]
  wire [31:0] _GEN_926 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_893; // @[stackmanage_35.scala 2991:69 stackmanage_35.scala 3036:29]
  wire [31:0] _GEN_927 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_894; // @[stackmanage_35.scala 2991:69 stackmanage_35.scala 3037:28]
  wire [31:0] _GEN_928 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_895; // @[stackmanage_35.scala 2991:69 stackmanage_35.scala 3038:29]
  wire [31:0] _GEN_929 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_896; // @[stackmanage_35.scala 2991:69 stackmanage_35.scala 3039:28]
  wire [31:0] _GEN_930 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_897; // @[stackmanage_35.scala 2991:69 stackmanage_35.scala 3040:29]
  wire [31:0] _GEN_931 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_898; // @[stackmanage_35.scala 2991:69 stackmanage_35.scala 3041:28]
  wire [31:0] _GEN_932 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_899; // @[stackmanage_35.scala 2991:69 stackmanage_35.scala 3042:29]
  wire [31:0] _GEN_933 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_900; // @[stackmanage_35.scala 2991:69 stackmanage_35.scala 3043:28]
  wire [31:0] _GEN_934 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_901; // @[stackmanage_35.scala 2991:69 stackmanage_35.scala 3044:29]
  wire [31:0] _GEN_935 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_902; // @[stackmanage_35.scala 2991:69 stackmanage_35.scala 3045:28]
  wire [31:0] _GEN_936 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_903; // @[stackmanage_35.scala 2991:69 stackmanage_35.scala 3046:29]
  wire [31:0] _GEN_937 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_904; // @[stackmanage_35.scala 2991:69 stackmanage_35.scala 3047:28]
  wire [31:0] _GEN_938 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_905; // @[stackmanage_35.scala 2991:69 stackmanage_35.scala 3048:29]
  wire [31:0] _GEN_939 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_906; // @[stackmanage_35.scala 2991:69 stackmanage_35.scala 3049:28]
  wire [31:0] _GEN_940 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_907; // @[stackmanage_35.scala 2991:69 stackmanage_35.scala 3050:29]
  wire [31:0] _GEN_941 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_908; // @[stackmanage_35.scala 2991:69 stackmanage_35.scala 3051:28]
  wire [31:0] _GEN_942 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_909; // @[stackmanage_35.scala 2991:69 stackmanage_35.scala 3052:29]
  wire [31:0] _GEN_943 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_910; // @[stackmanage_35.scala 2991:69 stackmanage_35.scala 3053:29]
  wire [31:0] _GEN_944 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_911; // @[stackmanage_35.scala 2991:69 stackmanage_35.scala 3054:29]
  wire [31:0] _GEN_945 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_912; // @[stackmanage_35.scala 2991:69 stackmanage_35.scala 3055:28]
  wire [31:0] _GEN_946 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_913; // @[stackmanage_35.scala 2991:69 stackmanage_35.scala 3056:29]
  wire [31:0] _GEN_947 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_914; // @[stackmanage_35.scala 2991:69 stackmanage_35.scala 3057:28]
  wire [31:0] _GEN_948 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_915; // @[stackmanage_35.scala 2991:69 stackmanage_35.scala 3058:29]
  wire [31:0] _GEN_949 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_916; // @[stackmanage_35.scala 2991:69 stackmanage_35.scala 3059:28]
  wire [31:0] _GEN_950 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_917; // @[stackmanage_35.scala 2991:69 stackmanage_35.scala 3060:29]
  wire [31:0] _GEN_951 = _T_105 & LUT_stack_io_pop_19 ? 32'h0 : _GEN_918; // @[stackmanage_35.scala 2991:69 stackmanage_35.scala 3061:28]
  wire [31:0] _GEN_952 = _T_105 & LUT_stack_io_pop_18 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 2920:69 stackmanage_35.scala 2921:29]
  wire [31:0] _GEN_953 = _T_105 & LUT_stack_io_pop_18 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 2920:69 stackmanage_35.scala 2922:28]
  wire [31:0] _GEN_955 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_919; // @[stackmanage_35.scala 2920:69 stackmanage_35.scala 2959:29]
  wire [31:0] _GEN_956 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_920; // @[stackmanage_35.scala 2920:69 stackmanage_35.scala 2960:28]
  wire [31:0] _GEN_957 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_922; // @[stackmanage_35.scala 2920:69 stackmanage_35.scala 2961:29]
  wire [31:0] _GEN_958 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_923; // @[stackmanage_35.scala 2920:69 stackmanage_35.scala 2962:29]
  wire [31:0] _GEN_959 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_924; // @[stackmanage_35.scala 2920:69 stackmanage_35.scala 2963:29]
  wire [31:0] _GEN_960 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_925; // @[stackmanage_35.scala 2920:69 stackmanage_35.scala 2964:28]
  wire [31:0] _GEN_961 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_926; // @[stackmanage_35.scala 2920:69 stackmanage_35.scala 2965:29]
  wire [31:0] _GEN_962 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_927; // @[stackmanage_35.scala 2920:69 stackmanage_35.scala 2966:28]
  wire [31:0] _GEN_963 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_928; // @[stackmanage_35.scala 2920:69 stackmanage_35.scala 2967:29]
  wire [31:0] _GEN_964 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_929; // @[stackmanage_35.scala 2920:69 stackmanage_35.scala 2968:28]
  wire [31:0] _GEN_965 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_930; // @[stackmanage_35.scala 2920:69 stackmanage_35.scala 2969:29]
  wire [31:0] _GEN_966 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_931; // @[stackmanage_35.scala 2920:69 stackmanage_35.scala 2970:28]
  wire [31:0] _GEN_967 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_932; // @[stackmanage_35.scala 2920:69 stackmanage_35.scala 2971:29]
  wire [31:0] _GEN_968 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_933; // @[stackmanage_35.scala 2920:69 stackmanage_35.scala 2972:28]
  wire [31:0] _GEN_969 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_934; // @[stackmanage_35.scala 2920:69 stackmanage_35.scala 2973:29]
  wire [31:0] _GEN_970 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_935; // @[stackmanage_35.scala 2920:69 stackmanage_35.scala 2974:28]
  wire [31:0] _GEN_971 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_936; // @[stackmanage_35.scala 2920:69 stackmanage_35.scala 2975:29]
  wire [31:0] _GEN_972 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_937; // @[stackmanage_35.scala 2920:69 stackmanage_35.scala 2976:28]
  wire [31:0] _GEN_973 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_938; // @[stackmanage_35.scala 2920:69 stackmanage_35.scala 2977:29]
  wire [31:0] _GEN_974 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_939; // @[stackmanage_35.scala 2920:69 stackmanage_35.scala 2978:28]
  wire [31:0] _GEN_975 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_940; // @[stackmanage_35.scala 2920:69 stackmanage_35.scala 2979:29]
  wire [31:0] _GEN_976 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_941; // @[stackmanage_35.scala 2920:69 stackmanage_35.scala 2980:28]
  wire [31:0] _GEN_977 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_942; // @[stackmanage_35.scala 2920:69 stackmanage_35.scala 2981:29]
  wire [31:0] _GEN_978 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_943; // @[stackmanage_35.scala 2920:69 stackmanage_35.scala 2982:29]
  wire [31:0] _GEN_979 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_944; // @[stackmanage_35.scala 2920:69 stackmanage_35.scala 2983:29]
  wire [31:0] _GEN_980 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_945; // @[stackmanage_35.scala 2920:69 stackmanage_35.scala 2984:28]
  wire [31:0] _GEN_981 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_946; // @[stackmanage_35.scala 2920:69 stackmanage_35.scala 2985:29]
  wire [31:0] _GEN_982 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_947; // @[stackmanage_35.scala 2920:69 stackmanage_35.scala 2986:28]
  wire [31:0] _GEN_983 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_948; // @[stackmanage_35.scala 2920:69 stackmanage_35.scala 2987:29]
  wire [31:0] _GEN_984 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_949; // @[stackmanage_35.scala 2920:69 stackmanage_35.scala 2988:28]
  wire [31:0] _GEN_985 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_950; // @[stackmanage_35.scala 2920:69 stackmanage_35.scala 2989:29]
  wire [31:0] _GEN_986 = _T_105 & LUT_stack_io_pop_18 ? 32'h0 : _GEN_951; // @[stackmanage_35.scala 2920:69 stackmanage_35.scala 2990:28]
  wire [31:0] _GEN_987 = _T_105 & LUT_stack_io_pop_17 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 2849:69 stackmanage_35.scala 2850:29]
  wire [31:0] _GEN_988 = _T_105 & LUT_stack_io_pop_17 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 2849:69 stackmanage_35.scala 2851:28]
  wire [31:0] _GEN_990 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_952; // @[stackmanage_35.scala 2849:69 stackmanage_35.scala 2886:29]
  wire [31:0] _GEN_991 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_953; // @[stackmanage_35.scala 2849:69 stackmanage_35.scala 2887:28]
  wire [31:0] _GEN_992 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_955; // @[stackmanage_35.scala 2849:69 stackmanage_35.scala 2888:29]
  wire [31:0] _GEN_993 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_956; // @[stackmanage_35.scala 2849:69 stackmanage_35.scala 2889:28]
  wire [31:0] _GEN_994 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_957; // @[stackmanage_35.scala 2849:69 stackmanage_35.scala 2890:29]
  wire [31:0] _GEN_995 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_958; // @[stackmanage_35.scala 2849:69 stackmanage_35.scala 2891:29]
  wire [31:0] _GEN_996 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_959; // @[stackmanage_35.scala 2849:69 stackmanage_35.scala 2892:29]
  wire [31:0] _GEN_997 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_960; // @[stackmanage_35.scala 2849:69 stackmanage_35.scala 2893:28]
  wire [31:0] _GEN_998 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_961; // @[stackmanage_35.scala 2849:69 stackmanage_35.scala 2894:29]
  wire [31:0] _GEN_999 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_962; // @[stackmanage_35.scala 2849:69 stackmanage_35.scala 2895:28]
  wire [31:0] _GEN_1000 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_963; // @[stackmanage_35.scala 2849:69 stackmanage_35.scala 2896:29]
  wire [31:0] _GEN_1001 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_964; // @[stackmanage_35.scala 2849:69 stackmanage_35.scala 2897:28]
  wire [31:0] _GEN_1002 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_965; // @[stackmanage_35.scala 2849:69 stackmanage_35.scala 2898:29]
  wire [31:0] _GEN_1003 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_966; // @[stackmanage_35.scala 2849:69 stackmanage_35.scala 2899:28]
  wire [31:0] _GEN_1004 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_967; // @[stackmanage_35.scala 2849:69 stackmanage_35.scala 2900:29]
  wire [31:0] _GEN_1005 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_968; // @[stackmanage_35.scala 2849:69 stackmanage_35.scala 2901:28]
  wire [31:0] _GEN_1006 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_969; // @[stackmanage_35.scala 2849:69 stackmanage_35.scala 2902:29]
  wire [31:0] _GEN_1007 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_970; // @[stackmanage_35.scala 2849:69 stackmanage_35.scala 2903:28]
  wire [31:0] _GEN_1008 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_971; // @[stackmanage_35.scala 2849:69 stackmanage_35.scala 2904:29]
  wire [31:0] _GEN_1009 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_972; // @[stackmanage_35.scala 2849:69 stackmanage_35.scala 2905:28]
  wire [31:0] _GEN_1010 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_973; // @[stackmanage_35.scala 2849:69 stackmanage_35.scala 2906:29]
  wire [31:0] _GEN_1011 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_974; // @[stackmanage_35.scala 2849:69 stackmanage_35.scala 2907:28]
  wire [31:0] _GEN_1012 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_975; // @[stackmanage_35.scala 2849:69 stackmanage_35.scala 2908:29]
  wire [31:0] _GEN_1013 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_976; // @[stackmanage_35.scala 2849:69 stackmanage_35.scala 2909:28]
  wire [31:0] _GEN_1014 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_977; // @[stackmanage_35.scala 2849:69 stackmanage_35.scala 2910:29]
  wire [31:0] _GEN_1015 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_978; // @[stackmanage_35.scala 2849:69 stackmanage_35.scala 2911:29]
  wire [31:0] _GEN_1016 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_979; // @[stackmanage_35.scala 2849:69 stackmanage_35.scala 2912:29]
  wire [31:0] _GEN_1017 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_980; // @[stackmanage_35.scala 2849:69 stackmanage_35.scala 2913:28]
  wire [31:0] _GEN_1018 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_981; // @[stackmanage_35.scala 2849:69 stackmanage_35.scala 2914:29]
  wire [31:0] _GEN_1019 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_982; // @[stackmanage_35.scala 2849:69 stackmanage_35.scala 2915:28]
  wire [31:0] _GEN_1020 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_983; // @[stackmanage_35.scala 2849:69 stackmanage_35.scala 2916:29]
  wire [31:0] _GEN_1021 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_984; // @[stackmanage_35.scala 2849:69 stackmanage_35.scala 2917:28]
  wire [31:0] _GEN_1022 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_985; // @[stackmanage_35.scala 2849:69 stackmanage_35.scala 2918:29]
  wire [31:0] _GEN_1023 = _T_105 & LUT_stack_io_pop_17 ? 32'h0 : _GEN_986; // @[stackmanage_35.scala 2849:69 stackmanage_35.scala 2919:28]
  wire [31:0] _GEN_1024 = _T_105 & LUT_stack_io_pop_16 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 2778:69 stackmanage_35.scala 2779:29]
  wire [31:0] _GEN_1025 = _T_105 & LUT_stack_io_pop_16 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 2778:69 stackmanage_35.scala 2780:28]
  wire [31:0] _GEN_1027 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_987; // @[stackmanage_35.scala 2778:69 stackmanage_35.scala 2813:29]
  wire [31:0] _GEN_1028 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_988; // @[stackmanage_35.scala 2778:69 stackmanage_35.scala 2814:28]
  wire [31:0] _GEN_1029 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_990; // @[stackmanage_35.scala 2778:69 stackmanage_35.scala 2815:29]
  wire [31:0] _GEN_1030 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_991; // @[stackmanage_35.scala 2778:69 stackmanage_35.scala 2816:28]
  wire [31:0] _GEN_1031 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_992; // @[stackmanage_35.scala 2778:69 stackmanage_35.scala 2817:29]
  wire [31:0] _GEN_1032 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_993; // @[stackmanage_35.scala 2778:69 stackmanage_35.scala 2818:28]
  wire [31:0] _GEN_1033 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_994; // @[stackmanage_35.scala 2778:69 stackmanage_35.scala 2819:29]
  wire [31:0] _GEN_1034 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_995; // @[stackmanage_35.scala 2778:69 stackmanage_35.scala 2820:29]
  wire [31:0] _GEN_1035 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_996; // @[stackmanage_35.scala 2778:69 stackmanage_35.scala 2821:29]
  wire [31:0] _GEN_1036 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_997; // @[stackmanage_35.scala 2778:69 stackmanage_35.scala 2822:28]
  wire [31:0] _GEN_1037 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_998; // @[stackmanage_35.scala 2778:69 stackmanage_35.scala 2823:29]
  wire [31:0] _GEN_1038 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_999; // @[stackmanage_35.scala 2778:69 stackmanage_35.scala 2824:28]
  wire [31:0] _GEN_1039 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1000; // @[stackmanage_35.scala 2778:69 stackmanage_35.scala 2825:29]
  wire [31:0] _GEN_1040 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1001; // @[stackmanage_35.scala 2778:69 stackmanage_35.scala 2826:28]
  wire [31:0] _GEN_1041 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1002; // @[stackmanage_35.scala 2778:69 stackmanage_35.scala 2827:29]
  wire [31:0] _GEN_1042 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1003; // @[stackmanage_35.scala 2778:69 stackmanage_35.scala 2828:28]
  wire [31:0] _GEN_1043 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1004; // @[stackmanage_35.scala 2778:69 stackmanage_35.scala 2829:29]
  wire [31:0] _GEN_1044 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1005; // @[stackmanage_35.scala 2778:69 stackmanage_35.scala 2830:28]
  wire [31:0] _GEN_1045 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1006; // @[stackmanage_35.scala 2778:69 stackmanage_35.scala 2831:29]
  wire [31:0] _GEN_1046 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1007; // @[stackmanage_35.scala 2778:69 stackmanage_35.scala 2832:28]
  wire [31:0] _GEN_1047 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1008; // @[stackmanage_35.scala 2778:69 stackmanage_35.scala 2833:29]
  wire [31:0] _GEN_1048 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1009; // @[stackmanage_35.scala 2778:69 stackmanage_35.scala 2834:28]
  wire [31:0] _GEN_1049 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1010; // @[stackmanage_35.scala 2778:69 stackmanage_35.scala 2835:29]
  wire [31:0] _GEN_1050 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1011; // @[stackmanage_35.scala 2778:69 stackmanage_35.scala 2836:28]
  wire [31:0] _GEN_1051 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1012; // @[stackmanage_35.scala 2778:69 stackmanage_35.scala 2837:29]
  wire [31:0] _GEN_1052 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1013; // @[stackmanage_35.scala 2778:69 stackmanage_35.scala 2838:28]
  wire [31:0] _GEN_1053 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1014; // @[stackmanage_35.scala 2778:69 stackmanage_35.scala 2839:29]
  wire [31:0] _GEN_1054 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1015; // @[stackmanage_35.scala 2778:69 stackmanage_35.scala 2840:29]
  wire [31:0] _GEN_1055 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1016; // @[stackmanage_35.scala 2778:69 stackmanage_35.scala 2841:29]
  wire [31:0] _GEN_1056 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1017; // @[stackmanage_35.scala 2778:69 stackmanage_35.scala 2842:28]
  wire [31:0] _GEN_1057 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1018; // @[stackmanage_35.scala 2778:69 stackmanage_35.scala 2843:29]
  wire [31:0] _GEN_1058 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1019; // @[stackmanage_35.scala 2778:69 stackmanage_35.scala 2844:28]
  wire [31:0] _GEN_1059 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1020; // @[stackmanage_35.scala 2778:69 stackmanage_35.scala 2845:29]
  wire [31:0] _GEN_1060 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1021; // @[stackmanage_35.scala 2778:69 stackmanage_35.scala 2846:28]
  wire [31:0] _GEN_1061 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1022; // @[stackmanage_35.scala 2778:69 stackmanage_35.scala 2847:29]
  wire [31:0] _GEN_1062 = _T_105 & LUT_stack_io_pop_16 ? 32'h0 : _GEN_1023; // @[stackmanage_35.scala 2778:69 stackmanage_35.scala 2848:28]
  wire [31:0] _GEN_1063 = _T_105 & LUT_stack_io_pop_15 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 2707:69 stackmanage_35.scala 2708:29]
  wire [31:0] _GEN_1064 = _T_105 & LUT_stack_io_pop_15 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 2707:69 stackmanage_35.scala 2709:28]
  wire [31:0] _GEN_1066 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1024; // @[stackmanage_35.scala 2707:69 stackmanage_35.scala 2740:29]
  wire [31:0] _GEN_1067 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1025; // @[stackmanage_35.scala 2707:69 stackmanage_35.scala 2741:28]
  wire [31:0] _GEN_1068 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1027; // @[stackmanage_35.scala 2707:69 stackmanage_35.scala 2742:29]
  wire [31:0] _GEN_1069 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1028; // @[stackmanage_35.scala 2707:69 stackmanage_35.scala 2743:28]
  wire [31:0] _GEN_1070 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1029; // @[stackmanage_35.scala 2707:69 stackmanage_35.scala 2744:29]
  wire [31:0] _GEN_1071 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1030; // @[stackmanage_35.scala 2707:69 stackmanage_35.scala 2745:28]
  wire [31:0] _GEN_1072 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1031; // @[stackmanage_35.scala 2707:69 stackmanage_35.scala 2746:29]
  wire [31:0] _GEN_1073 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1032; // @[stackmanage_35.scala 2707:69 stackmanage_35.scala 2747:28]
  wire [31:0] _GEN_1074 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1033; // @[stackmanage_35.scala 2707:69 stackmanage_35.scala 2748:29]
  wire [31:0] _GEN_1075 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1034; // @[stackmanage_35.scala 2707:69 stackmanage_35.scala 2749:29]
  wire [31:0] _GEN_1076 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1035; // @[stackmanage_35.scala 2707:69 stackmanage_35.scala 2750:29]
  wire [31:0] _GEN_1077 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1036; // @[stackmanage_35.scala 2707:69 stackmanage_35.scala 2751:28]
  wire [31:0] _GEN_1078 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1037; // @[stackmanage_35.scala 2707:69 stackmanage_35.scala 2752:29]
  wire [31:0] _GEN_1079 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1038; // @[stackmanage_35.scala 2707:69 stackmanage_35.scala 2753:28]
  wire [31:0] _GEN_1080 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1039; // @[stackmanage_35.scala 2707:69 stackmanage_35.scala 2754:29]
  wire [31:0] _GEN_1081 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1040; // @[stackmanage_35.scala 2707:69 stackmanage_35.scala 2755:28]
  wire [31:0] _GEN_1082 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1041; // @[stackmanage_35.scala 2707:69 stackmanage_35.scala 2756:29]
  wire [31:0] _GEN_1083 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1042; // @[stackmanage_35.scala 2707:69 stackmanage_35.scala 2757:28]
  wire [31:0] _GEN_1084 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1043; // @[stackmanage_35.scala 2707:69 stackmanage_35.scala 2758:29]
  wire [31:0] _GEN_1085 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1044; // @[stackmanage_35.scala 2707:69 stackmanage_35.scala 2759:28]
  wire [31:0] _GEN_1086 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1045; // @[stackmanage_35.scala 2707:69 stackmanage_35.scala 2760:29]
  wire [31:0] _GEN_1087 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1046; // @[stackmanage_35.scala 2707:69 stackmanage_35.scala 2761:28]
  wire [31:0] _GEN_1088 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1047; // @[stackmanage_35.scala 2707:69 stackmanage_35.scala 2762:29]
  wire [31:0] _GEN_1089 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1048; // @[stackmanage_35.scala 2707:69 stackmanage_35.scala 2763:28]
  wire [31:0] _GEN_1090 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1049; // @[stackmanage_35.scala 2707:69 stackmanage_35.scala 2764:29]
  wire [31:0] _GEN_1091 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1050; // @[stackmanage_35.scala 2707:69 stackmanage_35.scala 2765:28]
  wire [31:0] _GEN_1092 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1051; // @[stackmanage_35.scala 2707:69 stackmanage_35.scala 2766:29]
  wire [31:0] _GEN_1093 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1052; // @[stackmanage_35.scala 2707:69 stackmanage_35.scala 2767:28]
  wire [31:0] _GEN_1094 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1053; // @[stackmanage_35.scala 2707:69 stackmanage_35.scala 2768:29]
  wire [31:0] _GEN_1095 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1054; // @[stackmanage_35.scala 2707:69 stackmanage_35.scala 2769:29]
  wire [31:0] _GEN_1096 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1055; // @[stackmanage_35.scala 2707:69 stackmanage_35.scala 2770:29]
  wire [31:0] _GEN_1097 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1056; // @[stackmanage_35.scala 2707:69 stackmanage_35.scala 2771:28]
  wire [31:0] _GEN_1098 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1057; // @[stackmanage_35.scala 2707:69 stackmanage_35.scala 2772:29]
  wire [31:0] _GEN_1099 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1058; // @[stackmanage_35.scala 2707:69 stackmanage_35.scala 2773:28]
  wire [31:0] _GEN_1100 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1059; // @[stackmanage_35.scala 2707:69 stackmanage_35.scala 2774:29]
  wire [31:0] _GEN_1101 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1060; // @[stackmanage_35.scala 2707:69 stackmanage_35.scala 2775:28]
  wire [31:0] _GEN_1102 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1061; // @[stackmanage_35.scala 2707:69 stackmanage_35.scala 2776:29]
  wire [31:0] _GEN_1103 = _T_105 & LUT_stack_io_pop_15 ? 32'h0 : _GEN_1062; // @[stackmanage_35.scala 2707:69 stackmanage_35.scala 2777:28]
  wire [31:0] _GEN_1104 = _T_105 & LUT_stack_io_pop_14 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 2636:69 stackmanage_35.scala 2637:29]
  wire [31:0] _GEN_1105 = _T_105 & LUT_stack_io_pop_14 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 2636:69 stackmanage_35.scala 2638:28]
  wire [31:0] _GEN_1107 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1063; // @[stackmanage_35.scala 2636:69 stackmanage_35.scala 2667:29]
  wire [31:0] _GEN_1108 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1064; // @[stackmanage_35.scala 2636:69 stackmanage_35.scala 2668:28]
  wire [31:0] _GEN_1109 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1066; // @[stackmanage_35.scala 2636:69 stackmanage_35.scala 2669:29]
  wire [31:0] _GEN_1110 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1067; // @[stackmanage_35.scala 2636:69 stackmanage_35.scala 2670:28]
  wire [31:0] _GEN_1111 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1068; // @[stackmanage_35.scala 2636:69 stackmanage_35.scala 2671:29]
  wire [31:0] _GEN_1112 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1069; // @[stackmanage_35.scala 2636:69 stackmanage_35.scala 2672:28]
  wire [31:0] _GEN_1113 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1070; // @[stackmanage_35.scala 2636:69 stackmanage_35.scala 2673:29]
  wire [31:0] _GEN_1114 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1071; // @[stackmanage_35.scala 2636:69 stackmanage_35.scala 2674:28]
  wire [31:0] _GEN_1115 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1072; // @[stackmanage_35.scala 2636:69 stackmanage_35.scala 2675:29]
  wire [31:0] _GEN_1116 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1073; // @[stackmanage_35.scala 2636:69 stackmanage_35.scala 2676:28]
  wire [31:0] _GEN_1117 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1074; // @[stackmanage_35.scala 2636:69 stackmanage_35.scala 2677:29]
  wire [31:0] _GEN_1118 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1075; // @[stackmanage_35.scala 2636:69 stackmanage_35.scala 2678:29]
  wire [31:0] _GEN_1119 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1076; // @[stackmanage_35.scala 2636:69 stackmanage_35.scala 2679:29]
  wire [31:0] _GEN_1120 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1077; // @[stackmanage_35.scala 2636:69 stackmanage_35.scala 2680:28]
  wire [31:0] _GEN_1121 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1078; // @[stackmanage_35.scala 2636:69 stackmanage_35.scala 2681:29]
  wire [31:0] _GEN_1122 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1079; // @[stackmanage_35.scala 2636:69 stackmanage_35.scala 2682:28]
  wire [31:0] _GEN_1123 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1080; // @[stackmanage_35.scala 2636:69 stackmanage_35.scala 2683:29]
  wire [31:0] _GEN_1124 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1081; // @[stackmanage_35.scala 2636:69 stackmanage_35.scala 2684:28]
  wire [31:0] _GEN_1125 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1082; // @[stackmanage_35.scala 2636:69 stackmanage_35.scala 2685:29]
  wire [31:0] _GEN_1126 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1083; // @[stackmanage_35.scala 2636:69 stackmanage_35.scala 2686:28]
  wire [31:0] _GEN_1127 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1084; // @[stackmanage_35.scala 2636:69 stackmanage_35.scala 2687:29]
  wire [31:0] _GEN_1128 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1085; // @[stackmanage_35.scala 2636:69 stackmanage_35.scala 2688:28]
  wire [31:0] _GEN_1129 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1086; // @[stackmanage_35.scala 2636:69 stackmanage_35.scala 2689:29]
  wire [31:0] _GEN_1130 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1087; // @[stackmanage_35.scala 2636:69 stackmanage_35.scala 2690:28]
  wire [31:0] _GEN_1131 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1088; // @[stackmanage_35.scala 2636:69 stackmanage_35.scala 2691:29]
  wire [31:0] _GEN_1132 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1089; // @[stackmanage_35.scala 2636:69 stackmanage_35.scala 2692:28]
  wire [31:0] _GEN_1133 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1090; // @[stackmanage_35.scala 2636:69 stackmanage_35.scala 2693:29]
  wire [31:0] _GEN_1134 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1091; // @[stackmanage_35.scala 2636:69 stackmanage_35.scala 2694:28]
  wire [31:0] _GEN_1135 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1092; // @[stackmanage_35.scala 2636:69 stackmanage_35.scala 2695:29]
  wire [31:0] _GEN_1136 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1093; // @[stackmanage_35.scala 2636:69 stackmanage_35.scala 2696:28]
  wire [31:0] _GEN_1137 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1094; // @[stackmanage_35.scala 2636:69 stackmanage_35.scala 2697:29]
  wire [31:0] _GEN_1138 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1095; // @[stackmanage_35.scala 2636:69 stackmanage_35.scala 2698:29]
  wire [31:0] _GEN_1139 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1096; // @[stackmanage_35.scala 2636:69 stackmanage_35.scala 2699:29]
  wire [31:0] _GEN_1140 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1097; // @[stackmanage_35.scala 2636:69 stackmanage_35.scala 2700:28]
  wire [31:0] _GEN_1141 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1098; // @[stackmanage_35.scala 2636:69 stackmanage_35.scala 2701:29]
  wire [31:0] _GEN_1142 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1099; // @[stackmanage_35.scala 2636:69 stackmanage_35.scala 2702:28]
  wire [31:0] _GEN_1143 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1100; // @[stackmanage_35.scala 2636:69 stackmanage_35.scala 2703:29]
  wire [31:0] _GEN_1144 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1101; // @[stackmanage_35.scala 2636:69 stackmanage_35.scala 2704:28]
  wire [31:0] _GEN_1145 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1102; // @[stackmanage_35.scala 2636:69 stackmanage_35.scala 2705:29]
  wire [31:0] _GEN_1146 = _T_105 & LUT_stack_io_pop_14 ? 32'h0 : _GEN_1103; // @[stackmanage_35.scala 2636:69 stackmanage_35.scala 2706:28]
  wire [31:0] _GEN_1147 = _T_105 & LUT_stack_io_pop_13 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2566:29]
  wire [31:0] _GEN_1148 = _T_105 & LUT_stack_io_pop_13 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2567:28]
  wire [31:0] _GEN_1150 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1104; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2594:29]
  wire [31:0] _GEN_1151 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1105; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2595:28]
  wire [31:0] _GEN_1152 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1107; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2596:29]
  wire [31:0] _GEN_1153 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1108; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2597:28]
  wire [31:0] _GEN_1154 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1109; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2598:29]
  wire [31:0] _GEN_1155 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1110; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2599:28]
  wire [31:0] _GEN_1156 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1111; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2600:29]
  wire [31:0] _GEN_1157 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1112; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2601:28]
  wire [31:0] _GEN_1158 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1113; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2602:29]
  wire [31:0] _GEN_1159 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1114; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2603:28]
  wire [31:0] _GEN_1160 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1115; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2604:29]
  wire [31:0] _GEN_1161 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1116; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2605:28]
  wire [31:0] _GEN_1162 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1117; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2606:29]
  wire [31:0] _GEN_1163 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1118; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2607:29]
  wire [31:0] _GEN_1164 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1119; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2608:29]
  wire [31:0] _GEN_1165 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1120; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2609:28]
  wire [31:0] _GEN_1166 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1121; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2610:29]
  wire [31:0] _GEN_1167 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1122; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2611:28]
  wire [31:0] _GEN_1168 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1123; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2612:29]
  wire [31:0] _GEN_1169 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1124; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2613:28]
  wire [31:0] _GEN_1170 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1125; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2614:29]
  wire [31:0] _GEN_1171 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1126; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2615:28]
  wire [31:0] _GEN_1172 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1127; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2616:29]
  wire [31:0] _GEN_1173 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1128; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2617:28]
  wire [31:0] _GEN_1174 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1129; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2618:29]
  wire [31:0] _GEN_1175 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1130; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2619:28]
  wire [31:0] _GEN_1176 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1131; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2620:29]
  wire [31:0] _GEN_1177 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1132; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2621:28]
  wire [31:0] _GEN_1178 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1133; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2622:29]
  wire [31:0] _GEN_1179 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1134; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2623:28]
  wire [31:0] _GEN_1180 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1135; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2624:29]
  wire [31:0] _GEN_1181 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1136; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2625:28]
  wire [31:0] _GEN_1182 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1137; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2626:29]
  wire [31:0] _GEN_1183 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1138; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2627:29]
  wire [31:0] _GEN_1184 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1139; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2628:29]
  wire [31:0] _GEN_1185 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1140; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2629:28]
  wire [31:0] _GEN_1186 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1141; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2630:29]
  wire [31:0] _GEN_1187 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1142; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2631:28]
  wire [31:0] _GEN_1188 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1143; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2632:29]
  wire [31:0] _GEN_1189 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1144; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2633:28]
  wire [31:0] _GEN_1190 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1145; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2634:29]
  wire [31:0] _GEN_1191 = _T_105 & LUT_stack_io_pop_13 ? 32'h0 : _GEN_1146; // @[stackmanage_35.scala 2565:69 stackmanage_35.scala 2635:28]
  wire [31:0] _GEN_1192 = _T_105 & LUT_stack_io_pop_12 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2495:29]
  wire [31:0] _GEN_1193 = _T_105 & LUT_stack_io_pop_12 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2496:28]
  wire [31:0] _GEN_1195 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1147; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2521:29]
  wire [31:0] _GEN_1196 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1148; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2522:28]
  wire [31:0] _GEN_1197 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1150; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2523:29]
  wire [31:0] _GEN_1198 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1151; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2524:28]
  wire [31:0] _GEN_1199 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1152; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2525:29]
  wire [31:0] _GEN_1200 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1153; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2526:28]
  wire [31:0] _GEN_1201 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1154; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2527:29]
  wire [31:0] _GEN_1202 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1155; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2528:28]
  wire [31:0] _GEN_1203 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1156; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2529:29]
  wire [31:0] _GEN_1204 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1157; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2530:28]
  wire [31:0] _GEN_1205 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1158; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2531:29]
  wire [31:0] _GEN_1206 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1159; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2532:28]
  wire [31:0] _GEN_1207 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1160; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2533:29]
  wire [31:0] _GEN_1208 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1161; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2534:28]
  wire [31:0] _GEN_1209 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1162; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2535:29]
  wire [31:0] _GEN_1210 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1163; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2536:29]
  wire [31:0] _GEN_1211 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1164; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2537:29]
  wire [31:0] _GEN_1212 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1165; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2538:28]
  wire [31:0] _GEN_1213 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1166; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2539:29]
  wire [31:0] _GEN_1214 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1167; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2540:28]
  wire [31:0] _GEN_1215 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1168; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2541:29]
  wire [31:0] _GEN_1216 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1169; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2542:28]
  wire [31:0] _GEN_1217 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1170; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2543:29]
  wire [31:0] _GEN_1218 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1171; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2544:28]
  wire [31:0] _GEN_1219 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1172; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2545:29]
  wire [31:0] _GEN_1220 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1173; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2546:28]
  wire [31:0] _GEN_1221 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1174; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2547:29]
  wire [31:0] _GEN_1222 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1175; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2548:28]
  wire [31:0] _GEN_1223 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1176; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2549:29]
  wire [31:0] _GEN_1224 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1177; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2550:28]
  wire [31:0] _GEN_1225 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1178; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2551:29]
  wire [31:0] _GEN_1226 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1179; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2552:28]
  wire [31:0] _GEN_1227 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1180; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2553:29]
  wire [31:0] _GEN_1228 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1181; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2554:28]
  wire [31:0] _GEN_1229 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1182; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2555:29]
  wire [31:0] _GEN_1230 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1183; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2556:29]
  wire [31:0] _GEN_1231 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1184; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2557:29]
  wire [31:0] _GEN_1232 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1185; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2558:28]
  wire [31:0] _GEN_1233 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1186; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2559:29]
  wire [31:0] _GEN_1234 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1187; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2560:28]
  wire [31:0] _GEN_1235 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1188; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2561:29]
  wire [31:0] _GEN_1236 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1189; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2562:28]
  wire [31:0] _GEN_1237 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1190; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2563:29]
  wire [31:0] _GEN_1238 = _T_105 & LUT_stack_io_pop_12 ? 32'h0 : _GEN_1191; // @[stackmanage_35.scala 2494:69 stackmanage_35.scala 2564:28]
  wire [31:0] _GEN_1239 = _T_105 & LUT_stack_io_pop_11 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2424:29]
  wire [31:0] _GEN_1240 = _T_105 & LUT_stack_io_pop_11 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2425:28]
  wire [31:0] _GEN_1242 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1192; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2448:29]
  wire [31:0] _GEN_1243 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1193; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2449:28]
  wire [31:0] _GEN_1244 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1195; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2450:29]
  wire [31:0] _GEN_1245 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1196; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2451:28]
  wire [31:0] _GEN_1246 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1197; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2452:29]
  wire [31:0] _GEN_1247 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1198; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2453:28]
  wire [31:0] _GEN_1248 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1199; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2454:29]
  wire [31:0] _GEN_1249 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1200; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2455:28]
  wire [31:0] _GEN_1250 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1201; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2456:29]
  wire [31:0] _GEN_1251 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1202; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2457:28]
  wire [31:0] _GEN_1252 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1203; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2458:29]
  wire [31:0] _GEN_1253 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1204; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2459:28]
  wire [31:0] _GEN_1254 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1205; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2460:29]
  wire [31:0] _GEN_1255 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1206; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2461:28]
  wire [31:0] _GEN_1256 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1207; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2462:29]
  wire [31:0] _GEN_1257 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1208; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2463:28]
  wire [31:0] _GEN_1258 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1209; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2464:29]
  wire [31:0] _GEN_1259 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1210; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2465:29]
  wire [31:0] _GEN_1260 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1211; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2466:29]
  wire [31:0] _GEN_1261 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1212; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2467:28]
  wire [31:0] _GEN_1262 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1213; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2468:29]
  wire [31:0] _GEN_1263 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1214; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2469:28]
  wire [31:0] _GEN_1264 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1215; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2470:29]
  wire [31:0] _GEN_1265 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1216; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2471:28]
  wire [31:0] _GEN_1266 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1217; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2472:29]
  wire [31:0] _GEN_1267 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1218; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2473:28]
  wire [31:0] _GEN_1268 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1219; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2474:29]
  wire [31:0] _GEN_1269 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1220; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2475:28]
  wire [31:0] _GEN_1270 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1221; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2476:29]
  wire [31:0] _GEN_1271 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1222; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2477:28]
  wire [31:0] _GEN_1272 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1223; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2478:29]
  wire [31:0] _GEN_1273 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1224; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2479:28]
  wire [31:0] _GEN_1274 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1225; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2480:29]
  wire [31:0] _GEN_1275 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1226; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2481:28]
  wire [31:0] _GEN_1276 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1227; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2482:29]
  wire [31:0] _GEN_1277 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1228; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2483:28]
  wire [31:0] _GEN_1278 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1229; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2484:29]
  wire [31:0] _GEN_1279 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1230; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2485:29]
  wire [31:0] _GEN_1280 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1231; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2486:29]
  wire [31:0] _GEN_1281 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1232; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2487:28]
  wire [31:0] _GEN_1282 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1233; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2488:29]
  wire [31:0] _GEN_1283 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1234; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2489:28]
  wire [31:0] _GEN_1284 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1235; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2490:29]
  wire [31:0] _GEN_1285 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1236; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2491:28]
  wire [31:0] _GEN_1286 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1237; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2492:29]
  wire [31:0] _GEN_1287 = _T_105 & LUT_stack_io_pop_11 ? 32'h0 : _GEN_1238; // @[stackmanage_35.scala 2423:69 stackmanage_35.scala 2493:28]
  wire [31:0] _GEN_1288 = _T_105 & LUT_stack_io_pop_10 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2353:29]
  wire [31:0] _GEN_1289 = _T_105 & LUT_stack_io_pop_10 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2354:28]
  wire [31:0] _GEN_1291 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1239; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2375:29]
  wire [31:0] _GEN_1292 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1240; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2376:28]
  wire [31:0] _GEN_1293 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1242; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2377:29]
  wire [31:0] _GEN_1294 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1243; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2378:28]
  wire [31:0] _GEN_1295 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1244; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2379:29]
  wire [31:0] _GEN_1296 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1245; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2380:28]
  wire [31:0] _GEN_1297 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1246; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2381:29]
  wire [31:0] _GEN_1298 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1247; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2382:28]
  wire [31:0] _GEN_1299 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1248; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2383:29]
  wire [31:0] _GEN_1300 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1249; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2384:28]
  wire [31:0] _GEN_1301 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1250; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2385:29]
  wire [31:0] _GEN_1302 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1251; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2386:28]
  wire [31:0] _GEN_1303 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1252; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2387:29]
  wire [31:0] _GEN_1304 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1253; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2388:28]
  wire [31:0] _GEN_1305 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1254; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2389:29]
  wire [31:0] _GEN_1306 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1255; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2390:28]
  wire [31:0] _GEN_1307 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1256; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2391:29]
  wire [31:0] _GEN_1308 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1257; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2392:28]
  wire [31:0] _GEN_1309 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1258; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2393:29]
  wire [31:0] _GEN_1310 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1259; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2394:29]
  wire [31:0] _GEN_1311 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1260; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2395:29]
  wire [31:0] _GEN_1312 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1261; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2396:28]
  wire [31:0] _GEN_1313 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1262; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2397:29]
  wire [31:0] _GEN_1314 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1263; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2398:28]
  wire [31:0] _GEN_1315 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1264; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2399:29]
  wire [31:0] _GEN_1316 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1265; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2400:28]
  wire [31:0] _GEN_1317 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1266; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2401:29]
  wire [31:0] _GEN_1318 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1267; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2402:28]
  wire [31:0] _GEN_1319 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1268; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2403:29]
  wire [31:0] _GEN_1320 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1269; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2404:28]
  wire [31:0] _GEN_1321 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1270; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2405:29]
  wire [31:0] _GEN_1322 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1271; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2406:28]
  wire [31:0] _GEN_1323 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1272; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2407:29]
  wire [31:0] _GEN_1324 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1273; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2408:28]
  wire [31:0] _GEN_1325 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1274; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2409:29]
  wire [31:0] _GEN_1326 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1275; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2410:28]
  wire [31:0] _GEN_1327 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1276; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2411:29]
  wire [31:0] _GEN_1328 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1277; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2412:28]
  wire [31:0] _GEN_1329 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1278; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2413:29]
  wire [31:0] _GEN_1330 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1279; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2414:29]
  wire [31:0] _GEN_1331 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1280; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2415:29]
  wire [31:0] _GEN_1332 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1281; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2416:28]
  wire [31:0] _GEN_1333 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1282; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2417:29]
  wire [31:0] _GEN_1334 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1283; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2418:28]
  wire [31:0] _GEN_1335 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1284; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2419:29]
  wire [31:0] _GEN_1336 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1285; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2420:28]
  wire [31:0] _GEN_1337 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1286; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2421:29]
  wire [31:0] _GEN_1338 = _T_105 & LUT_stack_io_pop_10 ? 32'h0 : _GEN_1287; // @[stackmanage_35.scala 2352:69 stackmanage_35.scala 2422:28]
  wire [31:0] _GEN_1339 = _T_105 & LUT_stack_io_pop_9 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2282:28]
  wire [31:0] _GEN_1340 = _T_105 & LUT_stack_io_pop_9 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2283:27]
  wire [31:0] _GEN_1342 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1288; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2302:29]
  wire [31:0] _GEN_1343 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1289; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2303:29]
  wire [31:0] _GEN_1344 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1291; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2304:29]
  wire [31:0] _GEN_1345 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1292; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2305:28]
  wire [31:0] _GEN_1346 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1293; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2306:29]
  wire [31:0] _GEN_1347 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1294; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2307:28]
  wire [31:0] _GEN_1348 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1295; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2308:29]
  wire [31:0] _GEN_1349 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1296; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2309:28]
  wire [31:0] _GEN_1350 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1297; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2310:29]
  wire [31:0] _GEN_1351 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1298; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2311:28]
  wire [31:0] _GEN_1352 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1299; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2312:29]
  wire [31:0] _GEN_1353 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1300; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2313:28]
  wire [31:0] _GEN_1354 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1301; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2314:29]
  wire [31:0] _GEN_1355 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1302; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2315:28]
  wire [31:0] _GEN_1356 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1303; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2316:29]
  wire [31:0] _GEN_1357 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1304; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2317:28]
  wire [31:0] _GEN_1358 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1305; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2318:29]
  wire [31:0] _GEN_1359 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1306; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2319:28]
  wire [31:0] _GEN_1360 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1307; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2320:29]
  wire [31:0] _GEN_1361 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1308; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2321:28]
  wire [31:0] _GEN_1362 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1309; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2322:29]
  wire [31:0] _GEN_1363 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1310; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2323:29]
  wire [31:0] _GEN_1364 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1311; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2324:29]
  wire [31:0] _GEN_1365 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1312; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2325:28]
  wire [31:0] _GEN_1366 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1313; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2326:29]
  wire [31:0] _GEN_1367 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1314; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2327:28]
  wire [31:0] _GEN_1368 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1315; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2328:29]
  wire [31:0] _GEN_1369 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1316; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2329:28]
  wire [31:0] _GEN_1370 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1317; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2330:29]
  wire [31:0] _GEN_1371 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1318; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2331:28]
  wire [31:0] _GEN_1372 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1319; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2332:29]
  wire [31:0] _GEN_1373 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1320; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2333:28]
  wire [31:0] _GEN_1374 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1321; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2334:29]
  wire [31:0] _GEN_1375 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1322; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2335:28]
  wire [31:0] _GEN_1376 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1323; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2336:29]
  wire [31:0] _GEN_1377 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1324; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2337:28]
  wire [31:0] _GEN_1378 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1325; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2338:29]
  wire [31:0] _GEN_1379 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1326; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2339:28]
  wire [31:0] _GEN_1380 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1327; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2340:29]
  wire [31:0] _GEN_1381 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1328; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2341:28]
  wire [31:0] _GEN_1382 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1329; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2342:29]
  wire [31:0] _GEN_1383 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1330; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2343:29]
  wire [31:0] _GEN_1384 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1331; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2344:29]
  wire [31:0] _GEN_1385 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1332; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2345:28]
  wire [31:0] _GEN_1386 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1333; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2346:29]
  wire [31:0] _GEN_1387 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1334; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2347:28]
  wire [31:0] _GEN_1388 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1335; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2348:29]
  wire [31:0] _GEN_1389 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1336; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2349:28]
  wire [31:0] _GEN_1390 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1337; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2350:29]
  wire [31:0] _GEN_1391 = _T_105 & LUT_stack_io_pop_9 ? 32'h0 : _GEN_1338; // @[stackmanage_35.scala 2281:68 stackmanage_35.scala 2351:28]
  wire [31:0] _GEN_1392 = _T_105 & LUT_stack_io_pop_8 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2211:28]
  wire [31:0] _GEN_1393 = _T_105 & LUT_stack_io_pop_8 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2212:27]
  wire [31:0] _GEN_1395 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1339; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2229:28]
  wire [31:0] _GEN_1396 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1340; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2230:27]
  wire [31:0] _GEN_1397 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1342; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2231:29]
  wire [31:0] _GEN_1398 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1343; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2232:29]
  wire [31:0] _GEN_1399 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1344; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2233:29]
  wire [31:0] _GEN_1400 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1345; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2234:28]
  wire [31:0] _GEN_1401 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1346; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2235:29]
  wire [31:0] _GEN_1402 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1347; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2236:28]
  wire [31:0] _GEN_1403 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1348; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2237:29]
  wire [31:0] _GEN_1404 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1349; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2238:28]
  wire [31:0] _GEN_1405 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1350; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2239:29]
  wire [31:0] _GEN_1406 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1351; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2240:28]
  wire [31:0] _GEN_1407 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1352; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2241:29]
  wire [31:0] _GEN_1408 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1353; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2242:28]
  wire [31:0] _GEN_1409 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1354; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2243:29]
  wire [31:0] _GEN_1410 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1355; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2244:28]
  wire [31:0] _GEN_1411 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1356; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2245:29]
  wire [31:0] _GEN_1412 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1357; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2246:28]
  wire [31:0] _GEN_1413 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1358; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2247:29]
  wire [31:0] _GEN_1414 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1359; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2248:28]
  wire [31:0] _GEN_1415 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1360; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2249:29]
  wire [31:0] _GEN_1416 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1361; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2250:28]
  wire [31:0] _GEN_1417 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1362; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2251:29]
  wire [31:0] _GEN_1418 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1363; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2252:29]
  wire [31:0] _GEN_1419 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1364; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2253:29]
  wire [31:0] _GEN_1420 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1365; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2254:28]
  wire [31:0] _GEN_1421 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1366; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2255:29]
  wire [31:0] _GEN_1422 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1367; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2256:28]
  wire [31:0] _GEN_1423 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1368; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2257:29]
  wire [31:0] _GEN_1424 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1369; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2258:28]
  wire [31:0] _GEN_1425 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1370; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2259:29]
  wire [31:0] _GEN_1426 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1371; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2260:28]
  wire [31:0] _GEN_1427 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1372; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2261:29]
  wire [31:0] _GEN_1428 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1373; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2262:28]
  wire [31:0] _GEN_1429 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1374; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2263:29]
  wire [31:0] _GEN_1430 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1375; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2264:28]
  wire [31:0] _GEN_1431 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1376; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2265:29]
  wire [31:0] _GEN_1432 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1377; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2266:28]
  wire [31:0] _GEN_1433 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1378; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2267:29]
  wire [31:0] _GEN_1434 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1379; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2268:28]
  wire [31:0] _GEN_1435 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1380; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2269:29]
  wire [31:0] _GEN_1436 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1381; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2270:28]
  wire [31:0] _GEN_1437 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1382; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2271:29]
  wire [31:0] _GEN_1438 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1383; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2272:29]
  wire [31:0] _GEN_1439 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1384; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2273:29]
  wire [31:0] _GEN_1440 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1385; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2274:28]
  wire [31:0] _GEN_1441 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1386; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2275:29]
  wire [31:0] _GEN_1442 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1387; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2276:28]
  wire [31:0] _GEN_1443 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1388; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2277:29]
  wire [31:0] _GEN_1444 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1389; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2278:28]
  wire [31:0] _GEN_1445 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1390; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2279:29]
  wire [31:0] _GEN_1446 = _T_105 & LUT_stack_io_pop_8 ? 32'h0 : _GEN_1391; // @[stackmanage_35.scala 2210:68 stackmanage_35.scala 2280:28]
  wire [31:0] _GEN_1447 = _T_105 & LUT_stack_io_pop_7 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2140:28]
  wire [31:0] _GEN_1448 = _T_105 & LUT_stack_io_pop_7 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2141:27]
  wire [31:0] _GEN_1450 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1392; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2156:28]
  wire [31:0] _GEN_1451 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1393; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2157:27]
  wire [31:0] _GEN_1452 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1395; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2158:28]
  wire [31:0] _GEN_1453 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1396; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2159:27]
  wire [31:0] _GEN_1454 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1397; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2160:29]
  wire [31:0] _GEN_1455 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1398; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2161:29]
  wire [31:0] _GEN_1456 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1399; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2162:29]
  wire [31:0] _GEN_1457 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1400; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2163:28]
  wire [31:0] _GEN_1458 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1401; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2164:29]
  wire [31:0] _GEN_1459 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1402; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2165:28]
  wire [31:0] _GEN_1460 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1403; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2166:29]
  wire [31:0] _GEN_1461 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1404; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2167:28]
  wire [31:0] _GEN_1462 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1405; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2168:29]
  wire [31:0] _GEN_1463 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1406; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2169:28]
  wire [31:0] _GEN_1464 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1407; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2170:29]
  wire [31:0] _GEN_1465 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1408; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2171:28]
  wire [31:0] _GEN_1466 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1409; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2172:29]
  wire [31:0] _GEN_1467 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1410; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2173:28]
  wire [31:0] _GEN_1468 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1411; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2174:29]
  wire [31:0] _GEN_1469 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1412; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2175:28]
  wire [31:0] _GEN_1470 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1413; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2176:29]
  wire [31:0] _GEN_1471 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1414; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2177:28]
  wire [31:0] _GEN_1472 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1415; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2178:29]
  wire [31:0] _GEN_1473 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1416; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2179:28]
  wire [31:0] _GEN_1474 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1417; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2180:29]
  wire [31:0] _GEN_1475 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1418; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2181:29]
  wire [31:0] _GEN_1476 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1419; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2182:29]
  wire [31:0] _GEN_1477 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1420; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2183:28]
  wire [31:0] _GEN_1478 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1421; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2184:29]
  wire [31:0] _GEN_1479 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1422; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2185:28]
  wire [31:0] _GEN_1480 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1423; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2186:29]
  wire [31:0] _GEN_1481 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1424; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2187:28]
  wire [31:0] _GEN_1482 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1425; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2188:29]
  wire [31:0] _GEN_1483 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1426; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2189:28]
  wire [31:0] _GEN_1484 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1427; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2190:29]
  wire [31:0] _GEN_1485 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1428; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2191:28]
  wire [31:0] _GEN_1486 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1429; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2192:29]
  wire [31:0] _GEN_1487 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1430; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2193:28]
  wire [31:0] _GEN_1488 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1431; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2194:29]
  wire [31:0] _GEN_1489 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1432; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2195:28]
  wire [31:0] _GEN_1490 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1433; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2196:29]
  wire [31:0] _GEN_1491 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1434; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2197:28]
  wire [31:0] _GEN_1492 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1435; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2198:29]
  wire [31:0] _GEN_1493 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1436; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2199:28]
  wire [31:0] _GEN_1494 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1437; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2200:29]
  wire [31:0] _GEN_1495 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1438; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2201:29]
  wire [31:0] _GEN_1496 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1439; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2202:29]
  wire [31:0] _GEN_1497 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1440; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2203:28]
  wire [31:0] _GEN_1498 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1441; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2204:29]
  wire [31:0] _GEN_1499 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1442; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2205:28]
  wire [31:0] _GEN_1500 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1443; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2206:29]
  wire [31:0] _GEN_1501 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1444; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2207:28]
  wire [31:0] _GEN_1502 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1445; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2208:29]
  wire [31:0] _GEN_1503 = _T_105 & LUT_stack_io_pop_7 ? 32'h0 : _GEN_1446; // @[stackmanage_35.scala 2139:68 stackmanage_35.scala 2209:28]
  wire [31:0] _GEN_1504 = _T_105 & LUT_stack_io_pop_6 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2069:28]
  wire [31:0] _GEN_1505 = _T_105 & LUT_stack_io_pop_6 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2070:27]
  wire [31:0] _GEN_1507 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1447; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2083:28]
  wire [31:0] _GEN_1508 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1448; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2084:27]
  wire [31:0] _GEN_1509 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1450; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2085:28]
  wire [31:0] _GEN_1510 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1451; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2086:27]
  wire [31:0] _GEN_1511 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1452; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2087:28]
  wire [31:0] _GEN_1512 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1453; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2088:27]
  wire [31:0] _GEN_1513 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1454; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2089:29]
  wire [31:0] _GEN_1514 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1455; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2090:29]
  wire [31:0] _GEN_1515 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1456; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2091:29]
  wire [31:0] _GEN_1516 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1457; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2092:28]
  wire [31:0] _GEN_1517 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1458; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2093:29]
  wire [31:0] _GEN_1518 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1459; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2094:28]
  wire [31:0] _GEN_1519 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1460; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2095:29]
  wire [31:0] _GEN_1520 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1461; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2096:28]
  wire [31:0] _GEN_1521 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1462; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2097:29]
  wire [31:0] _GEN_1522 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1463; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2098:28]
  wire [31:0] _GEN_1523 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1464; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2099:29]
  wire [31:0] _GEN_1524 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1465; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2100:28]
  wire [31:0] _GEN_1525 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1466; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2101:29]
  wire [31:0] _GEN_1526 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1467; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2102:28]
  wire [31:0] _GEN_1527 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1468; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2103:29]
  wire [31:0] _GEN_1528 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1469; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2104:28]
  wire [31:0] _GEN_1529 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1470; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2105:29]
  wire [31:0] _GEN_1530 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1471; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2106:28]
  wire [31:0] _GEN_1531 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1472; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2107:29]
  wire [31:0] _GEN_1532 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1473; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2108:28]
  wire [31:0] _GEN_1533 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1474; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2109:29]
  wire [31:0] _GEN_1534 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1475; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2110:29]
  wire [31:0] _GEN_1535 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1476; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2111:29]
  wire [31:0] _GEN_1536 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1477; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2112:28]
  wire [31:0] _GEN_1537 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1478; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2113:29]
  wire [31:0] _GEN_1538 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1479; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2114:28]
  wire [31:0] _GEN_1539 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1480; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2115:29]
  wire [31:0] _GEN_1540 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1481; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2116:28]
  wire [31:0] _GEN_1541 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1482; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2117:29]
  wire [31:0] _GEN_1542 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1483; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2118:28]
  wire [31:0] _GEN_1543 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1484; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2119:29]
  wire [31:0] _GEN_1544 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1485; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2120:28]
  wire [31:0] _GEN_1545 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1486; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2121:29]
  wire [31:0] _GEN_1546 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1487; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2122:28]
  wire [31:0] _GEN_1547 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1488; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2123:29]
  wire [31:0] _GEN_1548 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1489; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2124:28]
  wire [31:0] _GEN_1549 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1490; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2125:29]
  wire [31:0] _GEN_1550 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1491; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2126:28]
  wire [31:0] _GEN_1551 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1492; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2127:29]
  wire [31:0] _GEN_1552 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1493; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2128:28]
  wire [31:0] _GEN_1553 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1494; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2129:29]
  wire [31:0] _GEN_1554 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1495; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2130:29]
  wire [31:0] _GEN_1555 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1496; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2131:29]
  wire [31:0] _GEN_1556 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1497; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2132:28]
  wire [31:0] _GEN_1557 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1498; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2133:29]
  wire [31:0] _GEN_1558 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1499; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2134:28]
  wire [31:0] _GEN_1559 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1500; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2135:29]
  wire [31:0] _GEN_1560 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1501; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2136:28]
  wire [31:0] _GEN_1561 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1502; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2137:29]
  wire [31:0] _GEN_1562 = _T_105 & LUT_stack_io_pop_6 ? 32'h0 : _GEN_1503; // @[stackmanage_35.scala 2068:68 stackmanage_35.scala 2138:28]
  wire [31:0] _GEN_1563 = _T_105 & LUT_stack_io_pop_5 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 1998:28]
  wire [31:0] _GEN_1564 = _T_105 & LUT_stack_io_pop_5 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 1999:27]
  wire [31:0] _GEN_1566 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1504; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2010:28]
  wire [31:0] _GEN_1567 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1505; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2011:27]
  wire [31:0] _GEN_1568 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1507; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2012:28]
  wire [31:0] _GEN_1569 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1508; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2013:27]
  wire [31:0] _GEN_1570 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1509; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2014:28]
  wire [31:0] _GEN_1571 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1510; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2015:27]
  wire [31:0] _GEN_1572 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1511; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2016:28]
  wire [31:0] _GEN_1573 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1512; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2017:27]
  wire [31:0] _GEN_1574 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1513; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2018:29]
  wire [31:0] _GEN_1575 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1514; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2019:29]
  wire [31:0] _GEN_1576 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1515; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2020:29]
  wire [31:0] _GEN_1577 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1516; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2021:28]
  wire [31:0] _GEN_1578 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1517; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2022:29]
  wire [31:0] _GEN_1579 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1518; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2023:28]
  wire [31:0] _GEN_1580 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1519; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2024:29]
  wire [31:0] _GEN_1581 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1520; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2025:28]
  wire [31:0] _GEN_1582 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1521; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2026:29]
  wire [31:0] _GEN_1583 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1522; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2027:28]
  wire [31:0] _GEN_1584 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1523; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2028:29]
  wire [31:0] _GEN_1585 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1524; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2029:28]
  wire [31:0] _GEN_1586 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1525; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2030:29]
  wire [31:0] _GEN_1587 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1526; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2031:28]
  wire [31:0] _GEN_1588 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1527; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2032:29]
  wire [31:0] _GEN_1589 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1528; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2033:28]
  wire [31:0] _GEN_1590 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1529; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2034:29]
  wire [31:0] _GEN_1591 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1530; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2035:28]
  wire [31:0] _GEN_1592 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1531; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2036:29]
  wire [31:0] _GEN_1593 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1532; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2037:28]
  wire [31:0] _GEN_1594 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1533; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2038:29]
  wire [31:0] _GEN_1595 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1534; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2039:29]
  wire [31:0] _GEN_1596 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1535; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2040:29]
  wire [31:0] _GEN_1597 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1536; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2041:28]
  wire [31:0] _GEN_1598 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1537; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2042:29]
  wire [31:0] _GEN_1599 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1538; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2043:28]
  wire [31:0] _GEN_1600 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1539; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2044:29]
  wire [31:0] _GEN_1601 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1540; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2045:28]
  wire [31:0] _GEN_1602 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1541; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2046:29]
  wire [31:0] _GEN_1603 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1542; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2047:28]
  wire [31:0] _GEN_1604 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1543; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2048:29]
  wire [31:0] _GEN_1605 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1544; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2049:28]
  wire [31:0] _GEN_1606 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1545; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2050:29]
  wire [31:0] _GEN_1607 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1546; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2051:28]
  wire [31:0] _GEN_1608 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1547; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2052:29]
  wire [31:0] _GEN_1609 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1548; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2053:28]
  wire [31:0] _GEN_1610 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1549; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2054:29]
  wire [31:0] _GEN_1611 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1550; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2055:28]
  wire [31:0] _GEN_1612 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1551; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2056:29]
  wire [31:0] _GEN_1613 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1552; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2057:28]
  wire [31:0] _GEN_1614 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1553; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2058:29]
  wire [31:0] _GEN_1615 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1554; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2059:29]
  wire [31:0] _GEN_1616 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1555; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2060:29]
  wire [31:0] _GEN_1617 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1556; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2061:28]
  wire [31:0] _GEN_1618 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1557; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2062:29]
  wire [31:0] _GEN_1619 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1558; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2063:28]
  wire [31:0] _GEN_1620 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1559; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2064:29]
  wire [31:0] _GEN_1621 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1560; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2065:28]
  wire [31:0] _GEN_1622 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1561; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2066:29]
  wire [31:0] _GEN_1623 = _T_105 & LUT_stack_io_pop_5 ? 32'h0 : _GEN_1562; // @[stackmanage_35.scala 1997:68 stackmanage_35.scala 2067:28]
  wire [31:0] _GEN_1624 = _T_105 & LUT_stack_io_pop_4 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1927:28]
  wire [31:0] _GEN_1625 = _T_105 & LUT_stack_io_pop_4 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1928:27]
  wire [31:0] _GEN_1627 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1563; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1937:28]
  wire [31:0] _GEN_1628 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1564; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1938:27]
  wire [31:0] _GEN_1629 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1566; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1939:28]
  wire [31:0] _GEN_1630 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1567; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1940:27]
  wire [31:0] _GEN_1631 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1568; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1941:28]
  wire [31:0] _GEN_1632 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1569; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1942:27]
  wire [31:0] _GEN_1633 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1570; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1943:28]
  wire [31:0] _GEN_1634 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1571; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1944:27]
  wire [31:0] _GEN_1635 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1572; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1945:28]
  wire [31:0] _GEN_1636 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1573; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1946:27]
  wire [31:0] _GEN_1637 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1574; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1947:29]
  wire [31:0] _GEN_1638 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1575; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1948:29]
  wire [31:0] _GEN_1639 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1576; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1949:29]
  wire [31:0] _GEN_1640 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1577; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1950:28]
  wire [31:0] _GEN_1641 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1578; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1951:29]
  wire [31:0] _GEN_1642 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1579; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1952:28]
  wire [31:0] _GEN_1643 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1580; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1953:29]
  wire [31:0] _GEN_1644 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1581; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1954:28]
  wire [31:0] _GEN_1645 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1582; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1955:29]
  wire [31:0] _GEN_1646 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1583; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1956:28]
  wire [31:0] _GEN_1647 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1584; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1957:29]
  wire [31:0] _GEN_1648 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1585; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1958:28]
  wire [31:0] _GEN_1649 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1586; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1959:29]
  wire [31:0] _GEN_1650 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1587; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1960:28]
  wire [31:0] _GEN_1651 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1588; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1961:29]
  wire [31:0] _GEN_1652 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1589; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1962:28]
  wire [31:0] _GEN_1653 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1590; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1963:29]
  wire [31:0] _GEN_1654 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1591; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1964:28]
  wire [31:0] _GEN_1655 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1592; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1965:29]
  wire [31:0] _GEN_1656 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1593; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1966:28]
  wire [31:0] _GEN_1657 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1594; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1967:29]
  wire [31:0] _GEN_1658 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1595; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1968:29]
  wire [31:0] _GEN_1659 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1596; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1969:29]
  wire [31:0] _GEN_1660 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1597; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1970:28]
  wire [31:0] _GEN_1661 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1598; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1971:29]
  wire [31:0] _GEN_1662 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1599; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1972:28]
  wire [31:0] _GEN_1663 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1600; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1973:29]
  wire [31:0] _GEN_1664 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1601; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1974:28]
  wire [31:0] _GEN_1665 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1602; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1975:29]
  wire [31:0] _GEN_1666 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1603; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1976:28]
  wire [31:0] _GEN_1667 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1604; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1977:29]
  wire [31:0] _GEN_1668 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1605; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1978:28]
  wire [31:0] _GEN_1669 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1606; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1979:29]
  wire [31:0] _GEN_1670 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1607; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1980:28]
  wire [31:0] _GEN_1671 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1608; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1981:29]
  wire [31:0] _GEN_1672 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1609; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1982:28]
  wire [31:0] _GEN_1673 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1610; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1983:29]
  wire [31:0] _GEN_1674 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1611; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1984:28]
  wire [31:0] _GEN_1675 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1612; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1985:29]
  wire [31:0] _GEN_1676 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1613; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1986:28]
  wire [31:0] _GEN_1677 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1614; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1987:29]
  wire [31:0] _GEN_1678 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1615; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1988:29]
  wire [31:0] _GEN_1679 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1616; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1989:29]
  wire [31:0] _GEN_1680 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1617; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1990:28]
  wire [31:0] _GEN_1681 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1618; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1991:29]
  wire [31:0] _GEN_1682 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1619; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1992:28]
  wire [31:0] _GEN_1683 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1620; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1993:29]
  wire [31:0] _GEN_1684 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1621; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1994:28]
  wire [31:0] _GEN_1685 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1622; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1995:29]
  wire [31:0] _GEN_1686 = _T_105 & LUT_stack_io_pop_4 ? 32'h0 : _GEN_1623; // @[stackmanage_35.scala 1926:68 stackmanage_35.scala 1996:28]
  wire [31:0] _GEN_1687 = _T_105 & LUT_stack_io_pop_3 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1856:28]
  wire [31:0] _GEN_1688 = _T_105 & LUT_stack_io_pop_3 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1857:27]
  wire [31:0] _GEN_1690 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1624; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1864:28]
  wire [31:0] _GEN_1691 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1625; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1865:27]
  wire [31:0] _GEN_1692 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1627; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1866:28]
  wire [31:0] _GEN_1693 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1628; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1867:27]
  wire [31:0] _GEN_1694 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1629; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1868:28]
  wire [31:0] _GEN_1695 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1630; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1869:27]
  wire [31:0] _GEN_1696 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1631; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1870:28]
  wire [31:0] _GEN_1697 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1632; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1871:27]
  wire [31:0] _GEN_1698 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1633; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1872:28]
  wire [31:0] _GEN_1699 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1634; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1873:27]
  wire [31:0] _GEN_1700 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1635; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1874:28]
  wire [31:0] _GEN_1701 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1636; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1875:27]
  wire [31:0] _GEN_1702 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1637; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1876:29]
  wire [31:0] _GEN_1703 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1638; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1877:29]
  wire [31:0] _GEN_1704 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1639; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1878:29]
  wire [31:0] _GEN_1705 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1640; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1879:28]
  wire [31:0] _GEN_1706 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1641; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1880:29]
  wire [31:0] _GEN_1707 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1642; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1881:28]
  wire [31:0] _GEN_1708 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1643; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1882:29]
  wire [31:0] _GEN_1709 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1644; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1883:28]
  wire [31:0] _GEN_1710 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1645; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1884:29]
  wire [31:0] _GEN_1711 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1646; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1885:28]
  wire [31:0] _GEN_1712 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1647; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1886:29]
  wire [31:0] _GEN_1713 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1648; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1887:28]
  wire [31:0] _GEN_1714 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1649; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1888:29]
  wire [31:0] _GEN_1715 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1650; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1889:28]
  wire [31:0] _GEN_1716 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1651; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1890:29]
  wire [31:0] _GEN_1717 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1652; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1891:28]
  wire [31:0] _GEN_1718 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1653; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1892:29]
  wire [31:0] _GEN_1719 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1654; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1893:28]
  wire [31:0] _GEN_1720 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1655; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1894:29]
  wire [31:0] _GEN_1721 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1656; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1895:28]
  wire [31:0] _GEN_1722 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1657; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1896:29]
  wire [31:0] _GEN_1723 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1658; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1897:29]
  wire [31:0] _GEN_1724 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1659; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1898:29]
  wire [31:0] _GEN_1725 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1660; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1899:28]
  wire [31:0] _GEN_1726 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1661; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1900:29]
  wire [31:0] _GEN_1727 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1662; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1901:28]
  wire [31:0] _GEN_1728 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1663; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1902:29]
  wire [31:0] _GEN_1729 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1664; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1903:28]
  wire [31:0] _GEN_1730 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1665; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1904:29]
  wire [31:0] _GEN_1731 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1666; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1905:28]
  wire [31:0] _GEN_1732 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1667; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1906:29]
  wire [31:0] _GEN_1733 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1668; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1907:28]
  wire [31:0] _GEN_1734 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1669; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1908:29]
  wire [31:0] _GEN_1735 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1670; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1909:28]
  wire [31:0] _GEN_1736 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1671; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1910:29]
  wire [31:0] _GEN_1737 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1672; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1911:28]
  wire [31:0] _GEN_1738 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1673; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1912:29]
  wire [31:0] _GEN_1739 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1674; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1913:28]
  wire [31:0] _GEN_1740 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1675; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1914:29]
  wire [31:0] _GEN_1741 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1676; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1915:28]
  wire [31:0] _GEN_1742 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1677; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1916:29]
  wire [31:0] _GEN_1743 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1678; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1917:29]
  wire [31:0] _GEN_1744 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1679; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1918:29]
  wire [31:0] _GEN_1745 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1680; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1919:28]
  wire [31:0] _GEN_1746 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1681; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1920:29]
  wire [31:0] _GEN_1747 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1682; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1921:28]
  wire [31:0] _GEN_1748 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1683; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1922:29]
  wire [31:0] _GEN_1749 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1684; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1923:28]
  wire [31:0] _GEN_1750 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1685; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1924:29]
  wire [31:0] _GEN_1751 = _T_105 & LUT_stack_io_pop_3 ? 32'h0 : _GEN_1686; // @[stackmanage_35.scala 1855:68 stackmanage_35.scala 1925:28]
  wire [31:0] _GEN_1752 = _T_105 & LUT_stack_io_pop_2 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1785:28]
  wire [31:0] _GEN_1753 = _T_105 & LUT_stack_io_pop_2 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1786:27]
  wire [31:0] _GEN_1755 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1687; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1791:28]
  wire [31:0] _GEN_1756 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1688; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1792:27]
  wire [31:0] _GEN_1757 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1690; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1793:28]
  wire [31:0] _GEN_1758 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1691; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1794:27]
  wire [31:0] _GEN_1759 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1692; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1795:28]
  wire [31:0] _GEN_1760 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1693; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1796:27]
  wire [31:0] _GEN_1761 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1694; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1797:28]
  wire [31:0] _GEN_1762 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1695; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1798:27]
  wire [31:0] _GEN_1763 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1696; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1799:28]
  wire [31:0] _GEN_1764 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1697; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1800:27]
  wire [31:0] _GEN_1765 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1698; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1801:28]
  wire [31:0] _GEN_1766 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1699; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1802:27]
  wire [31:0] _GEN_1767 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1700; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1803:28]
  wire [31:0] _GEN_1768 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1701; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1804:27]
  wire [31:0] _GEN_1769 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1702; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1805:29]
  wire [31:0] _GEN_1770 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1703; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1806:29]
  wire [31:0] _GEN_1771 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1704; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1807:29]
  wire [31:0] _GEN_1772 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1705; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1808:28]
  wire [31:0] _GEN_1773 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1706; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1809:29]
  wire [31:0] _GEN_1774 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1707; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1810:28]
  wire [31:0] _GEN_1775 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1708; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1811:29]
  wire [31:0] _GEN_1776 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1709; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1812:28]
  wire [31:0] _GEN_1777 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1710; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1813:29]
  wire [31:0] _GEN_1778 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1711; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1814:28]
  wire [31:0] _GEN_1779 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1712; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1815:29]
  wire [31:0] _GEN_1780 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1713; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1816:28]
  wire [31:0] _GEN_1781 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1714; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1817:29]
  wire [31:0] _GEN_1782 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1715; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1818:28]
  wire [31:0] _GEN_1783 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1716; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1819:29]
  wire [31:0] _GEN_1784 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1717; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1820:28]
  wire [31:0] _GEN_1785 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1718; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1821:29]
  wire [31:0] _GEN_1786 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1719; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1822:28]
  wire [31:0] _GEN_1787 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1720; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1823:29]
  wire [31:0] _GEN_1788 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1721; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1824:28]
  wire [31:0] _GEN_1789 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1722; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1825:29]
  wire [31:0] _GEN_1790 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1723; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1826:29]
  wire [31:0] _GEN_1791 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1724; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1827:29]
  wire [31:0] _GEN_1792 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1725; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1828:28]
  wire [31:0] _GEN_1793 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1726; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1829:29]
  wire [31:0] _GEN_1794 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1727; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1830:28]
  wire [31:0] _GEN_1795 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1728; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1831:29]
  wire [31:0] _GEN_1796 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1729; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1832:28]
  wire [31:0] _GEN_1797 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1730; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1833:29]
  wire [31:0] _GEN_1798 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1731; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1834:28]
  wire [31:0] _GEN_1799 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1732; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1835:29]
  wire [31:0] _GEN_1800 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1733; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1836:28]
  wire [31:0] _GEN_1801 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1734; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1837:29]
  wire [31:0] _GEN_1802 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1735; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1838:28]
  wire [31:0] _GEN_1803 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1736; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1839:29]
  wire [31:0] _GEN_1804 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1737; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1840:28]
  wire [31:0] _GEN_1805 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1738; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1841:29]
  wire [31:0] _GEN_1806 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1739; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1842:28]
  wire [31:0] _GEN_1807 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1740; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1843:29]
  wire [31:0] _GEN_1808 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1741; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1844:28]
  wire [31:0] _GEN_1809 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1742; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1845:29]
  wire [31:0] _GEN_1810 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1743; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1846:29]
  wire [31:0] _GEN_1811 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1744; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1847:29]
  wire [31:0] _GEN_1812 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1745; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1848:28]
  wire [31:0] _GEN_1813 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1746; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1849:29]
  wire [31:0] _GEN_1814 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1747; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1850:28]
  wire [31:0] _GEN_1815 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1748; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1851:29]
  wire [31:0] _GEN_1816 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1749; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1852:28]
  wire [31:0] _GEN_1817 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1750; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1853:29]
  wire [31:0] _GEN_1818 = _T_105 & LUT_stack_io_pop_2 ? 32'h0 : _GEN_1751; // @[stackmanage_35.scala 1784:68 stackmanage_35.scala 1854:28]
  wire [31:0] _GEN_1819 = _T_105 & LUT_stack_io_pop_1 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1714:28]
  wire [31:0] _GEN_1820 = _T_105 & LUT_stack_io_pop_1 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1715:27]
  wire [31:0] _GEN_1822 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1752; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1718:28]
  wire [31:0] _GEN_1823 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1753; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1719:27]
  wire [31:0] _GEN_1824 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1755; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1720:28]
  wire [31:0] _GEN_1825 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1756; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1721:27]
  wire [31:0] _GEN_1826 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1757; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1722:28]
  wire [31:0] _GEN_1827 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1758; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1723:27]
  wire [31:0] _GEN_1828 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1759; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1724:28]
  wire [31:0] _GEN_1829 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1760; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1725:27]
  wire [31:0] _GEN_1830 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1761; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1726:28]
  wire [31:0] _GEN_1831 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1762; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1727:27]
  wire [31:0] _GEN_1832 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1763; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1728:28]
  wire [31:0] _GEN_1833 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1764; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1729:27]
  wire [31:0] _GEN_1834 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1765; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1730:28]
  wire [31:0] _GEN_1835 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1766; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1731:27]
  wire [31:0] _GEN_1836 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1767; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1732:28]
  wire [31:0] _GEN_1837 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1768; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1733:27]
  wire [31:0] _GEN_1838 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1769; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1734:29]
  wire [31:0] _GEN_1839 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1770; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1735:29]
  wire [31:0] _GEN_1840 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1771; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1736:29]
  wire [31:0] _GEN_1841 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1772; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1737:28]
  wire [31:0] _GEN_1842 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1773; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1738:29]
  wire [31:0] _GEN_1843 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1774; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1739:28]
  wire [31:0] _GEN_1844 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1775; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1740:29]
  wire [31:0] _GEN_1845 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1776; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1741:28]
  wire [31:0] _GEN_1846 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1777; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1742:29]
  wire [31:0] _GEN_1847 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1778; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1743:28]
  wire [31:0] _GEN_1848 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1779; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1744:29]
  wire [31:0] _GEN_1849 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1780; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1745:28]
  wire [31:0] _GEN_1850 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1781; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1746:29]
  wire [31:0] _GEN_1851 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1782; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1747:28]
  wire [31:0] _GEN_1852 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1783; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1748:29]
  wire [31:0] _GEN_1853 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1784; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1749:28]
  wire [31:0] _GEN_1854 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1785; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1750:29]
  wire [31:0] _GEN_1855 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1786; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1751:28]
  wire [31:0] _GEN_1856 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1787; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1752:29]
  wire [31:0] _GEN_1857 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1788; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1753:28]
  wire [31:0] _GEN_1858 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1789; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1754:29]
  wire [31:0] _GEN_1859 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1790; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1755:29]
  wire [31:0] _GEN_1860 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1791; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1756:29]
  wire [31:0] _GEN_1861 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1792; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1757:28]
  wire [31:0] _GEN_1862 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1793; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1758:29]
  wire [31:0] _GEN_1863 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1794; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1759:28]
  wire [31:0] _GEN_1864 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1795; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1760:29]
  wire [31:0] _GEN_1865 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1796; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1761:28]
  wire [31:0] _GEN_1866 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1797; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1762:29]
  wire [31:0] _GEN_1867 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1798; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1763:28]
  wire [31:0] _GEN_1868 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1799; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1764:29]
  wire [31:0] _GEN_1869 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1800; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1765:28]
  wire [31:0] _GEN_1870 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1801; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1766:29]
  wire [31:0] _GEN_1871 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1802; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1767:28]
  wire [31:0] _GEN_1872 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1803; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1768:29]
  wire [31:0] _GEN_1873 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1804; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1769:28]
  wire [31:0] _GEN_1874 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1805; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1770:29]
  wire [31:0] _GEN_1875 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1806; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1771:28]
  wire [31:0] _GEN_1876 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1807; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1772:29]
  wire [31:0] _GEN_1877 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1808; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1773:28]
  wire [31:0] _GEN_1878 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1809; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1774:29]
  wire [31:0] _GEN_1879 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1810; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1775:29]
  wire [31:0] _GEN_1880 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1811; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1776:29]
  wire [31:0] _GEN_1881 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1812; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1777:28]
  wire [31:0] _GEN_1882 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1813; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1778:29]
  wire [31:0] _GEN_1883 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1814; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1779:28]
  wire [31:0] _GEN_1884 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1815; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1780:29]
  wire [31:0] _GEN_1885 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1816; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1781:28]
  wire [31:0] _GEN_1886 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1817; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1782:29]
  wire [31:0] _GEN_1887 = _T_105 & LUT_stack_io_pop_1 ? 32'h0 : _GEN_1818; // @[stackmanage_35.scala 1713:68 stackmanage_35.scala 1783:28]
  reg  pop_0; // @[stackmanage_35.scala 4201:46]
  reg  pop_1; // @[stackmanage_35.scala 4202:46]
  reg  pop_2; // @[stackmanage_35.scala 4203:46]
  reg  pop_3; // @[stackmanage_35.scala 4204:46]
  reg  pop_4; // @[stackmanage_35.scala 4205:46]
  reg  pop_5; // @[stackmanage_35.scala 4206:46]
  reg  pop_6; // @[stackmanage_35.scala 4207:46]
  reg  pop_7; // @[stackmanage_35.scala 4208:46]
  reg  pop_8; // @[stackmanage_35.scala 4209:46]
  reg  pop_9; // @[stackmanage_35.scala 4210:46]
  reg  pop_10; // @[stackmanage_35.scala 4212:47]
  reg  pop_11; // @[stackmanage_35.scala 4213:47]
  reg  pop_12; // @[stackmanage_35.scala 4214:47]
  reg  pop_13; // @[stackmanage_35.scala 4215:47]
  reg  pop_14; // @[stackmanage_35.scala 4216:47]
  reg  pop_15; // @[stackmanage_35.scala 4217:47]
  reg  pop_16; // @[stackmanage_35.scala 4218:47]
  reg  pop_17; // @[stackmanage_35.scala 4219:47]
  reg  pop_18; // @[stackmanage_35.scala 4220:47]
  reg  pop_19; // @[stackmanage_35.scala 4221:47]
  reg  pop_20; // @[stackmanage_35.scala 4223:47]
  reg  pop_21; // @[stackmanage_35.scala 4224:47]
  reg  pop_22; // @[stackmanage_35.scala 4225:47]
  reg  pop_23; // @[stackmanage_35.scala 4226:47]
  reg  pop_24; // @[stackmanage_35.scala 4227:47]
  reg  pop_25; // @[stackmanage_35.scala 4228:47]
  reg  pop_26; // @[stackmanage_35.scala 4229:47]
  reg  pop_27; // @[stackmanage_35.scala 4230:47]
  reg  pop_28; // @[stackmanage_35.scala 4231:47]
  reg  pop_29; // @[stackmanage_35.scala 4232:47]
  reg  pop_30; // @[stackmanage_35.scala 4234:47]
  reg  pop_31; // @[stackmanage_35.scala 4235:47]
  reg  pop_32; // @[stackmanage_35.scala 4236:47]
  reg  pop_33; // @[stackmanage_35.scala 4237:47]
  reg  pop_34; // @[stackmanage_35.scala 4238:47]
  wire  _T_314 = pop_34 & Stack_34_io_enable; // @[stackmanage_35.scala 4459:28]
  wire [31:0] _GEN_1958 = pop_34 & Stack_34_io_enable ? Stack_34_io_hit_out : 32'h0; // @[stackmanage_35.scala 4459:55 stackmanage_35.scala 4460:27 stackmanage_35.scala 4466:27]
  wire [31:0] _GEN_1959 = pop_34 & Stack_34_io_enable ? Stack_34_io_ray_out : 32'h0; // @[stackmanage_35.scala 4459:55 stackmanage_35.scala 4461:28 stackmanage_35.scala 4467:28]
  wire [31:0] _GEN_1960 = pop_34 & Stack_34_io_enable ? $signed(Stack_34_io_dataOut) : $signed(32'sh0); // @[stackmanage_35.scala 4459:55 stackmanage_35.scala 4462:25 stackmanage_35.scala 4468:25]
  wire [31:0] _GEN_1962 = pop_33 & Stack_33_io_enable ? Stack_33_io_hit_out : _GEN_1958; // @[stackmanage_35.scala 4454:55 stackmanage_35.scala 4455:27]
  wire [31:0] _GEN_1963 = pop_33 & Stack_33_io_enable ? Stack_33_io_ray_out : _GEN_1959; // @[stackmanage_35.scala 4454:55 stackmanage_35.scala 4456:28]
  wire [31:0] _GEN_1964 = pop_33 & Stack_33_io_enable ? $signed(Stack_33_io_dataOut) : $signed(_GEN_1960); // @[stackmanage_35.scala 4454:55 stackmanage_35.scala 4457:25]
  wire  _GEN_1965 = pop_33 & Stack_33_io_enable | _T_314; // @[stackmanage_35.scala 4454:55 stackmanage_35.scala 4458:31]
  wire [31:0] _GEN_1966 = pop_32 & Stack_32_io_enable ? Stack_32_io_hit_out : _GEN_1962; // @[stackmanage_35.scala 4449:55 stackmanage_35.scala 4450:27]
  wire [31:0] _GEN_1967 = pop_32 & Stack_32_io_enable ? Stack_32_io_ray_out : _GEN_1963; // @[stackmanage_35.scala 4449:55 stackmanage_35.scala 4451:28]
  wire [31:0] _GEN_1968 = pop_32 & Stack_32_io_enable ? $signed(Stack_32_io_dataOut) : $signed(_GEN_1964); // @[stackmanage_35.scala 4449:55 stackmanage_35.scala 4452:25]
  wire  _GEN_1969 = pop_32 & Stack_32_io_enable | _GEN_1965; // @[stackmanage_35.scala 4449:55 stackmanage_35.scala 4453:31]
  wire [31:0] _GEN_1970 = pop_31 & Stack_31_io_enable ? Stack_31_io_hit_out : _GEN_1966; // @[stackmanage_35.scala 4444:55 stackmanage_35.scala 4445:27]
  wire [31:0] _GEN_1971 = pop_31 & Stack_31_io_enable ? Stack_31_io_ray_out : _GEN_1967; // @[stackmanage_35.scala 4444:55 stackmanage_35.scala 4446:28]
  wire [31:0] _GEN_1972 = pop_31 & Stack_31_io_enable ? $signed(Stack_31_io_dataOut) : $signed(_GEN_1968); // @[stackmanage_35.scala 4444:55 stackmanage_35.scala 4447:25]
  wire  _GEN_1973 = pop_31 & Stack_31_io_enable | _GEN_1969; // @[stackmanage_35.scala 4444:55 stackmanage_35.scala 4448:31]
  wire [31:0] _GEN_1974 = pop_30 & Stack_30_io_enable ? Stack_30_io_hit_out : _GEN_1970; // @[stackmanage_35.scala 4439:55 stackmanage_35.scala 4440:27]
  wire [31:0] _GEN_1975 = pop_30 & Stack_30_io_enable ? Stack_30_io_ray_out : _GEN_1971; // @[stackmanage_35.scala 4439:55 stackmanage_35.scala 4441:28]
  wire [31:0] _GEN_1976 = pop_30 & Stack_30_io_enable ? $signed(Stack_30_io_dataOut) : $signed(_GEN_1972); // @[stackmanage_35.scala 4439:55 stackmanage_35.scala 4442:25]
  wire  _GEN_1977 = pop_30 & Stack_30_io_enable | _GEN_1973; // @[stackmanage_35.scala 4439:55 stackmanage_35.scala 4443:31]
  wire [31:0] _GEN_1978 = pop_29 & Stack_29_io_enable ? Stack_29_io_hit_out : _GEN_1974; // @[stackmanage_35.scala 4434:55 stackmanage_35.scala 4435:27]
  wire [31:0] _GEN_1979 = pop_29 & Stack_29_io_enable ? Stack_29_io_ray_out : _GEN_1975; // @[stackmanage_35.scala 4434:55 stackmanage_35.scala 4436:28]
  wire [31:0] _GEN_1980 = pop_29 & Stack_29_io_enable ? $signed(Stack_29_io_dataOut) : $signed(_GEN_1976); // @[stackmanage_35.scala 4434:55 stackmanage_35.scala 4437:25]
  wire  _GEN_1981 = pop_29 & Stack_29_io_enable | _GEN_1977; // @[stackmanage_35.scala 4434:55 stackmanage_35.scala 4438:31]
  wire [31:0] _GEN_1982 = pop_28 & Stack_28_io_enable ? Stack_28_io_hit_out : _GEN_1978; // @[stackmanage_35.scala 4429:55 stackmanage_35.scala 4430:27]
  wire [31:0] _GEN_1983 = pop_28 & Stack_28_io_enable ? Stack_28_io_ray_out : _GEN_1979; // @[stackmanage_35.scala 4429:55 stackmanage_35.scala 4431:28]
  wire [31:0] _GEN_1984 = pop_28 & Stack_28_io_enable ? $signed(Stack_28_io_dataOut) : $signed(_GEN_1980); // @[stackmanage_35.scala 4429:55 stackmanage_35.scala 4432:25]
  wire  _GEN_1985 = pop_28 & Stack_28_io_enable | _GEN_1981; // @[stackmanage_35.scala 4429:55 stackmanage_35.scala 4433:31]
  wire [31:0] _GEN_1986 = pop_27 & Stack_27_io_enable ? Stack_27_io_hit_out : _GEN_1982; // @[stackmanage_35.scala 4424:55 stackmanage_35.scala 4425:27]
  wire [31:0] _GEN_1987 = pop_27 & Stack_27_io_enable ? Stack_27_io_ray_out : _GEN_1983; // @[stackmanage_35.scala 4424:55 stackmanage_35.scala 4426:28]
  wire [31:0] _GEN_1988 = pop_27 & Stack_27_io_enable ? $signed(Stack_27_io_dataOut) : $signed(_GEN_1984); // @[stackmanage_35.scala 4424:55 stackmanage_35.scala 4427:25]
  wire  _GEN_1989 = pop_27 & Stack_27_io_enable | _GEN_1985; // @[stackmanage_35.scala 4424:55 stackmanage_35.scala 4428:31]
  wire [31:0] _GEN_1990 = pop_26 & Stack_26_io_enable ? Stack_26_io_hit_out : _GEN_1986; // @[stackmanage_35.scala 4419:55 stackmanage_35.scala 4420:27]
  wire [31:0] _GEN_1991 = pop_26 & Stack_26_io_enable ? Stack_26_io_ray_out : _GEN_1987; // @[stackmanage_35.scala 4419:55 stackmanage_35.scala 4421:28]
  wire [31:0] _GEN_1992 = pop_26 & Stack_26_io_enable ? $signed(Stack_26_io_dataOut) : $signed(_GEN_1988); // @[stackmanage_35.scala 4419:55 stackmanage_35.scala 4422:25]
  wire  _GEN_1993 = pop_26 & Stack_26_io_enable | _GEN_1989; // @[stackmanage_35.scala 4419:55 stackmanage_35.scala 4423:31]
  wire [31:0] _GEN_1994 = pop_25 & Stack_25_io_enable ? Stack_25_io_hit_out : _GEN_1990; // @[stackmanage_35.scala 4414:56 stackmanage_35.scala 4415:27]
  wire [31:0] _GEN_1995 = pop_25 & Stack_25_io_enable ? Stack_25_io_ray_out : _GEN_1991; // @[stackmanage_35.scala 4414:56 stackmanage_35.scala 4416:28]
  wire [31:0] _GEN_1996 = pop_25 & Stack_25_io_enable ? $signed(Stack_25_io_dataOut) : $signed(_GEN_1992); // @[stackmanage_35.scala 4414:56 stackmanage_35.scala 4417:25]
  wire  _GEN_1997 = pop_25 & Stack_25_io_enable | _GEN_1993; // @[stackmanage_35.scala 4414:56 stackmanage_35.scala 4418:31]
  wire [31:0] _GEN_1998 = pop_24 & Stack_24_io_enable ? Stack_24_io_hit_out : _GEN_1994; // @[stackmanage_35.scala 4409:55 stackmanage_35.scala 4410:27]
  wire [31:0] _GEN_1999 = pop_24 & Stack_24_io_enable ? Stack_24_io_ray_out : _GEN_1995; // @[stackmanage_35.scala 4409:55 stackmanage_35.scala 4411:28]
  wire [31:0] _GEN_2000 = pop_24 & Stack_24_io_enable ? $signed(Stack_24_io_dataOut) : $signed(_GEN_1996); // @[stackmanage_35.scala 4409:55 stackmanage_35.scala 4412:25]
  wire  _GEN_2001 = pop_24 & Stack_24_io_enable | _GEN_1997; // @[stackmanage_35.scala 4409:55 stackmanage_35.scala 4413:31]
  wire [31:0] _GEN_2002 = pop_23 & Stack_23_io_enable ? Stack_23_io_hit_out : _GEN_1998; // @[stackmanage_35.scala 4404:55 stackmanage_35.scala 4405:27]
  wire [31:0] _GEN_2003 = pop_23 & Stack_23_io_enable ? Stack_23_io_ray_out : _GEN_1999; // @[stackmanage_35.scala 4404:55 stackmanage_35.scala 4406:28]
  wire [31:0] _GEN_2004 = pop_23 & Stack_23_io_enable ? $signed(Stack_23_io_dataOut) : $signed(_GEN_2000); // @[stackmanage_35.scala 4404:55 stackmanage_35.scala 4407:25]
  wire  _GEN_2005 = pop_23 & Stack_23_io_enable | _GEN_2001; // @[stackmanage_35.scala 4404:55 stackmanage_35.scala 4408:31]
  wire [31:0] _GEN_2006 = pop_22 & Stack_22_io_enable ? Stack_22_io_hit_out : _GEN_2002; // @[stackmanage_35.scala 4399:55 stackmanage_35.scala 4400:27]
  wire [31:0] _GEN_2007 = pop_22 & Stack_22_io_enable ? Stack_22_io_ray_out : _GEN_2003; // @[stackmanage_35.scala 4399:55 stackmanage_35.scala 4401:28]
  wire [31:0] _GEN_2008 = pop_22 & Stack_22_io_enable ? $signed(Stack_22_io_dataOut) : $signed(_GEN_2004); // @[stackmanage_35.scala 4399:55 stackmanage_35.scala 4402:25]
  wire  _GEN_2009 = pop_22 & Stack_22_io_enable | _GEN_2005; // @[stackmanage_35.scala 4399:55 stackmanage_35.scala 4403:31]
  wire [31:0] _GEN_2010 = pop_21 & Stack_21_io_enable ? Stack_21_io_hit_out : _GEN_2006; // @[stackmanage_35.scala 4394:55 stackmanage_35.scala 4395:27]
  wire [31:0] _GEN_2011 = pop_21 & Stack_21_io_enable ? Stack_21_io_ray_out : _GEN_2007; // @[stackmanage_35.scala 4394:55 stackmanage_35.scala 4396:28]
  wire [31:0] _GEN_2012 = pop_21 & Stack_21_io_enable ? $signed(Stack_21_io_dataOut) : $signed(_GEN_2008); // @[stackmanage_35.scala 4394:55 stackmanage_35.scala 4397:25]
  wire  _GEN_2013 = pop_21 & Stack_21_io_enable | _GEN_2009; // @[stackmanage_35.scala 4394:55 stackmanage_35.scala 4398:31]
  wire [31:0] _GEN_2014 = pop_20 & Stack_20_io_enable ? Stack_20_io_hit_out : _GEN_2010; // @[stackmanage_35.scala 4389:55 stackmanage_35.scala 4390:27]
  wire [31:0] _GEN_2015 = pop_20 & Stack_20_io_enable ? Stack_20_io_ray_out : _GEN_2011; // @[stackmanage_35.scala 4389:55 stackmanage_35.scala 4391:28]
  wire [31:0] _GEN_2016 = pop_20 & Stack_20_io_enable ? $signed(Stack_20_io_dataOut) : $signed(_GEN_2012); // @[stackmanage_35.scala 4389:55 stackmanage_35.scala 4392:25]
  wire  _GEN_2017 = pop_20 & Stack_20_io_enable | _GEN_2013; // @[stackmanage_35.scala 4389:55 stackmanage_35.scala 4393:31]
  wire [31:0] _GEN_2018 = pop_19 & Stack_19_io_enable ? Stack_19_io_hit_out : _GEN_2014; // @[stackmanage_35.scala 4384:55 stackmanage_35.scala 4385:27]
  wire [31:0] _GEN_2019 = pop_19 & Stack_19_io_enable ? Stack_19_io_ray_out : _GEN_2015; // @[stackmanage_35.scala 4384:55 stackmanage_35.scala 4386:28]
  wire [31:0] _GEN_2020 = pop_19 & Stack_19_io_enable ? $signed(Stack_19_io_dataOut) : $signed(_GEN_2016); // @[stackmanage_35.scala 4384:55 stackmanage_35.scala 4387:25]
  wire  _GEN_2021 = pop_19 & Stack_19_io_enable | _GEN_2017; // @[stackmanage_35.scala 4384:55 stackmanage_35.scala 4388:31]
  wire [31:0] _GEN_2022 = pop_18 & Stack_18_io_enable ? Stack_18_io_hit_out : _GEN_2018; // @[stackmanage_35.scala 4379:55 stackmanage_35.scala 4380:27]
  wire [31:0] _GEN_2023 = pop_18 & Stack_18_io_enable ? Stack_18_io_ray_out : _GEN_2019; // @[stackmanage_35.scala 4379:55 stackmanage_35.scala 4381:28]
  wire [31:0] _GEN_2024 = pop_18 & Stack_18_io_enable ? $signed(Stack_18_io_dataOut) : $signed(_GEN_2020); // @[stackmanage_35.scala 4379:55 stackmanage_35.scala 4382:25]
  wire  _GEN_2025 = pop_18 & Stack_18_io_enable | _GEN_2021; // @[stackmanage_35.scala 4379:55 stackmanage_35.scala 4383:31]
  wire [31:0] _GEN_2026 = pop_17 & Stack_17_io_enable ? Stack_17_io_hit_out : _GEN_2022; // @[stackmanage_35.scala 4374:55 stackmanage_35.scala 4375:27]
  wire [31:0] _GEN_2027 = pop_17 & Stack_17_io_enable ? Stack_17_io_ray_out : _GEN_2023; // @[stackmanage_35.scala 4374:55 stackmanage_35.scala 4376:28]
  wire [31:0] _GEN_2028 = pop_17 & Stack_17_io_enable ? $signed(Stack_17_io_dataOut) : $signed(_GEN_2024); // @[stackmanage_35.scala 4374:55 stackmanage_35.scala 4377:25]
  wire  _GEN_2029 = pop_17 & Stack_17_io_enable | _GEN_2025; // @[stackmanage_35.scala 4374:55 stackmanage_35.scala 4378:31]
  wire [31:0] _GEN_2030 = pop_16 & Stack_16_io_enable ? Stack_16_io_hit_out : _GEN_2026; // @[stackmanage_35.scala 4369:55 stackmanage_35.scala 4370:27]
  wire [31:0] _GEN_2031 = pop_16 & Stack_16_io_enable ? Stack_16_io_ray_out : _GEN_2027; // @[stackmanage_35.scala 4369:55 stackmanage_35.scala 4371:28]
  wire [31:0] _GEN_2032 = pop_16 & Stack_16_io_enable ? $signed(Stack_16_io_dataOut) : $signed(_GEN_2028); // @[stackmanage_35.scala 4369:55 stackmanage_35.scala 4372:25]
  wire  _GEN_2033 = pop_16 & Stack_16_io_enable | _GEN_2029; // @[stackmanage_35.scala 4369:55 stackmanage_35.scala 4373:31]
  wire [31:0] _GEN_2034 = pop_15 & Stack_15_io_enable ? Stack_15_io_hit_out : _GEN_2030; // @[stackmanage_35.scala 4364:55 stackmanage_35.scala 4365:27]
  wire [31:0] _GEN_2035 = pop_15 & Stack_15_io_enable ? Stack_15_io_ray_out : _GEN_2031; // @[stackmanage_35.scala 4364:55 stackmanage_35.scala 4366:28]
  wire [31:0] _GEN_2036 = pop_15 & Stack_15_io_enable ? $signed(Stack_15_io_dataOut) : $signed(_GEN_2032); // @[stackmanage_35.scala 4364:55 stackmanage_35.scala 4367:25]
  wire  _GEN_2037 = pop_15 & Stack_15_io_enable | _GEN_2033; // @[stackmanage_35.scala 4364:55 stackmanage_35.scala 4368:31]
  wire [31:0] _GEN_2038 = pop_14 & Stack_14_io_enable ? Stack_14_io_hit_out : _GEN_2034; // @[stackmanage_35.scala 4359:55 stackmanage_35.scala 4360:27]
  wire [31:0] _GEN_2039 = pop_14 & Stack_14_io_enable ? Stack_14_io_ray_out : _GEN_2035; // @[stackmanage_35.scala 4359:55 stackmanage_35.scala 4361:28]
  wire [31:0] _GEN_2040 = pop_14 & Stack_14_io_enable ? $signed(Stack_14_io_dataOut) : $signed(_GEN_2036); // @[stackmanage_35.scala 4359:55 stackmanage_35.scala 4362:25]
  wire  _GEN_2041 = pop_14 & Stack_14_io_enable | _GEN_2037; // @[stackmanage_35.scala 4359:55 stackmanage_35.scala 4363:31]
  wire [31:0] _GEN_2042 = pop_13 & Stack_13_io_enable ? Stack_13_io_hit_out : _GEN_2038; // @[stackmanage_35.scala 4354:55 stackmanage_35.scala 4355:27]
  wire [31:0] _GEN_2043 = pop_13 & Stack_13_io_enable ? Stack_13_io_ray_out : _GEN_2039; // @[stackmanage_35.scala 4354:55 stackmanage_35.scala 4356:28]
  wire [31:0] _GEN_2044 = pop_13 & Stack_13_io_enable ? $signed(Stack_13_io_dataOut) : $signed(_GEN_2040); // @[stackmanage_35.scala 4354:55 stackmanage_35.scala 4357:25]
  wire  _GEN_2045 = pop_13 & Stack_13_io_enable | _GEN_2041; // @[stackmanage_35.scala 4354:55 stackmanage_35.scala 4358:31]
  wire [31:0] _GEN_2046 = pop_12 & Stack_12_io_enable ? Stack_12_io_hit_out : _GEN_2042; // @[stackmanage_35.scala 4349:55 stackmanage_35.scala 4350:27]
  wire [31:0] _GEN_2047 = pop_12 & Stack_12_io_enable ? Stack_12_io_ray_out : _GEN_2043; // @[stackmanage_35.scala 4349:55 stackmanage_35.scala 4351:28]
  wire [31:0] _GEN_2048 = pop_12 & Stack_12_io_enable ? $signed(Stack_12_io_dataOut) : $signed(_GEN_2044); // @[stackmanage_35.scala 4349:55 stackmanage_35.scala 4352:25]
  wire  _GEN_2049 = pop_12 & Stack_12_io_enable | _GEN_2045; // @[stackmanage_35.scala 4349:55 stackmanage_35.scala 4353:31]
  wire [31:0] _GEN_2050 = pop_11 & Stack_11_io_enable ? Stack_11_io_hit_out : _GEN_2046; // @[stackmanage_35.scala 4344:55 stackmanage_35.scala 4345:27]
  wire [31:0] _GEN_2051 = pop_11 & Stack_11_io_enable ? Stack_11_io_ray_out : _GEN_2047; // @[stackmanage_35.scala 4344:55 stackmanage_35.scala 4346:28]
  wire [31:0] _GEN_2052 = pop_11 & Stack_11_io_enable ? $signed(Stack_11_io_dataOut) : $signed(_GEN_2048); // @[stackmanage_35.scala 4344:55 stackmanage_35.scala 4347:25]
  wire  _GEN_2053 = pop_11 & Stack_11_io_enable | _GEN_2049; // @[stackmanage_35.scala 4344:55 stackmanage_35.scala 4348:31]
  wire [31:0] _GEN_2054 = pop_10 & Stack_10_io_enable ? Stack_10_io_hit_out : _GEN_2050; // @[stackmanage_35.scala 4339:55 stackmanage_35.scala 4340:27]
  wire [31:0] _GEN_2055 = pop_10 & Stack_10_io_enable ? Stack_10_io_ray_out : _GEN_2051; // @[stackmanage_35.scala 4339:55 stackmanage_35.scala 4341:28]
  wire [31:0] _GEN_2056 = pop_10 & Stack_10_io_enable ? $signed(Stack_10_io_dataOut) : $signed(_GEN_2052); // @[stackmanage_35.scala 4339:55 stackmanage_35.scala 4342:25]
  wire  _GEN_2057 = pop_10 & Stack_10_io_enable | _GEN_2053; // @[stackmanage_35.scala 4339:55 stackmanage_35.scala 4343:31]
  wire [31:0] _GEN_2058 = pop_9 & Stack_9_io_enable ? Stack_9_io_hit_out : _GEN_2054; // @[stackmanage_35.scala 4334:53 stackmanage_35.scala 4335:27]
  wire [31:0] _GEN_2059 = pop_9 & Stack_9_io_enable ? Stack_9_io_ray_out : _GEN_2055; // @[stackmanage_35.scala 4334:53 stackmanage_35.scala 4336:28]
  wire [31:0] _GEN_2060 = pop_9 & Stack_9_io_enable ? $signed(Stack_9_io_dataOut) : $signed(_GEN_2056); // @[stackmanage_35.scala 4334:53 stackmanage_35.scala 4337:25]
  wire  _GEN_2061 = pop_9 & Stack_9_io_enable | _GEN_2057; // @[stackmanage_35.scala 4334:53 stackmanage_35.scala 4338:31]
  wire [31:0] _GEN_2062 = pop_8 & Stack_8_io_enable ? Stack_8_io_hit_out : _GEN_2058; // @[stackmanage_35.scala 4329:53 stackmanage_35.scala 4330:27]
  wire [31:0] _GEN_2063 = pop_8 & Stack_8_io_enable ? Stack_8_io_ray_out : _GEN_2059; // @[stackmanage_35.scala 4329:53 stackmanage_35.scala 4331:28]
  wire [31:0] _GEN_2064 = pop_8 & Stack_8_io_enable ? $signed(Stack_8_io_dataOut) : $signed(_GEN_2060); // @[stackmanage_35.scala 4329:53 stackmanage_35.scala 4332:25]
  wire  _GEN_2065 = pop_8 & Stack_8_io_enable | _GEN_2061; // @[stackmanage_35.scala 4329:53 stackmanage_35.scala 4333:31]
  wire [31:0] _GEN_2066 = pop_7 & Stack_7_io_enable ? Stack_7_io_hit_out : _GEN_2062; // @[stackmanage_35.scala 4324:53 stackmanage_35.scala 4325:27]
  wire [31:0] _GEN_2067 = pop_7 & Stack_7_io_enable ? Stack_7_io_ray_out : _GEN_2063; // @[stackmanage_35.scala 4324:53 stackmanage_35.scala 4326:28]
  wire [31:0] _GEN_2068 = pop_7 & Stack_7_io_enable ? $signed(Stack_7_io_dataOut) : $signed(_GEN_2064); // @[stackmanage_35.scala 4324:53 stackmanage_35.scala 4327:25]
  wire  _GEN_2069 = pop_7 & Stack_7_io_enable | _GEN_2065; // @[stackmanage_35.scala 4324:53 stackmanage_35.scala 4328:31]
  wire [31:0] _GEN_2070 = pop_6 & Stack_6_io_enable ? Stack_6_io_hit_out : _GEN_2066; // @[stackmanage_35.scala 4319:53 stackmanage_35.scala 4320:27]
  wire [31:0] _GEN_2071 = pop_6 & Stack_6_io_enable ? Stack_6_io_ray_out : _GEN_2067; // @[stackmanage_35.scala 4319:53 stackmanage_35.scala 4321:28]
  wire [31:0] _GEN_2072 = pop_6 & Stack_6_io_enable ? $signed(Stack_6_io_dataOut) : $signed(_GEN_2068); // @[stackmanage_35.scala 4319:53 stackmanage_35.scala 4322:25]
  wire  _GEN_2073 = pop_6 & Stack_6_io_enable | _GEN_2069; // @[stackmanage_35.scala 4319:53 stackmanage_35.scala 4323:31]
  wire [31:0] _GEN_2074 = pop_5 & Stack_5_io_enable ? Stack_5_io_hit_out : _GEN_2070; // @[stackmanage_35.scala 4314:53 stackmanage_35.scala 4315:27]
  wire [31:0] _GEN_2075 = pop_5 & Stack_5_io_enable ? Stack_5_io_ray_out : _GEN_2071; // @[stackmanage_35.scala 4314:53 stackmanage_35.scala 4316:28]
  wire [31:0] _GEN_2076 = pop_5 & Stack_5_io_enable ? $signed(Stack_5_io_dataOut) : $signed(_GEN_2072); // @[stackmanage_35.scala 4314:53 stackmanage_35.scala 4317:25]
  wire  _GEN_2077 = pop_5 & Stack_5_io_enable | _GEN_2073; // @[stackmanage_35.scala 4314:53 stackmanage_35.scala 4318:31]
  wire [31:0] _GEN_2078 = pop_4 & Stack_4_io_enable ? Stack_4_io_hit_out : _GEN_2074; // @[stackmanage_35.scala 4309:53 stackmanage_35.scala 4310:27]
  wire [31:0] _GEN_2079 = pop_4 & Stack_4_io_enable ? Stack_4_io_ray_out : _GEN_2075; // @[stackmanage_35.scala 4309:53 stackmanage_35.scala 4311:28]
  wire [31:0] _GEN_2080 = pop_4 & Stack_4_io_enable ? $signed(Stack_4_io_dataOut) : $signed(_GEN_2076); // @[stackmanage_35.scala 4309:53 stackmanage_35.scala 4312:25]
  wire  _GEN_2081 = pop_4 & Stack_4_io_enable | _GEN_2077; // @[stackmanage_35.scala 4309:53 stackmanage_35.scala 4313:31]
  wire [31:0] _GEN_2082 = pop_3 & Stack_3_io_enable ? Stack_3_io_hit_out : _GEN_2078; // @[stackmanage_35.scala 4304:53 stackmanage_35.scala 4305:27]
  wire [31:0] _GEN_2083 = pop_3 & Stack_3_io_enable ? Stack_3_io_ray_out : _GEN_2079; // @[stackmanage_35.scala 4304:53 stackmanage_35.scala 4306:28]
  wire [31:0] _GEN_2084 = pop_3 & Stack_3_io_enable ? $signed(Stack_3_io_dataOut) : $signed(_GEN_2080); // @[stackmanage_35.scala 4304:53 stackmanage_35.scala 4307:25]
  wire  _GEN_2085 = pop_3 & Stack_3_io_enable | _GEN_2081; // @[stackmanage_35.scala 4304:53 stackmanage_35.scala 4308:31]
  wire  _GEN_2089 = pop_2 & Stack_2_io_enable | _GEN_2085; // @[stackmanage_35.scala 4299:53 stackmanage_35.scala 4303:31]
  wire  _GEN_2093 = pop_1 & Stack_1_io_enable | _GEN_2089; // @[stackmanage_35.scala 4294:53 stackmanage_35.scala 4298:31]
  wire  _GEN_2097 = pop_0 & Stack_0_io_enable | _GEN_2093; // @[stackmanage_35.scala 4288:48 stackmanage_35.scala 4293:31]
  reg  dispatch_0; // @[stackmanage_35.scala 4476:41]
  reg  dispatch_1; // @[stackmanage_35.scala 4477:41]
  reg  dispatch_2; // @[stackmanage_35.scala 4478:41]
  reg  dispatch_3; // @[stackmanage_35.scala 4479:41]
  reg  dispatch_4; // @[stackmanage_35.scala 4480:41]
  reg  dispatch_5; // @[stackmanage_35.scala 4481:41]
  reg  dispatch_6; // @[stackmanage_35.scala 4482:41]
  reg  dispatch_7; // @[stackmanage_35.scala 4483:41]
  reg  dispatch_8; // @[stackmanage_35.scala 4484:41]
  reg  dispatch_9; // @[stackmanage_35.scala 4485:41]
  reg  dispatch_10; // @[stackmanage_35.scala 4487:42]
  reg  dispatch_11; // @[stackmanage_35.scala 4488:42]
  reg  dispatch_12; // @[stackmanage_35.scala 4489:42]
  reg  dispatch_13; // @[stackmanage_35.scala 4490:42]
  reg  dispatch_14; // @[stackmanage_35.scala 4491:42]
  reg  dispatch_15; // @[stackmanage_35.scala 4492:42]
  reg  dispatch_16; // @[stackmanage_35.scala 4493:42]
  reg  dispatch_17; // @[stackmanage_35.scala 4494:42]
  reg  dispatch_18; // @[stackmanage_35.scala 4495:42]
  reg  dispatch_19; // @[stackmanage_35.scala 4496:42]
  reg  dispatch_20; // @[stackmanage_35.scala 4498:42]
  reg  dispatch_21; // @[stackmanage_35.scala 4499:42]
  reg  dispatch_22; // @[stackmanage_35.scala 4500:42]
  reg  dispatch_23; // @[stackmanage_35.scala 4501:42]
  reg  dispatch_24; // @[stackmanage_35.scala 4502:42]
  reg  dispatch_25; // @[stackmanage_35.scala 4503:42]
  reg  dispatch_26; // @[stackmanage_35.scala 4504:42]
  reg  dispatch_27; // @[stackmanage_35.scala 4505:42]
  reg  dispatch_28; // @[stackmanage_35.scala 4506:42]
  reg  dispatch_29; // @[stackmanage_35.scala 4507:42]
  reg  dispatch_30; // @[stackmanage_35.scala 4509:42]
  reg  dispatch_31; // @[stackmanage_35.scala 4510:42]
  reg  dispatch_32; // @[stackmanage_35.scala 4511:42]
  reg  dispatch_33; // @[stackmanage_35.scala 4512:42]
  reg  dispatch_34; // @[stackmanage_35.scala 4513:42]
  reg  dispatch_no_match; // @[stackmanage_35.scala 4514:42]
  reg  empty_0; // @[stackmanage_35.scala 4518:42]
  reg  empty_1; // @[stackmanage_35.scala 4519:42]
  reg  empty_2; // @[stackmanage_35.scala 4520:42]
  reg  empty_3; // @[stackmanage_35.scala 4521:42]
  reg  empty_4; // @[stackmanage_35.scala 4522:42]
  reg  empty_5; // @[stackmanage_35.scala 4523:42]
  reg  empty_6; // @[stackmanage_35.scala 4524:42]
  reg  empty_7; // @[stackmanage_35.scala 4525:42]
  reg  empty_8; // @[stackmanage_35.scala 4526:42]
  reg  empty_9; // @[stackmanage_35.scala 4527:42]
  reg  empty_10; // @[stackmanage_35.scala 4529:43]
  reg  empty_11; // @[stackmanage_35.scala 4530:43]
  reg  empty_12; // @[stackmanage_35.scala 4531:43]
  reg  empty_13; // @[stackmanage_35.scala 4532:43]
  reg  empty_14; // @[stackmanage_35.scala 4533:43]
  reg  empty_15; // @[stackmanage_35.scala 4534:43]
  reg  empty_16; // @[stackmanage_35.scala 4535:43]
  reg  empty_17; // @[stackmanage_35.scala 4536:43]
  reg  empty_18; // @[stackmanage_35.scala 4537:43]
  reg  empty_19; // @[stackmanage_35.scala 4538:43]
  reg  empty_20; // @[stackmanage_35.scala 4540:43]
  reg  empty_21; // @[stackmanage_35.scala 4541:43]
  reg  empty_22; // @[stackmanage_35.scala 4542:43]
  reg  empty_23; // @[stackmanage_35.scala 4543:43]
  reg  empty_24; // @[stackmanage_35.scala 4544:43]
  reg  empty_25; // @[stackmanage_35.scala 4545:43]
  reg  empty_26; // @[stackmanage_35.scala 4546:43]
  reg  empty_27; // @[stackmanage_35.scala 4547:43]
  reg  empty_28; // @[stackmanage_35.scala 4548:43]
  reg  empty_29; // @[stackmanage_35.scala 4549:43]
  reg  empty_30; // @[stackmanage_35.scala 4551:43]
  reg  empty_31; // @[stackmanage_35.scala 4552:43]
  reg  empty_32; // @[stackmanage_35.scala 4553:43]
  reg  empty_33; // @[stackmanage_35.scala 4554:43]
  reg  empty_34; // @[stackmanage_35.scala 4555:43]
  wire  _T_317 = pop_0 & empty_0; // @[stackmanage_35.scala 4599:22]
  wire  _T_320 = pop_1 & empty_1; // @[stackmanage_35.scala 4635:27]
  wire  _T_323 = pop_2 & empty_2; // @[stackmanage_35.scala 4672:27]
  wire  _T_326 = pop_3 & empty_3; // @[stackmanage_35.scala 4710:27]
  wire  _T_329 = pop_4 & empty_4; // @[stackmanage_35.scala 4748:27]
  wire  _T_332 = pop_5 & empty_5; // @[stackmanage_35.scala 4786:27]
  wire  _T_335 = pop_6 & empty_6; // @[stackmanage_35.scala 4824:27]
  wire  _T_338 = pop_7 & empty_7; // @[stackmanage_35.scala 4862:27]
  wire  _T_341 = pop_8 & empty_8; // @[stackmanage_35.scala 4900:27]
  wire  _T_344 = pop_9 & empty_9; // @[stackmanage_35.scala 4937:27]
  wire  _T_347 = pop_10 & empty_10; // @[stackmanage_35.scala 4975:28]
  wire  _T_350 = pop_11 & empty_11; // @[stackmanage_35.scala 5012:28]
  wire  _T_353 = pop_12 & empty_12; // @[stackmanage_35.scala 5049:28]
  wire  _T_356 = pop_13 & empty_13; // @[stackmanage_35.scala 5086:28]
  wire  _T_359 = pop_14 & empty_14; // @[stackmanage_35.scala 5123:28]
  wire  _T_362 = pop_15 & empty_15; // @[stackmanage_35.scala 5160:28]
  wire  _T_365 = pop_16 & empty_16; // @[stackmanage_35.scala 5197:28]
  wire  _T_368 = pop_17 & empty_17; // @[stackmanage_35.scala 5234:28]
  wire  _T_371 = pop_18 & empty_18; // @[stackmanage_35.scala 5271:28]
  wire  _T_374 = pop_19 & empty_19; // @[stackmanage_35.scala 5308:28]
  wire  _T_377 = pop_20 & empty_20; // @[stackmanage_35.scala 5345:28]
  wire  _T_380 = pop_21 & empty_21; // @[stackmanage_35.scala 5382:28]
  wire  _T_383 = pop_22 & empty_22; // @[stackmanage_35.scala 5419:28]
  wire  _T_386 = pop_23 & empty_23; // @[stackmanage_35.scala 5456:28]
  wire  _T_389 = pop_24 & empty_24; // @[stackmanage_35.scala 5493:28]
  wire  _T_392 = pop_25 & empty_25; // @[stackmanage_35.scala 5530:28]
  wire  _T_395 = pop_26 & empty_26; // @[stackmanage_35.scala 5567:30]
  wire  _T_398 = pop_27 & empty_27; // @[stackmanage_35.scala 5604:28]
  wire  _T_401 = pop_28 & empty_28; // @[stackmanage_35.scala 5641:28]
  wire  _T_404 = pop_29 & empty_29; // @[stackmanage_35.scala 5678:28]
  wire  _T_407 = pop_30 & empty_30; // @[stackmanage_35.scala 5715:29]
  wire  _T_410 = pop_31 & empty_31; // @[stackmanage_35.scala 5752:29]
  wire  _T_413 = pop_32 & empty_32; // @[stackmanage_35.scala 5789:29]
  wire  _T_416 = pop_33 & empty_33; // @[stackmanage_35.scala 5827:29]
  wire  _T_419 = pop_34 & empty_34; // @[stackmanage_35.scala 5864:29]
  wire  _GEN_2102 = pop_33 & empty_33 ? 1'h0 : _T_419; // @[stackmanage_35.scala 5827:46 stackmanage_35.scala 5863:34]
  wire  _GEN_2105 = pop_32 & empty_32 ? 1'h0 : _T_416; // @[stackmanage_35.scala 5789:46 stackmanage_35.scala 5824:34]
  wire  _GEN_2106 = pop_32 & empty_32 ? 1'h0 : _GEN_2102; // @[stackmanage_35.scala 5789:46 stackmanage_35.scala 5825:34]
  wire  _GEN_2109 = pop_31 & empty_31 ? 1'h0 : _T_413; // @[stackmanage_35.scala 5752:46 stackmanage_35.scala 5786:34]
  wire  _GEN_2110 = pop_31 & empty_31 ? 1'h0 : _GEN_2105; // @[stackmanage_35.scala 5752:46 stackmanage_35.scala 5787:34]
  wire  _GEN_2111 = pop_31 & empty_31 ? 1'h0 : _GEN_2106; // @[stackmanage_35.scala 5752:46 stackmanage_35.scala 5788:34]
  wire  _GEN_2114 = pop_30 & empty_30 ? 1'h0 : _T_410; // @[stackmanage_35.scala 5715:46 stackmanage_35.scala 5748:34]
  wire  _GEN_2115 = pop_30 & empty_30 ? 1'h0 : _GEN_2109; // @[stackmanage_35.scala 5715:46 stackmanage_35.scala 5749:34]
  wire  _GEN_2116 = pop_30 & empty_30 ? 1'h0 : _GEN_2110; // @[stackmanage_35.scala 5715:46 stackmanage_35.scala 5750:34]
  wire  _GEN_2117 = pop_30 & empty_30 ? 1'h0 : _GEN_2111; // @[stackmanage_35.scala 5715:46 stackmanage_35.scala 5751:34]
  wire  _GEN_2120 = pop_29 & empty_29 ? 1'h0 : _T_407; // @[stackmanage_35.scala 5678:45 stackmanage_35.scala 5710:34]
  wire  _GEN_2121 = pop_29 & empty_29 ? 1'h0 : _GEN_2114; // @[stackmanage_35.scala 5678:45 stackmanage_35.scala 5711:34]
  wire  _GEN_2122 = pop_29 & empty_29 ? 1'h0 : _GEN_2115; // @[stackmanage_35.scala 5678:45 stackmanage_35.scala 5712:34]
  wire  _GEN_2123 = pop_29 & empty_29 ? 1'h0 : _GEN_2116; // @[stackmanage_35.scala 5678:45 stackmanage_35.scala 5713:34]
  wire  _GEN_2124 = pop_29 & empty_29 ? 1'h0 : _GEN_2117; // @[stackmanage_35.scala 5678:45 stackmanage_35.scala 5714:34]
  wire  _GEN_2127 = pop_28 & empty_28 ? 1'h0 : _T_404; // @[stackmanage_35.scala 5641:45 stackmanage_35.scala 5672:34]
  wire  _GEN_2128 = pop_28 & empty_28 ? 1'h0 : _GEN_2120; // @[stackmanage_35.scala 5641:45 stackmanage_35.scala 5673:34]
  wire  _GEN_2129 = pop_28 & empty_28 ? 1'h0 : _GEN_2121; // @[stackmanage_35.scala 5641:45 stackmanage_35.scala 5674:34]
  wire  _GEN_2130 = pop_28 & empty_28 ? 1'h0 : _GEN_2122; // @[stackmanage_35.scala 5641:45 stackmanage_35.scala 5675:34]
  wire  _GEN_2131 = pop_28 & empty_28 ? 1'h0 : _GEN_2123; // @[stackmanage_35.scala 5641:45 stackmanage_35.scala 5676:34]
  wire  _GEN_2132 = pop_28 & empty_28 ? 1'h0 : _GEN_2124; // @[stackmanage_35.scala 5641:45 stackmanage_35.scala 5677:34]
  wire  _GEN_2135 = pop_27 & empty_27 ? 1'h0 : _T_401; // @[stackmanage_35.scala 5604:45 stackmanage_35.scala 5634:34]
  wire  _GEN_2136 = pop_27 & empty_27 ? 1'h0 : _GEN_2127; // @[stackmanage_35.scala 5604:45 stackmanage_35.scala 5635:34]
  wire  _GEN_2137 = pop_27 & empty_27 ? 1'h0 : _GEN_2128; // @[stackmanage_35.scala 5604:45 stackmanage_35.scala 5636:34]
  wire  _GEN_2138 = pop_27 & empty_27 ? 1'h0 : _GEN_2129; // @[stackmanage_35.scala 5604:45 stackmanage_35.scala 5637:34]
  wire  _GEN_2139 = pop_27 & empty_27 ? 1'h0 : _GEN_2130; // @[stackmanage_35.scala 5604:45 stackmanage_35.scala 5638:34]
  wire  _GEN_2140 = pop_27 & empty_27 ? 1'h0 : _GEN_2131; // @[stackmanage_35.scala 5604:45 stackmanage_35.scala 5639:34]
  wire  _GEN_2141 = pop_27 & empty_27 ? 1'h0 : _GEN_2132; // @[stackmanage_35.scala 5604:45 stackmanage_35.scala 5640:34]
  wire  _GEN_2144 = pop_26 & empty_26 ? 1'h0 : _T_398; // @[stackmanage_35.scala 5567:47 stackmanage_35.scala 5596:34]
  wire  _GEN_2145 = pop_26 & empty_26 ? 1'h0 : _GEN_2135; // @[stackmanage_35.scala 5567:47 stackmanage_35.scala 5597:34]
  wire  _GEN_2146 = pop_26 & empty_26 ? 1'h0 : _GEN_2136; // @[stackmanage_35.scala 5567:47 stackmanage_35.scala 5598:34]
  wire  _GEN_2147 = pop_26 & empty_26 ? 1'h0 : _GEN_2137; // @[stackmanage_35.scala 5567:47 stackmanage_35.scala 5599:34]
  wire  _GEN_2148 = pop_26 & empty_26 ? 1'h0 : _GEN_2138; // @[stackmanage_35.scala 5567:47 stackmanage_35.scala 5600:34]
  wire  _GEN_2149 = pop_26 & empty_26 ? 1'h0 : _GEN_2139; // @[stackmanage_35.scala 5567:47 stackmanage_35.scala 5601:34]
  wire  _GEN_2150 = pop_26 & empty_26 ? 1'h0 : _GEN_2140; // @[stackmanage_35.scala 5567:47 stackmanage_35.scala 5602:34]
  wire  _GEN_2151 = pop_26 & empty_26 ? 1'h0 : _GEN_2141; // @[stackmanage_35.scala 5567:47 stackmanage_35.scala 5603:34]
  wire  _GEN_2154 = pop_25 & empty_25 ? 1'h0 : _T_395; // @[stackmanage_35.scala 5530:45 stackmanage_35.scala 5558:34]
  wire  _GEN_2155 = pop_25 & empty_25 ? 1'h0 : _GEN_2144; // @[stackmanage_35.scala 5530:45 stackmanage_35.scala 5559:34]
  wire  _GEN_2156 = pop_25 & empty_25 ? 1'h0 : _GEN_2145; // @[stackmanage_35.scala 5530:45 stackmanage_35.scala 5560:34]
  wire  _GEN_2157 = pop_25 & empty_25 ? 1'h0 : _GEN_2146; // @[stackmanage_35.scala 5530:45 stackmanage_35.scala 5561:34]
  wire  _GEN_2158 = pop_25 & empty_25 ? 1'h0 : _GEN_2147; // @[stackmanage_35.scala 5530:45 stackmanage_35.scala 5562:34]
  wire  _GEN_2159 = pop_25 & empty_25 ? 1'h0 : _GEN_2148; // @[stackmanage_35.scala 5530:45 stackmanage_35.scala 5563:34]
  wire  _GEN_2160 = pop_25 & empty_25 ? 1'h0 : _GEN_2149; // @[stackmanage_35.scala 5530:45 stackmanage_35.scala 5564:34]
  wire  _GEN_2161 = pop_25 & empty_25 ? 1'h0 : _GEN_2150; // @[stackmanage_35.scala 5530:45 stackmanage_35.scala 5565:34]
  wire  _GEN_2162 = pop_25 & empty_25 ? 1'h0 : _GEN_2151; // @[stackmanage_35.scala 5530:45 stackmanage_35.scala 5566:34]
  wire  _GEN_2165 = pop_24 & empty_24 ? 1'h0 : _T_392; // @[stackmanage_35.scala 5493:45 stackmanage_35.scala 5520:34]
  wire  _GEN_2166 = pop_24 & empty_24 ? 1'h0 : _GEN_2154; // @[stackmanage_35.scala 5493:45 stackmanage_35.scala 5521:34]
  wire  _GEN_2167 = pop_24 & empty_24 ? 1'h0 : _GEN_2155; // @[stackmanage_35.scala 5493:45 stackmanage_35.scala 5522:34]
  wire  _GEN_2168 = pop_24 & empty_24 ? 1'h0 : _GEN_2156; // @[stackmanage_35.scala 5493:45 stackmanage_35.scala 5523:34]
  wire  _GEN_2169 = pop_24 & empty_24 ? 1'h0 : _GEN_2157; // @[stackmanage_35.scala 5493:45 stackmanage_35.scala 5524:34]
  wire  _GEN_2170 = pop_24 & empty_24 ? 1'h0 : _GEN_2158; // @[stackmanage_35.scala 5493:45 stackmanage_35.scala 5525:34]
  wire  _GEN_2171 = pop_24 & empty_24 ? 1'h0 : _GEN_2159; // @[stackmanage_35.scala 5493:45 stackmanage_35.scala 5526:34]
  wire  _GEN_2172 = pop_24 & empty_24 ? 1'h0 : _GEN_2160; // @[stackmanage_35.scala 5493:45 stackmanage_35.scala 5527:34]
  wire  _GEN_2173 = pop_24 & empty_24 ? 1'h0 : _GEN_2161; // @[stackmanage_35.scala 5493:45 stackmanage_35.scala 5528:34]
  wire  _GEN_2174 = pop_24 & empty_24 ? 1'h0 : _GEN_2162; // @[stackmanage_35.scala 5493:45 stackmanage_35.scala 5529:34]
  wire  _GEN_2177 = pop_23 & empty_23 ? 1'h0 : _T_389; // @[stackmanage_35.scala 5456:45 stackmanage_35.scala 5482:34]
  wire  _GEN_2178 = pop_23 & empty_23 ? 1'h0 : _GEN_2165; // @[stackmanage_35.scala 5456:45 stackmanage_35.scala 5483:34]
  wire  _GEN_2179 = pop_23 & empty_23 ? 1'h0 : _GEN_2166; // @[stackmanage_35.scala 5456:45 stackmanage_35.scala 5484:34]
  wire  _GEN_2180 = pop_23 & empty_23 ? 1'h0 : _GEN_2167; // @[stackmanage_35.scala 5456:45 stackmanage_35.scala 5485:34]
  wire  _GEN_2181 = pop_23 & empty_23 ? 1'h0 : _GEN_2168; // @[stackmanage_35.scala 5456:45 stackmanage_35.scala 5486:34]
  wire  _GEN_2182 = pop_23 & empty_23 ? 1'h0 : _GEN_2169; // @[stackmanage_35.scala 5456:45 stackmanage_35.scala 5487:34]
  wire  _GEN_2183 = pop_23 & empty_23 ? 1'h0 : _GEN_2170; // @[stackmanage_35.scala 5456:45 stackmanage_35.scala 5488:34]
  wire  _GEN_2184 = pop_23 & empty_23 ? 1'h0 : _GEN_2171; // @[stackmanage_35.scala 5456:45 stackmanage_35.scala 5489:34]
  wire  _GEN_2185 = pop_23 & empty_23 ? 1'h0 : _GEN_2172; // @[stackmanage_35.scala 5456:45 stackmanage_35.scala 5490:34]
  wire  _GEN_2186 = pop_23 & empty_23 ? 1'h0 : _GEN_2173; // @[stackmanage_35.scala 5456:45 stackmanage_35.scala 5491:34]
  wire  _GEN_2187 = pop_23 & empty_23 ? 1'h0 : _GEN_2174; // @[stackmanage_35.scala 5456:45 stackmanage_35.scala 5492:34]
  wire  _GEN_2190 = pop_22 & empty_22 ? 1'h0 : _T_386; // @[stackmanage_35.scala 5419:45 stackmanage_35.scala 5444:34]
  wire  _GEN_2191 = pop_22 & empty_22 ? 1'h0 : _GEN_2177; // @[stackmanage_35.scala 5419:45 stackmanage_35.scala 5445:34]
  wire  _GEN_2192 = pop_22 & empty_22 ? 1'h0 : _GEN_2178; // @[stackmanage_35.scala 5419:45 stackmanage_35.scala 5446:34]
  wire  _GEN_2193 = pop_22 & empty_22 ? 1'h0 : _GEN_2179; // @[stackmanage_35.scala 5419:45 stackmanage_35.scala 5447:34]
  wire  _GEN_2194 = pop_22 & empty_22 ? 1'h0 : _GEN_2180; // @[stackmanage_35.scala 5419:45 stackmanage_35.scala 5448:34]
  wire  _GEN_2195 = pop_22 & empty_22 ? 1'h0 : _GEN_2181; // @[stackmanage_35.scala 5419:45 stackmanage_35.scala 5449:34]
  wire  _GEN_2196 = pop_22 & empty_22 ? 1'h0 : _GEN_2182; // @[stackmanage_35.scala 5419:45 stackmanage_35.scala 5450:34]
  wire  _GEN_2197 = pop_22 & empty_22 ? 1'h0 : _GEN_2183; // @[stackmanage_35.scala 5419:45 stackmanage_35.scala 5451:34]
  wire  _GEN_2198 = pop_22 & empty_22 ? 1'h0 : _GEN_2184; // @[stackmanage_35.scala 5419:45 stackmanage_35.scala 5452:34]
  wire  _GEN_2199 = pop_22 & empty_22 ? 1'h0 : _GEN_2185; // @[stackmanage_35.scala 5419:45 stackmanage_35.scala 5453:34]
  wire  _GEN_2200 = pop_22 & empty_22 ? 1'h0 : _GEN_2186; // @[stackmanage_35.scala 5419:45 stackmanage_35.scala 5454:34]
  wire  _GEN_2201 = pop_22 & empty_22 ? 1'h0 : _GEN_2187; // @[stackmanage_35.scala 5419:45 stackmanage_35.scala 5455:34]
  wire  _GEN_2204 = pop_21 & empty_21 ? 1'h0 : _T_383; // @[stackmanage_35.scala 5382:45 stackmanage_35.scala 5406:34]
  wire  _GEN_2205 = pop_21 & empty_21 ? 1'h0 : _GEN_2190; // @[stackmanage_35.scala 5382:45 stackmanage_35.scala 5407:34]
  wire  _GEN_2206 = pop_21 & empty_21 ? 1'h0 : _GEN_2191; // @[stackmanage_35.scala 5382:45 stackmanage_35.scala 5408:34]
  wire  _GEN_2207 = pop_21 & empty_21 ? 1'h0 : _GEN_2192; // @[stackmanage_35.scala 5382:45 stackmanage_35.scala 5409:34]
  wire  _GEN_2208 = pop_21 & empty_21 ? 1'h0 : _GEN_2193; // @[stackmanage_35.scala 5382:45 stackmanage_35.scala 5410:34]
  wire  _GEN_2209 = pop_21 & empty_21 ? 1'h0 : _GEN_2194; // @[stackmanage_35.scala 5382:45 stackmanage_35.scala 5411:34]
  wire  _GEN_2210 = pop_21 & empty_21 ? 1'h0 : _GEN_2195; // @[stackmanage_35.scala 5382:45 stackmanage_35.scala 5412:34]
  wire  _GEN_2211 = pop_21 & empty_21 ? 1'h0 : _GEN_2196; // @[stackmanage_35.scala 5382:45 stackmanage_35.scala 5413:34]
  wire  _GEN_2212 = pop_21 & empty_21 ? 1'h0 : _GEN_2197; // @[stackmanage_35.scala 5382:45 stackmanage_35.scala 5414:34]
  wire  _GEN_2213 = pop_21 & empty_21 ? 1'h0 : _GEN_2198; // @[stackmanage_35.scala 5382:45 stackmanage_35.scala 5415:34]
  wire  _GEN_2214 = pop_21 & empty_21 ? 1'h0 : _GEN_2199; // @[stackmanage_35.scala 5382:45 stackmanage_35.scala 5416:34]
  wire  _GEN_2215 = pop_21 & empty_21 ? 1'h0 : _GEN_2200; // @[stackmanage_35.scala 5382:45 stackmanage_35.scala 5417:34]
  wire  _GEN_2216 = pop_21 & empty_21 ? 1'h0 : _GEN_2201; // @[stackmanage_35.scala 5382:45 stackmanage_35.scala 5418:34]
  wire  _GEN_2219 = pop_20 & empty_20 ? 1'h0 : _T_380; // @[stackmanage_35.scala 5345:45 stackmanage_35.scala 5368:34]
  wire  _GEN_2220 = pop_20 & empty_20 ? 1'h0 : _GEN_2204; // @[stackmanage_35.scala 5345:45 stackmanage_35.scala 5369:34]
  wire  _GEN_2221 = pop_20 & empty_20 ? 1'h0 : _GEN_2205; // @[stackmanage_35.scala 5345:45 stackmanage_35.scala 5370:34]
  wire  _GEN_2222 = pop_20 & empty_20 ? 1'h0 : _GEN_2206; // @[stackmanage_35.scala 5345:45 stackmanage_35.scala 5371:34]
  wire  _GEN_2223 = pop_20 & empty_20 ? 1'h0 : _GEN_2207; // @[stackmanage_35.scala 5345:45 stackmanage_35.scala 5372:34]
  wire  _GEN_2224 = pop_20 & empty_20 ? 1'h0 : _GEN_2208; // @[stackmanage_35.scala 5345:45 stackmanage_35.scala 5373:34]
  wire  _GEN_2225 = pop_20 & empty_20 ? 1'h0 : _GEN_2209; // @[stackmanage_35.scala 5345:45 stackmanage_35.scala 5374:34]
  wire  _GEN_2226 = pop_20 & empty_20 ? 1'h0 : _GEN_2210; // @[stackmanage_35.scala 5345:45 stackmanage_35.scala 5375:34]
  wire  _GEN_2227 = pop_20 & empty_20 ? 1'h0 : _GEN_2211; // @[stackmanage_35.scala 5345:45 stackmanage_35.scala 5376:34]
  wire  _GEN_2228 = pop_20 & empty_20 ? 1'h0 : _GEN_2212; // @[stackmanage_35.scala 5345:45 stackmanage_35.scala 5377:34]
  wire  _GEN_2229 = pop_20 & empty_20 ? 1'h0 : _GEN_2213; // @[stackmanage_35.scala 5345:45 stackmanage_35.scala 5378:34]
  wire  _GEN_2230 = pop_20 & empty_20 ? 1'h0 : _GEN_2214; // @[stackmanage_35.scala 5345:45 stackmanage_35.scala 5379:34]
  wire  _GEN_2231 = pop_20 & empty_20 ? 1'h0 : _GEN_2215; // @[stackmanage_35.scala 5345:45 stackmanage_35.scala 5380:34]
  wire  _GEN_2232 = pop_20 & empty_20 ? 1'h0 : _GEN_2216; // @[stackmanage_35.scala 5345:45 stackmanage_35.scala 5381:34]
  wire  _GEN_2235 = pop_19 & empty_19 ? 1'h0 : _T_377; // @[stackmanage_35.scala 5308:45 stackmanage_35.scala 5330:34]
  wire  _GEN_2236 = pop_19 & empty_19 ? 1'h0 : _GEN_2219; // @[stackmanage_35.scala 5308:45 stackmanage_35.scala 5331:34]
  wire  _GEN_2237 = pop_19 & empty_19 ? 1'h0 : _GEN_2220; // @[stackmanage_35.scala 5308:45 stackmanage_35.scala 5332:34]
  wire  _GEN_2238 = pop_19 & empty_19 ? 1'h0 : _GEN_2221; // @[stackmanage_35.scala 5308:45 stackmanage_35.scala 5333:34]
  wire  _GEN_2239 = pop_19 & empty_19 ? 1'h0 : _GEN_2222; // @[stackmanage_35.scala 5308:45 stackmanage_35.scala 5334:34]
  wire  _GEN_2240 = pop_19 & empty_19 ? 1'h0 : _GEN_2223; // @[stackmanage_35.scala 5308:45 stackmanage_35.scala 5335:34]
  wire  _GEN_2241 = pop_19 & empty_19 ? 1'h0 : _GEN_2224; // @[stackmanage_35.scala 5308:45 stackmanage_35.scala 5336:34]
  wire  _GEN_2242 = pop_19 & empty_19 ? 1'h0 : _GEN_2225; // @[stackmanage_35.scala 5308:45 stackmanage_35.scala 5337:34]
  wire  _GEN_2243 = pop_19 & empty_19 ? 1'h0 : _GEN_2226; // @[stackmanage_35.scala 5308:45 stackmanage_35.scala 5338:34]
  wire  _GEN_2244 = pop_19 & empty_19 ? 1'h0 : _GEN_2227; // @[stackmanage_35.scala 5308:45 stackmanage_35.scala 5339:34]
  wire  _GEN_2245 = pop_19 & empty_19 ? 1'h0 : _GEN_2228; // @[stackmanage_35.scala 5308:45 stackmanage_35.scala 5340:34]
  wire  _GEN_2246 = pop_19 & empty_19 ? 1'h0 : _GEN_2229; // @[stackmanage_35.scala 5308:45 stackmanage_35.scala 5341:34]
  wire  _GEN_2247 = pop_19 & empty_19 ? 1'h0 : _GEN_2230; // @[stackmanage_35.scala 5308:45 stackmanage_35.scala 5342:34]
  wire  _GEN_2248 = pop_19 & empty_19 ? 1'h0 : _GEN_2231; // @[stackmanage_35.scala 5308:45 stackmanage_35.scala 5343:34]
  wire  _GEN_2249 = pop_19 & empty_19 ? 1'h0 : _GEN_2232; // @[stackmanage_35.scala 5308:45 stackmanage_35.scala 5344:34]
  wire  _GEN_2252 = pop_18 & empty_18 ? 1'h0 : _T_374; // @[stackmanage_35.scala 5271:45 stackmanage_35.scala 5292:34]
  wire  _GEN_2253 = pop_18 & empty_18 ? 1'h0 : _GEN_2235; // @[stackmanage_35.scala 5271:45 stackmanage_35.scala 5293:34]
  wire  _GEN_2254 = pop_18 & empty_18 ? 1'h0 : _GEN_2236; // @[stackmanage_35.scala 5271:45 stackmanage_35.scala 5294:34]
  wire  _GEN_2255 = pop_18 & empty_18 ? 1'h0 : _GEN_2237; // @[stackmanage_35.scala 5271:45 stackmanage_35.scala 5295:34]
  wire  _GEN_2256 = pop_18 & empty_18 ? 1'h0 : _GEN_2238; // @[stackmanage_35.scala 5271:45 stackmanage_35.scala 5296:34]
  wire  _GEN_2257 = pop_18 & empty_18 ? 1'h0 : _GEN_2239; // @[stackmanage_35.scala 5271:45 stackmanage_35.scala 5297:34]
  wire  _GEN_2258 = pop_18 & empty_18 ? 1'h0 : _GEN_2240; // @[stackmanage_35.scala 5271:45 stackmanage_35.scala 5298:34]
  wire  _GEN_2259 = pop_18 & empty_18 ? 1'h0 : _GEN_2241; // @[stackmanage_35.scala 5271:45 stackmanage_35.scala 5299:34]
  wire  _GEN_2260 = pop_18 & empty_18 ? 1'h0 : _GEN_2242; // @[stackmanage_35.scala 5271:45 stackmanage_35.scala 5300:34]
  wire  _GEN_2261 = pop_18 & empty_18 ? 1'h0 : _GEN_2243; // @[stackmanage_35.scala 5271:45 stackmanage_35.scala 5301:34]
  wire  _GEN_2262 = pop_18 & empty_18 ? 1'h0 : _GEN_2244; // @[stackmanage_35.scala 5271:45 stackmanage_35.scala 5302:34]
  wire  _GEN_2263 = pop_18 & empty_18 ? 1'h0 : _GEN_2245; // @[stackmanage_35.scala 5271:45 stackmanage_35.scala 5303:34]
  wire  _GEN_2264 = pop_18 & empty_18 ? 1'h0 : _GEN_2246; // @[stackmanage_35.scala 5271:45 stackmanage_35.scala 5304:34]
  wire  _GEN_2265 = pop_18 & empty_18 ? 1'h0 : _GEN_2247; // @[stackmanage_35.scala 5271:45 stackmanage_35.scala 5305:34]
  wire  _GEN_2266 = pop_18 & empty_18 ? 1'h0 : _GEN_2248; // @[stackmanage_35.scala 5271:45 stackmanage_35.scala 5306:34]
  wire  _GEN_2267 = pop_18 & empty_18 ? 1'h0 : _GEN_2249; // @[stackmanage_35.scala 5271:45 stackmanage_35.scala 5307:34]
  wire  _GEN_2270 = pop_17 & empty_17 ? 1'h0 : _T_371; // @[stackmanage_35.scala 5234:45 stackmanage_35.scala 5254:34]
  wire  _GEN_2271 = pop_17 & empty_17 ? 1'h0 : _GEN_2252; // @[stackmanage_35.scala 5234:45 stackmanage_35.scala 5255:34]
  wire  _GEN_2272 = pop_17 & empty_17 ? 1'h0 : _GEN_2253; // @[stackmanage_35.scala 5234:45 stackmanage_35.scala 5256:34]
  wire  _GEN_2273 = pop_17 & empty_17 ? 1'h0 : _GEN_2254; // @[stackmanage_35.scala 5234:45 stackmanage_35.scala 5257:34]
  wire  _GEN_2274 = pop_17 & empty_17 ? 1'h0 : _GEN_2255; // @[stackmanage_35.scala 5234:45 stackmanage_35.scala 5258:34]
  wire  _GEN_2275 = pop_17 & empty_17 ? 1'h0 : _GEN_2256; // @[stackmanage_35.scala 5234:45 stackmanage_35.scala 5259:34]
  wire  _GEN_2276 = pop_17 & empty_17 ? 1'h0 : _GEN_2257; // @[stackmanage_35.scala 5234:45 stackmanage_35.scala 5260:34]
  wire  _GEN_2277 = pop_17 & empty_17 ? 1'h0 : _GEN_2258; // @[stackmanage_35.scala 5234:45 stackmanage_35.scala 5261:34]
  wire  _GEN_2278 = pop_17 & empty_17 ? 1'h0 : _GEN_2259; // @[stackmanage_35.scala 5234:45 stackmanage_35.scala 5262:34]
  wire  _GEN_2279 = pop_17 & empty_17 ? 1'h0 : _GEN_2260; // @[stackmanage_35.scala 5234:45 stackmanage_35.scala 5263:34]
  wire  _GEN_2280 = pop_17 & empty_17 ? 1'h0 : _GEN_2261; // @[stackmanage_35.scala 5234:45 stackmanage_35.scala 5264:34]
  wire  _GEN_2281 = pop_17 & empty_17 ? 1'h0 : _GEN_2262; // @[stackmanage_35.scala 5234:45 stackmanage_35.scala 5265:34]
  wire  _GEN_2282 = pop_17 & empty_17 ? 1'h0 : _GEN_2263; // @[stackmanage_35.scala 5234:45 stackmanage_35.scala 5266:34]
  wire  _GEN_2283 = pop_17 & empty_17 ? 1'h0 : _GEN_2264; // @[stackmanage_35.scala 5234:45 stackmanage_35.scala 5267:34]
  wire  _GEN_2284 = pop_17 & empty_17 ? 1'h0 : _GEN_2265; // @[stackmanage_35.scala 5234:45 stackmanage_35.scala 5268:34]
  wire  _GEN_2285 = pop_17 & empty_17 ? 1'h0 : _GEN_2266; // @[stackmanage_35.scala 5234:45 stackmanage_35.scala 5269:34]
  wire  _GEN_2286 = pop_17 & empty_17 ? 1'h0 : _GEN_2267; // @[stackmanage_35.scala 5234:45 stackmanage_35.scala 5270:34]
  wire  _GEN_2289 = pop_16 & empty_16 ? 1'h0 : _T_368; // @[stackmanage_35.scala 5197:45 stackmanage_35.scala 5216:34]
  wire  _GEN_2290 = pop_16 & empty_16 ? 1'h0 : _GEN_2270; // @[stackmanage_35.scala 5197:45 stackmanage_35.scala 5217:34]
  wire  _GEN_2291 = pop_16 & empty_16 ? 1'h0 : _GEN_2271; // @[stackmanage_35.scala 5197:45 stackmanage_35.scala 5218:34]
  wire  _GEN_2292 = pop_16 & empty_16 ? 1'h0 : _GEN_2272; // @[stackmanage_35.scala 5197:45 stackmanage_35.scala 5219:34]
  wire  _GEN_2293 = pop_16 & empty_16 ? 1'h0 : _GEN_2273; // @[stackmanage_35.scala 5197:45 stackmanage_35.scala 5220:34]
  wire  _GEN_2294 = pop_16 & empty_16 ? 1'h0 : _GEN_2274; // @[stackmanage_35.scala 5197:45 stackmanage_35.scala 5221:34]
  wire  _GEN_2295 = pop_16 & empty_16 ? 1'h0 : _GEN_2275; // @[stackmanage_35.scala 5197:45 stackmanage_35.scala 5222:34]
  wire  _GEN_2296 = pop_16 & empty_16 ? 1'h0 : _GEN_2276; // @[stackmanage_35.scala 5197:45 stackmanage_35.scala 5223:34]
  wire  _GEN_2297 = pop_16 & empty_16 ? 1'h0 : _GEN_2277; // @[stackmanage_35.scala 5197:45 stackmanage_35.scala 5224:34]
  wire  _GEN_2298 = pop_16 & empty_16 ? 1'h0 : _GEN_2278; // @[stackmanage_35.scala 5197:45 stackmanage_35.scala 5225:34]
  wire  _GEN_2299 = pop_16 & empty_16 ? 1'h0 : _GEN_2279; // @[stackmanage_35.scala 5197:45 stackmanage_35.scala 5226:34]
  wire  _GEN_2300 = pop_16 & empty_16 ? 1'h0 : _GEN_2280; // @[stackmanage_35.scala 5197:45 stackmanage_35.scala 5227:34]
  wire  _GEN_2301 = pop_16 & empty_16 ? 1'h0 : _GEN_2281; // @[stackmanage_35.scala 5197:45 stackmanage_35.scala 5228:34]
  wire  _GEN_2302 = pop_16 & empty_16 ? 1'h0 : _GEN_2282; // @[stackmanage_35.scala 5197:45 stackmanage_35.scala 5229:34]
  wire  _GEN_2303 = pop_16 & empty_16 ? 1'h0 : _GEN_2283; // @[stackmanage_35.scala 5197:45 stackmanage_35.scala 5230:34]
  wire  _GEN_2304 = pop_16 & empty_16 ? 1'h0 : _GEN_2284; // @[stackmanage_35.scala 5197:45 stackmanage_35.scala 5231:34]
  wire  _GEN_2305 = pop_16 & empty_16 ? 1'h0 : _GEN_2285; // @[stackmanage_35.scala 5197:45 stackmanage_35.scala 5232:34]
  wire  _GEN_2306 = pop_16 & empty_16 ? 1'h0 : _GEN_2286; // @[stackmanage_35.scala 5197:45 stackmanage_35.scala 5233:34]
  wire  _GEN_2309 = pop_15 & empty_15 ? 1'h0 : _T_365; // @[stackmanage_35.scala 5160:45 stackmanage_35.scala 5178:34]
  wire  _GEN_2310 = pop_15 & empty_15 ? 1'h0 : _GEN_2289; // @[stackmanage_35.scala 5160:45 stackmanage_35.scala 5179:34]
  wire  _GEN_2311 = pop_15 & empty_15 ? 1'h0 : _GEN_2290; // @[stackmanage_35.scala 5160:45 stackmanage_35.scala 5180:34]
  wire  _GEN_2312 = pop_15 & empty_15 ? 1'h0 : _GEN_2291; // @[stackmanage_35.scala 5160:45 stackmanage_35.scala 5181:34]
  wire  _GEN_2313 = pop_15 & empty_15 ? 1'h0 : _GEN_2292; // @[stackmanage_35.scala 5160:45 stackmanage_35.scala 5182:34]
  wire  _GEN_2314 = pop_15 & empty_15 ? 1'h0 : _GEN_2293; // @[stackmanage_35.scala 5160:45 stackmanage_35.scala 5183:34]
  wire  _GEN_2315 = pop_15 & empty_15 ? 1'h0 : _GEN_2294; // @[stackmanage_35.scala 5160:45 stackmanage_35.scala 5184:34]
  wire  _GEN_2316 = pop_15 & empty_15 ? 1'h0 : _GEN_2295; // @[stackmanage_35.scala 5160:45 stackmanage_35.scala 5185:34]
  wire  _GEN_2317 = pop_15 & empty_15 ? 1'h0 : _GEN_2296; // @[stackmanage_35.scala 5160:45 stackmanage_35.scala 5186:34]
  wire  _GEN_2318 = pop_15 & empty_15 ? 1'h0 : _GEN_2297; // @[stackmanage_35.scala 5160:45 stackmanage_35.scala 5187:34]
  wire  _GEN_2319 = pop_15 & empty_15 ? 1'h0 : _GEN_2298; // @[stackmanage_35.scala 5160:45 stackmanage_35.scala 5188:34]
  wire  _GEN_2320 = pop_15 & empty_15 ? 1'h0 : _GEN_2299; // @[stackmanage_35.scala 5160:45 stackmanage_35.scala 5189:34]
  wire  _GEN_2321 = pop_15 & empty_15 ? 1'h0 : _GEN_2300; // @[stackmanage_35.scala 5160:45 stackmanage_35.scala 5190:34]
  wire  _GEN_2322 = pop_15 & empty_15 ? 1'h0 : _GEN_2301; // @[stackmanage_35.scala 5160:45 stackmanage_35.scala 5191:34]
  wire  _GEN_2323 = pop_15 & empty_15 ? 1'h0 : _GEN_2302; // @[stackmanage_35.scala 5160:45 stackmanage_35.scala 5192:34]
  wire  _GEN_2324 = pop_15 & empty_15 ? 1'h0 : _GEN_2303; // @[stackmanage_35.scala 5160:45 stackmanage_35.scala 5193:34]
  wire  _GEN_2325 = pop_15 & empty_15 ? 1'h0 : _GEN_2304; // @[stackmanage_35.scala 5160:45 stackmanage_35.scala 5194:34]
  wire  _GEN_2326 = pop_15 & empty_15 ? 1'h0 : _GEN_2305; // @[stackmanage_35.scala 5160:45 stackmanage_35.scala 5195:34]
  wire  _GEN_2327 = pop_15 & empty_15 ? 1'h0 : _GEN_2306; // @[stackmanage_35.scala 5160:45 stackmanage_35.scala 5196:34]
  wire  _GEN_2330 = pop_14 & empty_14 ? 1'h0 : _T_362; // @[stackmanage_35.scala 5123:45 stackmanage_35.scala 5140:34]
  wire  _GEN_2331 = pop_14 & empty_14 ? 1'h0 : _GEN_2309; // @[stackmanage_35.scala 5123:45 stackmanage_35.scala 5141:34]
  wire  _GEN_2332 = pop_14 & empty_14 ? 1'h0 : _GEN_2310; // @[stackmanage_35.scala 5123:45 stackmanage_35.scala 5142:34]
  wire  _GEN_2333 = pop_14 & empty_14 ? 1'h0 : _GEN_2311; // @[stackmanage_35.scala 5123:45 stackmanage_35.scala 5143:34]
  wire  _GEN_2334 = pop_14 & empty_14 ? 1'h0 : _GEN_2312; // @[stackmanage_35.scala 5123:45 stackmanage_35.scala 5144:34]
  wire  _GEN_2335 = pop_14 & empty_14 ? 1'h0 : _GEN_2313; // @[stackmanage_35.scala 5123:45 stackmanage_35.scala 5145:34]
  wire  _GEN_2336 = pop_14 & empty_14 ? 1'h0 : _GEN_2314; // @[stackmanage_35.scala 5123:45 stackmanage_35.scala 5146:34]
  wire  _GEN_2337 = pop_14 & empty_14 ? 1'h0 : _GEN_2315; // @[stackmanage_35.scala 5123:45 stackmanage_35.scala 5147:34]
  wire  _GEN_2338 = pop_14 & empty_14 ? 1'h0 : _GEN_2316; // @[stackmanage_35.scala 5123:45 stackmanage_35.scala 5148:34]
  wire  _GEN_2339 = pop_14 & empty_14 ? 1'h0 : _GEN_2317; // @[stackmanage_35.scala 5123:45 stackmanage_35.scala 5149:34]
  wire  _GEN_2340 = pop_14 & empty_14 ? 1'h0 : _GEN_2318; // @[stackmanage_35.scala 5123:45 stackmanage_35.scala 5150:34]
  wire  _GEN_2341 = pop_14 & empty_14 ? 1'h0 : _GEN_2319; // @[stackmanage_35.scala 5123:45 stackmanage_35.scala 5151:34]
  wire  _GEN_2342 = pop_14 & empty_14 ? 1'h0 : _GEN_2320; // @[stackmanage_35.scala 5123:45 stackmanage_35.scala 5152:34]
  wire  _GEN_2343 = pop_14 & empty_14 ? 1'h0 : _GEN_2321; // @[stackmanage_35.scala 5123:45 stackmanage_35.scala 5153:34]
  wire  _GEN_2344 = pop_14 & empty_14 ? 1'h0 : _GEN_2322; // @[stackmanage_35.scala 5123:45 stackmanage_35.scala 5154:34]
  wire  _GEN_2345 = pop_14 & empty_14 ? 1'h0 : _GEN_2323; // @[stackmanage_35.scala 5123:45 stackmanage_35.scala 5155:34]
  wire  _GEN_2346 = pop_14 & empty_14 ? 1'h0 : _GEN_2324; // @[stackmanage_35.scala 5123:45 stackmanage_35.scala 5156:34]
  wire  _GEN_2347 = pop_14 & empty_14 ? 1'h0 : _GEN_2325; // @[stackmanage_35.scala 5123:45 stackmanage_35.scala 5157:34]
  wire  _GEN_2348 = pop_14 & empty_14 ? 1'h0 : _GEN_2326; // @[stackmanage_35.scala 5123:45 stackmanage_35.scala 5158:34]
  wire  _GEN_2349 = pop_14 & empty_14 ? 1'h0 : _GEN_2327; // @[stackmanage_35.scala 5123:45 stackmanage_35.scala 5159:34]
  wire  _GEN_2352 = pop_13 & empty_13 ? 1'h0 : _T_359; // @[stackmanage_35.scala 5086:45 stackmanage_35.scala 5102:34]
  wire  _GEN_2353 = pop_13 & empty_13 ? 1'h0 : _GEN_2330; // @[stackmanage_35.scala 5086:45 stackmanage_35.scala 5103:34]
  wire  _GEN_2354 = pop_13 & empty_13 ? 1'h0 : _GEN_2331; // @[stackmanage_35.scala 5086:45 stackmanage_35.scala 5104:34]
  wire  _GEN_2355 = pop_13 & empty_13 ? 1'h0 : _GEN_2332; // @[stackmanage_35.scala 5086:45 stackmanage_35.scala 5105:34]
  wire  _GEN_2356 = pop_13 & empty_13 ? 1'h0 : _GEN_2333; // @[stackmanage_35.scala 5086:45 stackmanage_35.scala 5106:34]
  wire  _GEN_2357 = pop_13 & empty_13 ? 1'h0 : _GEN_2334; // @[stackmanage_35.scala 5086:45 stackmanage_35.scala 5107:34]
  wire  _GEN_2358 = pop_13 & empty_13 ? 1'h0 : _GEN_2335; // @[stackmanage_35.scala 5086:45 stackmanage_35.scala 5108:34]
  wire  _GEN_2359 = pop_13 & empty_13 ? 1'h0 : _GEN_2336; // @[stackmanage_35.scala 5086:45 stackmanage_35.scala 5109:34]
  wire  _GEN_2360 = pop_13 & empty_13 ? 1'h0 : _GEN_2337; // @[stackmanage_35.scala 5086:45 stackmanage_35.scala 5110:34]
  wire  _GEN_2361 = pop_13 & empty_13 ? 1'h0 : _GEN_2338; // @[stackmanage_35.scala 5086:45 stackmanage_35.scala 5111:34]
  wire  _GEN_2362 = pop_13 & empty_13 ? 1'h0 : _GEN_2339; // @[stackmanage_35.scala 5086:45 stackmanage_35.scala 5112:34]
  wire  _GEN_2363 = pop_13 & empty_13 ? 1'h0 : _GEN_2340; // @[stackmanage_35.scala 5086:45 stackmanage_35.scala 5113:34]
  wire  _GEN_2364 = pop_13 & empty_13 ? 1'h0 : _GEN_2341; // @[stackmanage_35.scala 5086:45 stackmanage_35.scala 5114:34]
  wire  _GEN_2365 = pop_13 & empty_13 ? 1'h0 : _GEN_2342; // @[stackmanage_35.scala 5086:45 stackmanage_35.scala 5115:34]
  wire  _GEN_2366 = pop_13 & empty_13 ? 1'h0 : _GEN_2343; // @[stackmanage_35.scala 5086:45 stackmanage_35.scala 5116:34]
  wire  _GEN_2367 = pop_13 & empty_13 ? 1'h0 : _GEN_2344; // @[stackmanage_35.scala 5086:45 stackmanage_35.scala 5117:34]
  wire  _GEN_2368 = pop_13 & empty_13 ? 1'h0 : _GEN_2345; // @[stackmanage_35.scala 5086:45 stackmanage_35.scala 5118:34]
  wire  _GEN_2369 = pop_13 & empty_13 ? 1'h0 : _GEN_2346; // @[stackmanage_35.scala 5086:45 stackmanage_35.scala 5119:34]
  wire  _GEN_2370 = pop_13 & empty_13 ? 1'h0 : _GEN_2347; // @[stackmanage_35.scala 5086:45 stackmanage_35.scala 5120:34]
  wire  _GEN_2371 = pop_13 & empty_13 ? 1'h0 : _GEN_2348; // @[stackmanage_35.scala 5086:45 stackmanage_35.scala 5121:34]
  wire  _GEN_2372 = pop_13 & empty_13 ? 1'h0 : _GEN_2349; // @[stackmanage_35.scala 5086:45 stackmanage_35.scala 5122:34]
  wire  _GEN_2375 = pop_12 & empty_12 ? 1'h0 : _T_356; // @[stackmanage_35.scala 5049:45 stackmanage_35.scala 5064:34]
  wire  _GEN_2376 = pop_12 & empty_12 ? 1'h0 : _GEN_2352; // @[stackmanage_35.scala 5049:45 stackmanage_35.scala 5065:34]
  wire  _GEN_2377 = pop_12 & empty_12 ? 1'h0 : _GEN_2353; // @[stackmanage_35.scala 5049:45 stackmanage_35.scala 5066:34]
  wire  _GEN_2378 = pop_12 & empty_12 ? 1'h0 : _GEN_2354; // @[stackmanage_35.scala 5049:45 stackmanage_35.scala 5067:34]
  wire  _GEN_2379 = pop_12 & empty_12 ? 1'h0 : _GEN_2355; // @[stackmanage_35.scala 5049:45 stackmanage_35.scala 5068:34]
  wire  _GEN_2380 = pop_12 & empty_12 ? 1'h0 : _GEN_2356; // @[stackmanage_35.scala 5049:45 stackmanage_35.scala 5069:34]
  wire  _GEN_2381 = pop_12 & empty_12 ? 1'h0 : _GEN_2357; // @[stackmanage_35.scala 5049:45 stackmanage_35.scala 5070:34]
  wire  _GEN_2382 = pop_12 & empty_12 ? 1'h0 : _GEN_2358; // @[stackmanage_35.scala 5049:45 stackmanage_35.scala 5071:34]
  wire  _GEN_2383 = pop_12 & empty_12 ? 1'h0 : _GEN_2359; // @[stackmanage_35.scala 5049:45 stackmanage_35.scala 5072:34]
  wire  _GEN_2384 = pop_12 & empty_12 ? 1'h0 : _GEN_2360; // @[stackmanage_35.scala 5049:45 stackmanage_35.scala 5073:34]
  wire  _GEN_2385 = pop_12 & empty_12 ? 1'h0 : _GEN_2361; // @[stackmanage_35.scala 5049:45 stackmanage_35.scala 5074:34]
  wire  _GEN_2386 = pop_12 & empty_12 ? 1'h0 : _GEN_2362; // @[stackmanage_35.scala 5049:45 stackmanage_35.scala 5075:34]
  wire  _GEN_2387 = pop_12 & empty_12 ? 1'h0 : _GEN_2363; // @[stackmanage_35.scala 5049:45 stackmanage_35.scala 5076:34]
  wire  _GEN_2388 = pop_12 & empty_12 ? 1'h0 : _GEN_2364; // @[stackmanage_35.scala 5049:45 stackmanage_35.scala 5077:34]
  wire  _GEN_2389 = pop_12 & empty_12 ? 1'h0 : _GEN_2365; // @[stackmanage_35.scala 5049:45 stackmanage_35.scala 5078:34]
  wire  _GEN_2390 = pop_12 & empty_12 ? 1'h0 : _GEN_2366; // @[stackmanage_35.scala 5049:45 stackmanage_35.scala 5079:34]
  wire  _GEN_2391 = pop_12 & empty_12 ? 1'h0 : _GEN_2367; // @[stackmanage_35.scala 5049:45 stackmanage_35.scala 5080:34]
  wire  _GEN_2392 = pop_12 & empty_12 ? 1'h0 : _GEN_2368; // @[stackmanage_35.scala 5049:45 stackmanage_35.scala 5081:34]
  wire  _GEN_2393 = pop_12 & empty_12 ? 1'h0 : _GEN_2369; // @[stackmanage_35.scala 5049:45 stackmanage_35.scala 5082:34]
  wire  _GEN_2394 = pop_12 & empty_12 ? 1'h0 : _GEN_2370; // @[stackmanage_35.scala 5049:45 stackmanage_35.scala 5083:34]
  wire  _GEN_2395 = pop_12 & empty_12 ? 1'h0 : _GEN_2371; // @[stackmanage_35.scala 5049:45 stackmanage_35.scala 5084:34]
  wire  _GEN_2396 = pop_12 & empty_12 ? 1'h0 : _GEN_2372; // @[stackmanage_35.scala 5049:45 stackmanage_35.scala 5085:34]
  wire  _GEN_2399 = pop_11 & empty_11 ? 1'h0 : _T_353; // @[stackmanage_35.scala 5012:45 stackmanage_35.scala 5026:34]
  wire  _GEN_2400 = pop_11 & empty_11 ? 1'h0 : _GEN_2375; // @[stackmanage_35.scala 5012:45 stackmanage_35.scala 5027:34]
  wire  _GEN_2401 = pop_11 & empty_11 ? 1'h0 : _GEN_2376; // @[stackmanage_35.scala 5012:45 stackmanage_35.scala 5028:34]
  wire  _GEN_2402 = pop_11 & empty_11 ? 1'h0 : _GEN_2377; // @[stackmanage_35.scala 5012:45 stackmanage_35.scala 5029:34]
  wire  _GEN_2403 = pop_11 & empty_11 ? 1'h0 : _GEN_2378; // @[stackmanage_35.scala 5012:45 stackmanage_35.scala 5030:34]
  wire  _GEN_2404 = pop_11 & empty_11 ? 1'h0 : _GEN_2379; // @[stackmanage_35.scala 5012:45 stackmanage_35.scala 5031:34]
  wire  _GEN_2405 = pop_11 & empty_11 ? 1'h0 : _GEN_2380; // @[stackmanage_35.scala 5012:45 stackmanage_35.scala 5032:34]
  wire  _GEN_2406 = pop_11 & empty_11 ? 1'h0 : _GEN_2381; // @[stackmanage_35.scala 5012:45 stackmanage_35.scala 5033:34]
  wire  _GEN_2407 = pop_11 & empty_11 ? 1'h0 : _GEN_2382; // @[stackmanage_35.scala 5012:45 stackmanage_35.scala 5034:34]
  wire  _GEN_2408 = pop_11 & empty_11 ? 1'h0 : _GEN_2383; // @[stackmanage_35.scala 5012:45 stackmanage_35.scala 5035:34]
  wire  _GEN_2409 = pop_11 & empty_11 ? 1'h0 : _GEN_2384; // @[stackmanage_35.scala 5012:45 stackmanage_35.scala 5036:34]
  wire  _GEN_2410 = pop_11 & empty_11 ? 1'h0 : _GEN_2385; // @[stackmanage_35.scala 5012:45 stackmanage_35.scala 5037:34]
  wire  _GEN_2411 = pop_11 & empty_11 ? 1'h0 : _GEN_2386; // @[stackmanage_35.scala 5012:45 stackmanage_35.scala 5038:34]
  wire  _GEN_2412 = pop_11 & empty_11 ? 1'h0 : _GEN_2387; // @[stackmanage_35.scala 5012:45 stackmanage_35.scala 5039:34]
  wire  _GEN_2413 = pop_11 & empty_11 ? 1'h0 : _GEN_2388; // @[stackmanage_35.scala 5012:45 stackmanage_35.scala 5040:34]
  wire  _GEN_2414 = pop_11 & empty_11 ? 1'h0 : _GEN_2389; // @[stackmanage_35.scala 5012:45 stackmanage_35.scala 5041:34]
  wire  _GEN_2415 = pop_11 & empty_11 ? 1'h0 : _GEN_2390; // @[stackmanage_35.scala 5012:45 stackmanage_35.scala 5042:34]
  wire  _GEN_2416 = pop_11 & empty_11 ? 1'h0 : _GEN_2391; // @[stackmanage_35.scala 5012:45 stackmanage_35.scala 5043:34]
  wire  _GEN_2417 = pop_11 & empty_11 ? 1'h0 : _GEN_2392; // @[stackmanage_35.scala 5012:45 stackmanage_35.scala 5044:34]
  wire  _GEN_2418 = pop_11 & empty_11 ? 1'h0 : _GEN_2393; // @[stackmanage_35.scala 5012:45 stackmanage_35.scala 5045:34]
  wire  _GEN_2419 = pop_11 & empty_11 ? 1'h0 : _GEN_2394; // @[stackmanage_35.scala 5012:45 stackmanage_35.scala 5046:34]
  wire  _GEN_2420 = pop_11 & empty_11 ? 1'h0 : _GEN_2395; // @[stackmanage_35.scala 5012:45 stackmanage_35.scala 5047:34]
  wire  _GEN_2421 = pop_11 & empty_11 ? 1'h0 : _GEN_2396; // @[stackmanage_35.scala 5012:45 stackmanage_35.scala 5048:34]
  wire  _GEN_2424 = pop_10 & empty_10 ? 1'h0 : _T_350; // @[stackmanage_35.scala 4975:45 stackmanage_35.scala 4988:34]
  wire  _GEN_2425 = pop_10 & empty_10 ? 1'h0 : _GEN_2399; // @[stackmanage_35.scala 4975:45 stackmanage_35.scala 4989:34]
  wire  _GEN_2426 = pop_10 & empty_10 ? 1'h0 : _GEN_2400; // @[stackmanage_35.scala 4975:45 stackmanage_35.scala 4990:34]
  wire  _GEN_2427 = pop_10 & empty_10 ? 1'h0 : _GEN_2401; // @[stackmanage_35.scala 4975:45 stackmanage_35.scala 4991:34]
  wire  _GEN_2428 = pop_10 & empty_10 ? 1'h0 : _GEN_2402; // @[stackmanage_35.scala 4975:45 stackmanage_35.scala 4992:34]
  wire  _GEN_2429 = pop_10 & empty_10 ? 1'h0 : _GEN_2403; // @[stackmanage_35.scala 4975:45 stackmanage_35.scala 4993:34]
  wire  _GEN_2430 = pop_10 & empty_10 ? 1'h0 : _GEN_2404; // @[stackmanage_35.scala 4975:45 stackmanage_35.scala 4994:34]
  wire  _GEN_2431 = pop_10 & empty_10 ? 1'h0 : _GEN_2405; // @[stackmanage_35.scala 4975:45 stackmanage_35.scala 4995:34]
  wire  _GEN_2432 = pop_10 & empty_10 ? 1'h0 : _GEN_2406; // @[stackmanage_35.scala 4975:45 stackmanage_35.scala 4996:34]
  wire  _GEN_2433 = pop_10 & empty_10 ? 1'h0 : _GEN_2407; // @[stackmanage_35.scala 4975:45 stackmanage_35.scala 4997:34]
  wire  _GEN_2434 = pop_10 & empty_10 ? 1'h0 : _GEN_2408; // @[stackmanage_35.scala 4975:45 stackmanage_35.scala 4998:34]
  wire  _GEN_2435 = pop_10 & empty_10 ? 1'h0 : _GEN_2409; // @[stackmanage_35.scala 4975:45 stackmanage_35.scala 4999:34]
  wire  _GEN_2436 = pop_10 & empty_10 ? 1'h0 : _GEN_2410; // @[stackmanage_35.scala 4975:45 stackmanage_35.scala 5000:34]
  wire  _GEN_2437 = pop_10 & empty_10 ? 1'h0 : _GEN_2411; // @[stackmanage_35.scala 4975:45 stackmanage_35.scala 5001:34]
  wire  _GEN_2438 = pop_10 & empty_10 ? 1'h0 : _GEN_2412; // @[stackmanage_35.scala 4975:45 stackmanage_35.scala 5002:34]
  wire  _GEN_2439 = pop_10 & empty_10 ? 1'h0 : _GEN_2413; // @[stackmanage_35.scala 4975:45 stackmanage_35.scala 5003:34]
  wire  _GEN_2440 = pop_10 & empty_10 ? 1'h0 : _GEN_2414; // @[stackmanage_35.scala 4975:45 stackmanage_35.scala 5004:34]
  wire  _GEN_2441 = pop_10 & empty_10 ? 1'h0 : _GEN_2415; // @[stackmanage_35.scala 4975:45 stackmanage_35.scala 5005:34]
  wire  _GEN_2442 = pop_10 & empty_10 ? 1'h0 : _GEN_2416; // @[stackmanage_35.scala 4975:45 stackmanage_35.scala 5006:34]
  wire  _GEN_2443 = pop_10 & empty_10 ? 1'h0 : _GEN_2417; // @[stackmanage_35.scala 4975:45 stackmanage_35.scala 5007:34]
  wire  _GEN_2444 = pop_10 & empty_10 ? 1'h0 : _GEN_2418; // @[stackmanage_35.scala 4975:45 stackmanage_35.scala 5008:34]
  wire  _GEN_2445 = pop_10 & empty_10 ? 1'h0 : _GEN_2419; // @[stackmanage_35.scala 4975:45 stackmanage_35.scala 5009:34]
  wire  _GEN_2446 = pop_10 & empty_10 ? 1'h0 : _GEN_2420; // @[stackmanage_35.scala 4975:45 stackmanage_35.scala 5010:34]
  wire  _GEN_2447 = pop_10 & empty_10 ? 1'h0 : _GEN_2421; // @[stackmanage_35.scala 4975:45 stackmanage_35.scala 5011:34]
  wire  _GEN_2450 = pop_9 & empty_9 ? 1'h0 : _T_347; // @[stackmanage_35.scala 4937:43 stackmanage_35.scala 4949:34]
  wire  _GEN_2451 = pop_9 & empty_9 ? 1'h0 : _GEN_2424; // @[stackmanage_35.scala 4937:43 stackmanage_35.scala 4950:34]
  wire  _GEN_2452 = pop_9 & empty_9 ? 1'h0 : _GEN_2425; // @[stackmanage_35.scala 4937:43 stackmanage_35.scala 4951:34]
  wire  _GEN_2453 = pop_9 & empty_9 ? 1'h0 : _GEN_2426; // @[stackmanage_35.scala 4937:43 stackmanage_35.scala 4952:34]
  wire  _GEN_2454 = pop_9 & empty_9 ? 1'h0 : _GEN_2427; // @[stackmanage_35.scala 4937:43 stackmanage_35.scala 4953:34]
  wire  _GEN_2455 = pop_9 & empty_9 ? 1'h0 : _GEN_2428; // @[stackmanage_35.scala 4937:43 stackmanage_35.scala 4954:34]
  wire  _GEN_2456 = pop_9 & empty_9 ? 1'h0 : _GEN_2429; // @[stackmanage_35.scala 4937:43 stackmanage_35.scala 4955:34]
  wire  _GEN_2457 = pop_9 & empty_9 ? 1'h0 : _GEN_2430; // @[stackmanage_35.scala 4937:43 stackmanage_35.scala 4956:34]
  wire  _GEN_2458 = pop_9 & empty_9 ? 1'h0 : _GEN_2431; // @[stackmanage_35.scala 4937:43 stackmanage_35.scala 4957:34]
  wire  _GEN_2459 = pop_9 & empty_9 ? 1'h0 : _GEN_2432; // @[stackmanage_35.scala 4937:43 stackmanage_35.scala 4958:34]
  wire  _GEN_2460 = pop_9 & empty_9 ? 1'h0 : _GEN_2433; // @[stackmanage_35.scala 4937:43 stackmanage_35.scala 4959:34]
  wire  _GEN_2461 = pop_9 & empty_9 ? 1'h0 : _GEN_2434; // @[stackmanage_35.scala 4937:43 stackmanage_35.scala 4960:34]
  wire  _GEN_2462 = pop_9 & empty_9 ? 1'h0 : _GEN_2435; // @[stackmanage_35.scala 4937:43 stackmanage_35.scala 4961:34]
  wire  _GEN_2463 = pop_9 & empty_9 ? 1'h0 : _GEN_2436; // @[stackmanage_35.scala 4937:43 stackmanage_35.scala 4962:34]
  wire  _GEN_2464 = pop_9 & empty_9 ? 1'h0 : _GEN_2437; // @[stackmanage_35.scala 4937:43 stackmanage_35.scala 4963:34]
  wire  _GEN_2465 = pop_9 & empty_9 ? 1'h0 : _GEN_2438; // @[stackmanage_35.scala 4937:43 stackmanage_35.scala 4964:34]
  wire  _GEN_2466 = pop_9 & empty_9 ? 1'h0 : _GEN_2439; // @[stackmanage_35.scala 4937:43 stackmanage_35.scala 4965:34]
  wire  _GEN_2467 = pop_9 & empty_9 ? 1'h0 : _GEN_2440; // @[stackmanage_35.scala 4937:43 stackmanage_35.scala 4966:34]
  wire  _GEN_2468 = pop_9 & empty_9 ? 1'h0 : _GEN_2441; // @[stackmanage_35.scala 4937:43 stackmanage_35.scala 4967:34]
  wire  _GEN_2469 = pop_9 & empty_9 ? 1'h0 : _GEN_2442; // @[stackmanage_35.scala 4937:43 stackmanage_35.scala 4968:34]
  wire  _GEN_2470 = pop_9 & empty_9 ? 1'h0 : _GEN_2443; // @[stackmanage_35.scala 4937:43 stackmanage_35.scala 4969:34]
  wire  _GEN_2471 = pop_9 & empty_9 ? 1'h0 : _GEN_2444; // @[stackmanage_35.scala 4937:43 stackmanage_35.scala 4970:34]
  wire  _GEN_2472 = pop_9 & empty_9 ? 1'h0 : _GEN_2445; // @[stackmanage_35.scala 4937:43 stackmanage_35.scala 4971:34]
  wire  _GEN_2473 = pop_9 & empty_9 ? 1'h0 : _GEN_2446; // @[stackmanage_35.scala 4937:43 stackmanage_35.scala 4972:34]
  wire  _GEN_2474 = pop_9 & empty_9 ? 1'h0 : _GEN_2447; // @[stackmanage_35.scala 4937:43 stackmanage_35.scala 4973:34]
  wire  _GEN_2477 = pop_8 & empty_8 ? 1'h0 : _T_344; // @[stackmanage_35.scala 4900:43 stackmanage_35.scala 4911:33]
  wire  _GEN_2478 = pop_8 & empty_8 ? 1'h0 : _GEN_2450; // @[stackmanage_35.scala 4900:43 stackmanage_35.scala 4912:34]
  wire  _GEN_2479 = pop_8 & empty_8 ? 1'h0 : _GEN_2451; // @[stackmanage_35.scala 4900:43 stackmanage_35.scala 4913:34]
  wire  _GEN_2480 = pop_8 & empty_8 ? 1'h0 : _GEN_2452; // @[stackmanage_35.scala 4900:43 stackmanage_35.scala 4914:34]
  wire  _GEN_2481 = pop_8 & empty_8 ? 1'h0 : _GEN_2453; // @[stackmanage_35.scala 4900:43 stackmanage_35.scala 4915:34]
  wire  _GEN_2482 = pop_8 & empty_8 ? 1'h0 : _GEN_2454; // @[stackmanage_35.scala 4900:43 stackmanage_35.scala 4916:34]
  wire  _GEN_2483 = pop_8 & empty_8 ? 1'h0 : _GEN_2455; // @[stackmanage_35.scala 4900:43 stackmanage_35.scala 4917:34]
  wire  _GEN_2484 = pop_8 & empty_8 ? 1'h0 : _GEN_2456; // @[stackmanage_35.scala 4900:43 stackmanage_35.scala 4918:34]
  wire  _GEN_2485 = pop_8 & empty_8 ? 1'h0 : _GEN_2457; // @[stackmanage_35.scala 4900:43 stackmanage_35.scala 4919:34]
  wire  _GEN_2486 = pop_8 & empty_8 ? 1'h0 : _GEN_2458; // @[stackmanage_35.scala 4900:43 stackmanage_35.scala 4920:34]
  wire  _GEN_2487 = pop_8 & empty_8 ? 1'h0 : _GEN_2459; // @[stackmanage_35.scala 4900:43 stackmanage_35.scala 4921:34]
  wire  _GEN_2488 = pop_8 & empty_8 ? 1'h0 : _GEN_2460; // @[stackmanage_35.scala 4900:43 stackmanage_35.scala 4922:34]
  wire  _GEN_2489 = pop_8 & empty_8 ? 1'h0 : _GEN_2461; // @[stackmanage_35.scala 4900:43 stackmanage_35.scala 4923:34]
  wire  _GEN_2490 = pop_8 & empty_8 ? 1'h0 : _GEN_2462; // @[stackmanage_35.scala 4900:43 stackmanage_35.scala 4924:34]
  wire  _GEN_2491 = pop_8 & empty_8 ? 1'h0 : _GEN_2463; // @[stackmanage_35.scala 4900:43 stackmanage_35.scala 4925:34]
  wire  _GEN_2492 = pop_8 & empty_8 ? 1'h0 : _GEN_2464; // @[stackmanage_35.scala 4900:43 stackmanage_35.scala 4926:34]
  wire  _GEN_2493 = pop_8 & empty_8 ? 1'h0 : _GEN_2465; // @[stackmanage_35.scala 4900:43 stackmanage_35.scala 4927:34]
  wire  _GEN_2494 = pop_8 & empty_8 ? 1'h0 : _GEN_2466; // @[stackmanage_35.scala 4900:43 stackmanage_35.scala 4928:34]
  wire  _GEN_2495 = pop_8 & empty_8 ? 1'h0 : _GEN_2467; // @[stackmanage_35.scala 4900:43 stackmanage_35.scala 4929:34]
  wire  _GEN_2496 = pop_8 & empty_8 ? 1'h0 : _GEN_2468; // @[stackmanage_35.scala 4900:43 stackmanage_35.scala 4930:34]
  wire  _GEN_2497 = pop_8 & empty_8 ? 1'h0 : _GEN_2469; // @[stackmanage_35.scala 4900:43 stackmanage_35.scala 4931:34]
  wire  _GEN_2498 = pop_8 & empty_8 ? 1'h0 : _GEN_2470; // @[stackmanage_35.scala 4900:43 stackmanage_35.scala 4932:34]
  wire  _GEN_2499 = pop_8 & empty_8 ? 1'h0 : _GEN_2471; // @[stackmanage_35.scala 4900:43 stackmanage_35.scala 4933:34]
  wire  _GEN_2500 = pop_8 & empty_8 ? 1'h0 : _GEN_2472; // @[stackmanage_35.scala 4900:43 stackmanage_35.scala 4934:34]
  wire  _GEN_2501 = pop_8 & empty_8 ? 1'h0 : _GEN_2473; // @[stackmanage_35.scala 4900:43 stackmanage_35.scala 4935:34]
  wire  _GEN_2502 = pop_8 & empty_8 ? 1'h0 : _GEN_2474; // @[stackmanage_35.scala 4900:43 stackmanage_35.scala 4936:34]
  wire  _GEN_2505 = pop_7 & empty_7 ? 1'h0 : _T_341; // @[stackmanage_35.scala 4862:43 stackmanage_35.scala 4872:33]
  wire  _GEN_2506 = pop_7 & empty_7 ? 1'h0 : _GEN_2477; // @[stackmanage_35.scala 4862:43 stackmanage_35.scala 4873:33]
  wire  _GEN_2507 = pop_7 & empty_7 ? 1'h0 : _GEN_2478; // @[stackmanage_35.scala 4862:43 stackmanage_35.scala 4874:34]
  wire  _GEN_2508 = pop_7 & empty_7 ? 1'h0 : _GEN_2479; // @[stackmanage_35.scala 4862:43 stackmanage_35.scala 4875:34]
  wire  _GEN_2509 = pop_7 & empty_7 ? 1'h0 : _GEN_2480; // @[stackmanage_35.scala 4862:43 stackmanage_35.scala 4876:34]
  wire  _GEN_2510 = pop_7 & empty_7 ? 1'h0 : _GEN_2481; // @[stackmanage_35.scala 4862:43 stackmanage_35.scala 4877:34]
  wire  _GEN_2511 = pop_7 & empty_7 ? 1'h0 : _GEN_2482; // @[stackmanage_35.scala 4862:43 stackmanage_35.scala 4878:34]
  wire  _GEN_2512 = pop_7 & empty_7 ? 1'h0 : _GEN_2483; // @[stackmanage_35.scala 4862:43 stackmanage_35.scala 4879:34]
  wire  _GEN_2513 = pop_7 & empty_7 ? 1'h0 : _GEN_2484; // @[stackmanage_35.scala 4862:43 stackmanage_35.scala 4880:34]
  wire  _GEN_2514 = pop_7 & empty_7 ? 1'h0 : _GEN_2485; // @[stackmanage_35.scala 4862:43 stackmanage_35.scala 4881:34]
  wire  _GEN_2515 = pop_7 & empty_7 ? 1'h0 : _GEN_2486; // @[stackmanage_35.scala 4862:43 stackmanage_35.scala 4882:34]
  wire  _GEN_2516 = pop_7 & empty_7 ? 1'h0 : _GEN_2487; // @[stackmanage_35.scala 4862:43 stackmanage_35.scala 4883:34]
  wire  _GEN_2517 = pop_7 & empty_7 ? 1'h0 : _GEN_2488; // @[stackmanage_35.scala 4862:43 stackmanage_35.scala 4884:34]
  wire  _GEN_2518 = pop_7 & empty_7 ? 1'h0 : _GEN_2489; // @[stackmanage_35.scala 4862:43 stackmanage_35.scala 4885:34]
  wire  _GEN_2519 = pop_7 & empty_7 ? 1'h0 : _GEN_2490; // @[stackmanage_35.scala 4862:43 stackmanage_35.scala 4886:34]
  wire  _GEN_2520 = pop_7 & empty_7 ? 1'h0 : _GEN_2491; // @[stackmanage_35.scala 4862:43 stackmanage_35.scala 4887:34]
  wire  _GEN_2521 = pop_7 & empty_7 ? 1'h0 : _GEN_2492; // @[stackmanage_35.scala 4862:43 stackmanage_35.scala 4888:34]
  wire  _GEN_2522 = pop_7 & empty_7 ? 1'h0 : _GEN_2493; // @[stackmanage_35.scala 4862:43 stackmanage_35.scala 4889:34]
  wire  _GEN_2523 = pop_7 & empty_7 ? 1'h0 : _GEN_2494; // @[stackmanage_35.scala 4862:43 stackmanage_35.scala 4890:34]
  wire  _GEN_2524 = pop_7 & empty_7 ? 1'h0 : _GEN_2495; // @[stackmanage_35.scala 4862:43 stackmanage_35.scala 4891:34]
  wire  _GEN_2525 = pop_7 & empty_7 ? 1'h0 : _GEN_2496; // @[stackmanage_35.scala 4862:43 stackmanage_35.scala 4892:34]
  wire  _GEN_2526 = pop_7 & empty_7 ? 1'h0 : _GEN_2497; // @[stackmanage_35.scala 4862:43 stackmanage_35.scala 4893:34]
  wire  _GEN_2527 = pop_7 & empty_7 ? 1'h0 : _GEN_2498; // @[stackmanage_35.scala 4862:43 stackmanage_35.scala 4894:34]
  wire  _GEN_2528 = pop_7 & empty_7 ? 1'h0 : _GEN_2499; // @[stackmanage_35.scala 4862:43 stackmanage_35.scala 4895:34]
  wire  _GEN_2529 = pop_7 & empty_7 ? 1'h0 : _GEN_2500; // @[stackmanage_35.scala 4862:43 stackmanage_35.scala 4896:34]
  wire  _GEN_2530 = pop_7 & empty_7 ? 1'h0 : _GEN_2501; // @[stackmanage_35.scala 4862:43 stackmanage_35.scala 4897:34]
  wire  _GEN_2531 = pop_7 & empty_7 ? 1'h0 : _GEN_2502; // @[stackmanage_35.scala 4862:43 stackmanage_35.scala 4898:34]
  wire  _GEN_2534 = pop_6 & empty_6 ? 1'h0 : _T_338; // @[stackmanage_35.scala 4824:43 stackmanage_35.scala 4833:33]
  wire  _GEN_2535 = pop_6 & empty_6 ? 1'h0 : _GEN_2505; // @[stackmanage_35.scala 4824:43 stackmanage_35.scala 4834:33]
  wire  _GEN_2536 = pop_6 & empty_6 ? 1'h0 : _GEN_2506; // @[stackmanage_35.scala 4824:43 stackmanage_35.scala 4835:33]
  wire  _GEN_2537 = pop_6 & empty_6 ? 1'h0 : _GEN_2507; // @[stackmanage_35.scala 4824:43 stackmanage_35.scala 4836:34]
  wire  _GEN_2538 = pop_6 & empty_6 ? 1'h0 : _GEN_2508; // @[stackmanage_35.scala 4824:43 stackmanage_35.scala 4837:34]
  wire  _GEN_2539 = pop_6 & empty_6 ? 1'h0 : _GEN_2509; // @[stackmanage_35.scala 4824:43 stackmanage_35.scala 4838:34]
  wire  _GEN_2540 = pop_6 & empty_6 ? 1'h0 : _GEN_2510; // @[stackmanage_35.scala 4824:43 stackmanage_35.scala 4839:34]
  wire  _GEN_2541 = pop_6 & empty_6 ? 1'h0 : _GEN_2511; // @[stackmanage_35.scala 4824:43 stackmanage_35.scala 4840:34]
  wire  _GEN_2542 = pop_6 & empty_6 ? 1'h0 : _GEN_2512; // @[stackmanage_35.scala 4824:43 stackmanage_35.scala 4841:34]
  wire  _GEN_2543 = pop_6 & empty_6 ? 1'h0 : _GEN_2513; // @[stackmanage_35.scala 4824:43 stackmanage_35.scala 4842:34]
  wire  _GEN_2544 = pop_6 & empty_6 ? 1'h0 : _GEN_2514; // @[stackmanage_35.scala 4824:43 stackmanage_35.scala 4843:34]
  wire  _GEN_2545 = pop_6 & empty_6 ? 1'h0 : _GEN_2515; // @[stackmanage_35.scala 4824:43 stackmanage_35.scala 4844:34]
  wire  _GEN_2546 = pop_6 & empty_6 ? 1'h0 : _GEN_2516; // @[stackmanage_35.scala 4824:43 stackmanage_35.scala 4845:34]
  wire  _GEN_2547 = pop_6 & empty_6 ? 1'h0 : _GEN_2517; // @[stackmanage_35.scala 4824:43 stackmanage_35.scala 4846:34]
  wire  _GEN_2548 = pop_6 & empty_6 ? 1'h0 : _GEN_2518; // @[stackmanage_35.scala 4824:43 stackmanage_35.scala 4847:34]
  wire  _GEN_2549 = pop_6 & empty_6 ? 1'h0 : _GEN_2519; // @[stackmanage_35.scala 4824:43 stackmanage_35.scala 4848:34]
  wire  _GEN_2550 = pop_6 & empty_6 ? 1'h0 : _GEN_2520; // @[stackmanage_35.scala 4824:43 stackmanage_35.scala 4849:34]
  wire  _GEN_2551 = pop_6 & empty_6 ? 1'h0 : _GEN_2521; // @[stackmanage_35.scala 4824:43 stackmanage_35.scala 4850:34]
  wire  _GEN_2552 = pop_6 & empty_6 ? 1'h0 : _GEN_2522; // @[stackmanage_35.scala 4824:43 stackmanage_35.scala 4851:34]
  wire  _GEN_2553 = pop_6 & empty_6 ? 1'h0 : _GEN_2523; // @[stackmanage_35.scala 4824:43 stackmanage_35.scala 4852:34]
  wire  _GEN_2554 = pop_6 & empty_6 ? 1'h0 : _GEN_2524; // @[stackmanage_35.scala 4824:43 stackmanage_35.scala 4853:34]
  wire  _GEN_2555 = pop_6 & empty_6 ? 1'h0 : _GEN_2525; // @[stackmanage_35.scala 4824:43 stackmanage_35.scala 4854:34]
  wire  _GEN_2556 = pop_6 & empty_6 ? 1'h0 : _GEN_2526; // @[stackmanage_35.scala 4824:43 stackmanage_35.scala 4855:34]
  wire  _GEN_2557 = pop_6 & empty_6 ? 1'h0 : _GEN_2527; // @[stackmanage_35.scala 4824:43 stackmanage_35.scala 4856:34]
  wire  _GEN_2558 = pop_6 & empty_6 ? 1'h0 : _GEN_2528; // @[stackmanage_35.scala 4824:43 stackmanage_35.scala 4857:34]
  wire  _GEN_2559 = pop_6 & empty_6 ? 1'h0 : _GEN_2529; // @[stackmanage_35.scala 4824:43 stackmanage_35.scala 4858:34]
  wire  _GEN_2560 = pop_6 & empty_6 ? 1'h0 : _GEN_2530; // @[stackmanage_35.scala 4824:43 stackmanage_35.scala 4859:34]
  wire  _GEN_2561 = pop_6 & empty_6 ? 1'h0 : _GEN_2531; // @[stackmanage_35.scala 4824:43 stackmanage_35.scala 4860:34]
  wire  _GEN_2564 = pop_5 & empty_5 ? 1'h0 : _T_335; // @[stackmanage_35.scala 4786:43 stackmanage_35.scala 4794:33]
  wire  _GEN_2565 = pop_5 & empty_5 ? 1'h0 : _GEN_2534; // @[stackmanage_35.scala 4786:43 stackmanage_35.scala 4795:33]
  wire  _GEN_2566 = pop_5 & empty_5 ? 1'h0 : _GEN_2535; // @[stackmanage_35.scala 4786:43 stackmanage_35.scala 4796:33]
  wire  _GEN_2567 = pop_5 & empty_5 ? 1'h0 : _GEN_2536; // @[stackmanage_35.scala 4786:43 stackmanage_35.scala 4797:33]
  wire  _GEN_2568 = pop_5 & empty_5 ? 1'h0 : _GEN_2537; // @[stackmanage_35.scala 4786:43 stackmanage_35.scala 4798:34]
  wire  _GEN_2569 = pop_5 & empty_5 ? 1'h0 : _GEN_2538; // @[stackmanage_35.scala 4786:43 stackmanage_35.scala 4799:34]
  wire  _GEN_2570 = pop_5 & empty_5 ? 1'h0 : _GEN_2539; // @[stackmanage_35.scala 4786:43 stackmanage_35.scala 4800:34]
  wire  _GEN_2571 = pop_5 & empty_5 ? 1'h0 : _GEN_2540; // @[stackmanage_35.scala 4786:43 stackmanage_35.scala 4801:34]
  wire  _GEN_2572 = pop_5 & empty_5 ? 1'h0 : _GEN_2541; // @[stackmanage_35.scala 4786:43 stackmanage_35.scala 4802:34]
  wire  _GEN_2573 = pop_5 & empty_5 ? 1'h0 : _GEN_2542; // @[stackmanage_35.scala 4786:43 stackmanage_35.scala 4803:34]
  wire  _GEN_2574 = pop_5 & empty_5 ? 1'h0 : _GEN_2543; // @[stackmanage_35.scala 4786:43 stackmanage_35.scala 4804:34]
  wire  _GEN_2575 = pop_5 & empty_5 ? 1'h0 : _GEN_2544; // @[stackmanage_35.scala 4786:43 stackmanage_35.scala 4805:34]
  wire  _GEN_2576 = pop_5 & empty_5 ? 1'h0 : _GEN_2545; // @[stackmanage_35.scala 4786:43 stackmanage_35.scala 4806:34]
  wire  _GEN_2577 = pop_5 & empty_5 ? 1'h0 : _GEN_2546; // @[stackmanage_35.scala 4786:43 stackmanage_35.scala 4807:34]
  wire  _GEN_2578 = pop_5 & empty_5 ? 1'h0 : _GEN_2547; // @[stackmanage_35.scala 4786:43 stackmanage_35.scala 4808:34]
  wire  _GEN_2579 = pop_5 & empty_5 ? 1'h0 : _GEN_2548; // @[stackmanage_35.scala 4786:43 stackmanage_35.scala 4809:34]
  wire  _GEN_2580 = pop_5 & empty_5 ? 1'h0 : _GEN_2549; // @[stackmanage_35.scala 4786:43 stackmanage_35.scala 4810:34]
  wire  _GEN_2581 = pop_5 & empty_5 ? 1'h0 : _GEN_2550; // @[stackmanage_35.scala 4786:43 stackmanage_35.scala 4811:34]
  wire  _GEN_2582 = pop_5 & empty_5 ? 1'h0 : _GEN_2551; // @[stackmanage_35.scala 4786:43 stackmanage_35.scala 4812:34]
  wire  _GEN_2583 = pop_5 & empty_5 ? 1'h0 : _GEN_2552; // @[stackmanage_35.scala 4786:43 stackmanage_35.scala 4813:34]
  wire  _GEN_2584 = pop_5 & empty_5 ? 1'h0 : _GEN_2553; // @[stackmanage_35.scala 4786:43 stackmanage_35.scala 4814:34]
  wire  _GEN_2585 = pop_5 & empty_5 ? 1'h0 : _GEN_2554; // @[stackmanage_35.scala 4786:43 stackmanage_35.scala 4815:34]
  wire  _GEN_2586 = pop_5 & empty_5 ? 1'h0 : _GEN_2555; // @[stackmanage_35.scala 4786:43 stackmanage_35.scala 4816:34]
  wire  _GEN_2587 = pop_5 & empty_5 ? 1'h0 : _GEN_2556; // @[stackmanage_35.scala 4786:43 stackmanage_35.scala 4817:34]
  wire  _GEN_2588 = pop_5 & empty_5 ? 1'h0 : _GEN_2557; // @[stackmanage_35.scala 4786:43 stackmanage_35.scala 4818:34]
  wire  _GEN_2589 = pop_5 & empty_5 ? 1'h0 : _GEN_2558; // @[stackmanage_35.scala 4786:43 stackmanage_35.scala 4819:34]
  wire  _GEN_2590 = pop_5 & empty_5 ? 1'h0 : _GEN_2559; // @[stackmanage_35.scala 4786:43 stackmanage_35.scala 4820:34]
  wire  _GEN_2591 = pop_5 & empty_5 ? 1'h0 : _GEN_2560; // @[stackmanage_35.scala 4786:43 stackmanage_35.scala 4821:34]
  wire  _GEN_2592 = pop_5 & empty_5 ? 1'h0 : _GEN_2561; // @[stackmanage_35.scala 4786:43 stackmanage_35.scala 4822:34]
  wire  _GEN_2595 = pop_4 & empty_4 ? 1'h0 : _T_332; // @[stackmanage_35.scala 4748:43 stackmanage_35.scala 4755:33]
  wire  _GEN_2596 = pop_4 & empty_4 ? 1'h0 : _GEN_2564; // @[stackmanage_35.scala 4748:43 stackmanage_35.scala 4756:33]
  wire  _GEN_2597 = pop_4 & empty_4 ? 1'h0 : _GEN_2565; // @[stackmanage_35.scala 4748:43 stackmanage_35.scala 4757:33]
  wire  _GEN_2598 = pop_4 & empty_4 ? 1'h0 : _GEN_2566; // @[stackmanage_35.scala 4748:43 stackmanage_35.scala 4758:33]
  wire  _GEN_2599 = pop_4 & empty_4 ? 1'h0 : _GEN_2567; // @[stackmanage_35.scala 4748:43 stackmanage_35.scala 4759:33]
  wire  _GEN_2600 = pop_4 & empty_4 ? 1'h0 : _GEN_2568; // @[stackmanage_35.scala 4748:43 stackmanage_35.scala 4760:34]
  wire  _GEN_2601 = pop_4 & empty_4 ? 1'h0 : _GEN_2569; // @[stackmanage_35.scala 4748:43 stackmanage_35.scala 4761:34]
  wire  _GEN_2602 = pop_4 & empty_4 ? 1'h0 : _GEN_2570; // @[stackmanage_35.scala 4748:43 stackmanage_35.scala 4762:34]
  wire  _GEN_2603 = pop_4 & empty_4 ? 1'h0 : _GEN_2571; // @[stackmanage_35.scala 4748:43 stackmanage_35.scala 4763:34]
  wire  _GEN_2604 = pop_4 & empty_4 ? 1'h0 : _GEN_2572; // @[stackmanage_35.scala 4748:43 stackmanage_35.scala 4764:34]
  wire  _GEN_2605 = pop_4 & empty_4 ? 1'h0 : _GEN_2573; // @[stackmanage_35.scala 4748:43 stackmanage_35.scala 4765:34]
  wire  _GEN_2606 = pop_4 & empty_4 ? 1'h0 : _GEN_2574; // @[stackmanage_35.scala 4748:43 stackmanage_35.scala 4766:34]
  wire  _GEN_2607 = pop_4 & empty_4 ? 1'h0 : _GEN_2575; // @[stackmanage_35.scala 4748:43 stackmanage_35.scala 4767:34]
  wire  _GEN_2608 = pop_4 & empty_4 ? 1'h0 : _GEN_2576; // @[stackmanage_35.scala 4748:43 stackmanage_35.scala 4768:34]
  wire  _GEN_2609 = pop_4 & empty_4 ? 1'h0 : _GEN_2577; // @[stackmanage_35.scala 4748:43 stackmanage_35.scala 4769:34]
  wire  _GEN_2610 = pop_4 & empty_4 ? 1'h0 : _GEN_2578; // @[stackmanage_35.scala 4748:43 stackmanage_35.scala 4770:34]
  wire  _GEN_2611 = pop_4 & empty_4 ? 1'h0 : _GEN_2579; // @[stackmanage_35.scala 4748:43 stackmanage_35.scala 4771:34]
  wire  _GEN_2612 = pop_4 & empty_4 ? 1'h0 : _GEN_2580; // @[stackmanage_35.scala 4748:43 stackmanage_35.scala 4772:34]
  wire  _GEN_2613 = pop_4 & empty_4 ? 1'h0 : _GEN_2581; // @[stackmanage_35.scala 4748:43 stackmanage_35.scala 4773:34]
  wire  _GEN_2614 = pop_4 & empty_4 ? 1'h0 : _GEN_2582; // @[stackmanage_35.scala 4748:43 stackmanage_35.scala 4774:34]
  wire  _GEN_2615 = pop_4 & empty_4 ? 1'h0 : _GEN_2583; // @[stackmanage_35.scala 4748:43 stackmanage_35.scala 4775:34]
  wire  _GEN_2616 = pop_4 & empty_4 ? 1'h0 : _GEN_2584; // @[stackmanage_35.scala 4748:43 stackmanage_35.scala 4776:34]
  wire  _GEN_2617 = pop_4 & empty_4 ? 1'h0 : _GEN_2585; // @[stackmanage_35.scala 4748:43 stackmanage_35.scala 4777:34]
  wire  _GEN_2618 = pop_4 & empty_4 ? 1'h0 : _GEN_2586; // @[stackmanage_35.scala 4748:43 stackmanage_35.scala 4778:34]
  wire  _GEN_2619 = pop_4 & empty_4 ? 1'h0 : _GEN_2587; // @[stackmanage_35.scala 4748:43 stackmanage_35.scala 4779:34]
  wire  _GEN_2620 = pop_4 & empty_4 ? 1'h0 : _GEN_2588; // @[stackmanage_35.scala 4748:43 stackmanage_35.scala 4780:34]
  wire  _GEN_2621 = pop_4 & empty_4 ? 1'h0 : _GEN_2589; // @[stackmanage_35.scala 4748:43 stackmanage_35.scala 4781:34]
  wire  _GEN_2622 = pop_4 & empty_4 ? 1'h0 : _GEN_2590; // @[stackmanage_35.scala 4748:43 stackmanage_35.scala 4782:34]
  wire  _GEN_2623 = pop_4 & empty_4 ? 1'h0 : _GEN_2591; // @[stackmanage_35.scala 4748:43 stackmanage_35.scala 4783:34]
  wire  _GEN_2624 = pop_4 & empty_4 ? 1'h0 : _GEN_2592; // @[stackmanage_35.scala 4748:43 stackmanage_35.scala 4784:34]
  wire  _GEN_2627 = pop_3 & empty_3 ? 1'h0 : _T_329; // @[stackmanage_35.scala 4710:43 stackmanage_35.scala 4716:33]
  wire  _GEN_2628 = pop_3 & empty_3 ? 1'h0 : _GEN_2595; // @[stackmanage_35.scala 4710:43 stackmanage_35.scala 4717:33]
  wire  _GEN_2629 = pop_3 & empty_3 ? 1'h0 : _GEN_2596; // @[stackmanage_35.scala 4710:43 stackmanage_35.scala 4718:33]
  wire  _GEN_2630 = pop_3 & empty_3 ? 1'h0 : _GEN_2597; // @[stackmanage_35.scala 4710:43 stackmanage_35.scala 4719:33]
  wire  _GEN_2631 = pop_3 & empty_3 ? 1'h0 : _GEN_2598; // @[stackmanage_35.scala 4710:43 stackmanage_35.scala 4720:33]
  wire  _GEN_2632 = pop_3 & empty_3 ? 1'h0 : _GEN_2599; // @[stackmanage_35.scala 4710:43 stackmanage_35.scala 4721:33]
  wire  _GEN_2633 = pop_3 & empty_3 ? 1'h0 : _GEN_2600; // @[stackmanage_35.scala 4710:43 stackmanage_35.scala 4722:34]
  wire  _GEN_2634 = pop_3 & empty_3 ? 1'h0 : _GEN_2601; // @[stackmanage_35.scala 4710:43 stackmanage_35.scala 4723:34]
  wire  _GEN_2635 = pop_3 & empty_3 ? 1'h0 : _GEN_2602; // @[stackmanage_35.scala 4710:43 stackmanage_35.scala 4724:34]
  wire  _GEN_2636 = pop_3 & empty_3 ? 1'h0 : _GEN_2603; // @[stackmanage_35.scala 4710:43 stackmanage_35.scala 4725:34]
  wire  _GEN_2637 = pop_3 & empty_3 ? 1'h0 : _GEN_2604; // @[stackmanage_35.scala 4710:43 stackmanage_35.scala 4726:34]
  wire  _GEN_2638 = pop_3 & empty_3 ? 1'h0 : _GEN_2605; // @[stackmanage_35.scala 4710:43 stackmanage_35.scala 4727:34]
  wire  _GEN_2639 = pop_3 & empty_3 ? 1'h0 : _GEN_2606; // @[stackmanage_35.scala 4710:43 stackmanage_35.scala 4728:34]
  wire  _GEN_2640 = pop_3 & empty_3 ? 1'h0 : _GEN_2607; // @[stackmanage_35.scala 4710:43 stackmanage_35.scala 4729:34]
  wire  _GEN_2641 = pop_3 & empty_3 ? 1'h0 : _GEN_2608; // @[stackmanage_35.scala 4710:43 stackmanage_35.scala 4730:34]
  wire  _GEN_2642 = pop_3 & empty_3 ? 1'h0 : _GEN_2609; // @[stackmanage_35.scala 4710:43 stackmanage_35.scala 4731:34]
  wire  _GEN_2643 = pop_3 & empty_3 ? 1'h0 : _GEN_2610; // @[stackmanage_35.scala 4710:43 stackmanage_35.scala 4732:34]
  wire  _GEN_2644 = pop_3 & empty_3 ? 1'h0 : _GEN_2611; // @[stackmanage_35.scala 4710:43 stackmanage_35.scala 4733:34]
  wire  _GEN_2645 = pop_3 & empty_3 ? 1'h0 : _GEN_2612; // @[stackmanage_35.scala 4710:43 stackmanage_35.scala 4734:34]
  wire  _GEN_2646 = pop_3 & empty_3 ? 1'h0 : _GEN_2613; // @[stackmanage_35.scala 4710:43 stackmanage_35.scala 4735:34]
  wire  _GEN_2647 = pop_3 & empty_3 ? 1'h0 : _GEN_2614; // @[stackmanage_35.scala 4710:43 stackmanage_35.scala 4736:34]
  wire  _GEN_2648 = pop_3 & empty_3 ? 1'h0 : _GEN_2615; // @[stackmanage_35.scala 4710:43 stackmanage_35.scala 4737:34]
  wire  _GEN_2649 = pop_3 & empty_3 ? 1'h0 : _GEN_2616; // @[stackmanage_35.scala 4710:43 stackmanage_35.scala 4738:34]
  wire  _GEN_2650 = pop_3 & empty_3 ? 1'h0 : _GEN_2617; // @[stackmanage_35.scala 4710:43 stackmanage_35.scala 4739:34]
  wire  _GEN_2651 = pop_3 & empty_3 ? 1'h0 : _GEN_2618; // @[stackmanage_35.scala 4710:43 stackmanage_35.scala 4740:34]
  wire  _GEN_2652 = pop_3 & empty_3 ? 1'h0 : _GEN_2619; // @[stackmanage_35.scala 4710:43 stackmanage_35.scala 4741:34]
  wire  _GEN_2653 = pop_3 & empty_3 ? 1'h0 : _GEN_2620; // @[stackmanage_35.scala 4710:43 stackmanage_35.scala 4742:34]
  wire  _GEN_2654 = pop_3 & empty_3 ? 1'h0 : _GEN_2621; // @[stackmanage_35.scala 4710:43 stackmanage_35.scala 4743:34]
  wire  _GEN_2655 = pop_3 & empty_3 ? 1'h0 : _GEN_2622; // @[stackmanage_35.scala 4710:43 stackmanage_35.scala 4744:34]
  wire  _GEN_2656 = pop_3 & empty_3 ? 1'h0 : _GEN_2623; // @[stackmanage_35.scala 4710:43 stackmanage_35.scala 4745:34]
  wire  _GEN_2657 = pop_3 & empty_3 ? 1'h0 : _GEN_2624; // @[stackmanage_35.scala 4710:43 stackmanage_35.scala 4746:34]
  wire  _T_468 = dispatch_0 | dispatch_1 | dispatch_2 | dispatch_3 | dispatch_4 | dispatch_5 | dispatch_6 | dispatch_7
     | dispatch_8 | dispatch_9 | dispatch_10 | dispatch_11 | dispatch_12 | dispatch_13 | dispatch_14 | dispatch_15 |
    dispatch_16 | dispatch_17 | dispatch_18 | dispatch_19 | dispatch_20 | dispatch_21 | dispatch_22 | dispatch_23 |
    dispatch_24; // @[stackmanage_35.scala 5944:538]
  wire  _T_514 = Stack_0_io_empty & Stack_1_io_empty & Stack_2_io_empty & Stack_3_io_empty & Stack_4_io_empty &
    Stack_5_io_empty & Stack_6_io_empty & Stack_7_io_empty & Stack_8_io_empty & Stack_9_io_empty & Stack_10_io_empty &
    Stack_11_io_empty & Stack_12_io_empty & Stack_13_io_empty & Stack_14_io_empty & Stack_15_io_empty &
    Stack_16_io_empty & Stack_17_io_empty & Stack_18_io_empty & Stack_19_io_empty & Stack_20_io_empty &
    Stack_21_io_empty & Stack_22_io_empty & Stack_23_io_empty & Stack_24_io_empty; // @[stackmanage_35.scala 5946:496]
  LUT LUT_stack ( // @[stackmanage_35.scala 33:45]
    .clock(LUT_stack_clock),
    .reset(LUT_stack_reset),
    .io_push(LUT_stack_io_push),
    .io_push_valid(LUT_stack_io_push_valid),
    .io_pop(LUT_stack_io_pop),
    .io_pop_valid(LUT_stack_io_pop_valid),
    .io_empty_0(LUT_stack_io_empty_0),
    .io_empty_1(LUT_stack_io_empty_1),
    .io_empty_2(LUT_stack_io_empty_2),
    .io_empty_3(LUT_stack_io_empty_3),
    .io_empty_4(LUT_stack_io_empty_4),
    .io_empty_5(LUT_stack_io_empty_5),
    .io_empty_6(LUT_stack_io_empty_6),
    .io_empty_7(LUT_stack_io_empty_7),
    .io_empty_8(LUT_stack_io_empty_8),
    .io_empty_9(LUT_stack_io_empty_9),
    .io_empty_10(LUT_stack_io_empty_10),
    .io_empty_11(LUT_stack_io_empty_11),
    .io_empty_12(LUT_stack_io_empty_12),
    .io_empty_13(LUT_stack_io_empty_13),
    .io_empty_14(LUT_stack_io_empty_14),
    .io_empty_15(LUT_stack_io_empty_15),
    .io_empty_16(LUT_stack_io_empty_16),
    .io_empty_17(LUT_stack_io_empty_17),
    .io_empty_18(LUT_stack_io_empty_18),
    .io_empty_19(LUT_stack_io_empty_19),
    .io_empty_20(LUT_stack_io_empty_20),
    .io_empty_21(LUT_stack_io_empty_21),
    .io_empty_22(LUT_stack_io_empty_22),
    .io_empty_23(LUT_stack_io_empty_23),
    .io_empty_24(LUT_stack_io_empty_24),
    .io_empty_25(LUT_stack_io_empty_25),
    .io_empty_26(LUT_stack_io_empty_26),
    .io_empty_27(LUT_stack_io_empty_27),
    .io_empty_28(LUT_stack_io_empty_28),
    .io_empty_29(LUT_stack_io_empty_29),
    .io_empty_30(LUT_stack_io_empty_30),
    .io_empty_31(LUT_stack_io_empty_31),
    .io_empty_32(LUT_stack_io_empty_32),
    .io_empty_33(LUT_stack_io_empty_33),
    .io_empty_34(LUT_stack_io_empty_34),
    .io_dispatch_0(LUT_stack_io_dispatch_0),
    .io_dispatch_1(LUT_stack_io_dispatch_1),
    .io_dispatch_2(LUT_stack_io_dispatch_2),
    .io_dispatch_3(LUT_stack_io_dispatch_3),
    .io_dispatch_4(LUT_stack_io_dispatch_4),
    .io_dispatch_5(LUT_stack_io_dispatch_5),
    .io_dispatch_6(LUT_stack_io_dispatch_6),
    .io_dispatch_7(LUT_stack_io_dispatch_7),
    .io_dispatch_8(LUT_stack_io_dispatch_8),
    .io_dispatch_9(LUT_stack_io_dispatch_9),
    .io_dispatch_10(LUT_stack_io_dispatch_10),
    .io_dispatch_11(LUT_stack_io_dispatch_11),
    .io_dispatch_12(LUT_stack_io_dispatch_12),
    .io_dispatch_13(LUT_stack_io_dispatch_13),
    .io_dispatch_14(LUT_stack_io_dispatch_14),
    .io_dispatch_15(LUT_stack_io_dispatch_15),
    .io_dispatch_16(LUT_stack_io_dispatch_16),
    .io_dispatch_17(LUT_stack_io_dispatch_17),
    .io_dispatch_18(LUT_stack_io_dispatch_18),
    .io_dispatch_19(LUT_stack_io_dispatch_19),
    .io_dispatch_20(LUT_stack_io_dispatch_20),
    .io_dispatch_21(LUT_stack_io_dispatch_21),
    .io_dispatch_22(LUT_stack_io_dispatch_22),
    .io_dispatch_23(LUT_stack_io_dispatch_23),
    .io_dispatch_24(LUT_stack_io_dispatch_24),
    .io_dispatch_25(LUT_stack_io_dispatch_25),
    .io_dispatch_26(LUT_stack_io_dispatch_26),
    .io_dispatch_27(LUT_stack_io_dispatch_27),
    .io_dispatch_28(LUT_stack_io_dispatch_28),
    .io_dispatch_29(LUT_stack_io_dispatch_29),
    .io_dispatch_30(LUT_stack_io_dispatch_30),
    .io_dispatch_31(LUT_stack_io_dispatch_31),
    .io_dispatch_32(LUT_stack_io_dispatch_32),
    .io_dispatch_33(LUT_stack_io_dispatch_33),
    .io_dispatch_34(LUT_stack_io_dispatch_34),
    .io_ray_id_push(LUT_stack_io_ray_id_push),
    .io_ray_id_pop(LUT_stack_io_ray_id_pop),
    .io_node_id_push_in(LUT_stack_io_node_id_push_in),
    .io_hitT_in(LUT_stack_io_hitT_in),
    .io_ray_id_pop_out(LUT_stack_io_ray_id_pop_out),
    .io_hitT_out(LUT_stack_io_hitT_out),
    .io_pop_0(LUT_stack_io_pop_0),
    .io_pop_1(LUT_stack_io_pop_1),
    .io_pop_2(LUT_stack_io_pop_2),
    .io_pop_3(LUT_stack_io_pop_3),
    .io_pop_4(LUT_stack_io_pop_4),
    .io_pop_5(LUT_stack_io_pop_5),
    .io_pop_6(LUT_stack_io_pop_6),
    .io_pop_7(LUT_stack_io_pop_7),
    .io_pop_8(LUT_stack_io_pop_8),
    .io_pop_9(LUT_stack_io_pop_9),
    .io_pop_10(LUT_stack_io_pop_10),
    .io_pop_11(LUT_stack_io_pop_11),
    .io_pop_12(LUT_stack_io_pop_12),
    .io_pop_13(LUT_stack_io_pop_13),
    .io_pop_14(LUT_stack_io_pop_14),
    .io_pop_15(LUT_stack_io_pop_15),
    .io_pop_16(LUT_stack_io_pop_16),
    .io_pop_17(LUT_stack_io_pop_17),
    .io_pop_18(LUT_stack_io_pop_18),
    .io_pop_19(LUT_stack_io_pop_19),
    .io_pop_20(LUT_stack_io_pop_20),
    .io_pop_21(LUT_stack_io_pop_21),
    .io_pop_22(LUT_stack_io_pop_22),
    .io_pop_23(LUT_stack_io_pop_23),
    .io_pop_24(LUT_stack_io_pop_24),
    .io_pop_25(LUT_stack_io_pop_25),
    .io_pop_26(LUT_stack_io_pop_26),
    .io_pop_27(LUT_stack_io_pop_27),
    .io_pop_28(LUT_stack_io_pop_28),
    .io_pop_29(LUT_stack_io_pop_29),
    .io_pop_30(LUT_stack_io_pop_30),
    .io_pop_31(LUT_stack_io_pop_31),
    .io_pop_32(LUT_stack_io_pop_32),
    .io_pop_33(LUT_stack_io_pop_33),
    .io_pop_34(LUT_stack_io_pop_34),
    .io_pop_en(LUT_stack_io_pop_en),
    .io_push_0(LUT_stack_io_push_0),
    .io_push_1(LUT_stack_io_push_1),
    .io_push_2(LUT_stack_io_push_2),
    .io_push_3(LUT_stack_io_push_3),
    .io_push_4(LUT_stack_io_push_4),
    .io_push_5(LUT_stack_io_push_5),
    .io_push_6(LUT_stack_io_push_6),
    .io_push_7(LUT_stack_io_push_7),
    .io_push_8(LUT_stack_io_push_8),
    .io_push_9(LUT_stack_io_push_9),
    .io_push_10(LUT_stack_io_push_10),
    .io_push_11(LUT_stack_io_push_11),
    .io_push_12(LUT_stack_io_push_12),
    .io_push_13(LUT_stack_io_push_13),
    .io_push_14(LUT_stack_io_push_14),
    .io_push_15(LUT_stack_io_push_15),
    .io_push_16(LUT_stack_io_push_16),
    .io_push_17(LUT_stack_io_push_17),
    .io_push_18(LUT_stack_io_push_18),
    .io_push_19(LUT_stack_io_push_19),
    .io_push_20(LUT_stack_io_push_20),
    .io_push_21(LUT_stack_io_push_21),
    .io_push_22(LUT_stack_io_push_22),
    .io_push_23(LUT_stack_io_push_23),
    .io_push_24(LUT_stack_io_push_24),
    .io_push_25(LUT_stack_io_push_25),
    .io_push_26(LUT_stack_io_push_26),
    .io_push_27(LUT_stack_io_push_27),
    .io_push_28(LUT_stack_io_push_28),
    .io_push_29(LUT_stack_io_push_29),
    .io_push_30(LUT_stack_io_push_30),
    .io_push_31(LUT_stack_io_push_31),
    .io_push_32(LUT_stack_io_push_32),
    .io_push_33(LUT_stack_io_push_33),
    .io_push_34(LUT_stack_io_push_34),
    .io_push_en(LUT_stack_io_push_en),
    .io_no_match(LUT_stack_io_no_match)
  );
  Stack Stack_0 ( // @[stackmanage_35.scala 34:48]
    .clock(Stack_0_clock),
    .reset(Stack_0_reset),
    .io_push(Stack_0_io_push),
    .io_pop(Stack_0_io_pop),
    .io_dataIn(Stack_0_io_dataIn),
    .io_ray_id(Stack_0_io_ray_id),
    .io_dataOut(Stack_0_io_dataOut),
    .io_empty(Stack_0_io_empty),
    .io_hit_in(Stack_0_io_hit_in),
    .io_hit_out(Stack_0_io_hit_out),
    .io_ray_out(Stack_0_io_ray_out),
    .io_enable(Stack_0_io_enable)
  );
  Stack Stack_1 ( // @[stackmanage_35.scala 35:48]
    .clock(Stack_1_clock),
    .reset(Stack_1_reset),
    .io_push(Stack_1_io_push),
    .io_pop(Stack_1_io_pop),
    .io_dataIn(Stack_1_io_dataIn),
    .io_ray_id(Stack_1_io_ray_id),
    .io_dataOut(Stack_1_io_dataOut),
    .io_empty(Stack_1_io_empty),
    .io_hit_in(Stack_1_io_hit_in),
    .io_hit_out(Stack_1_io_hit_out),
    .io_ray_out(Stack_1_io_ray_out),
    .io_enable(Stack_1_io_enable)
  );
  Stack Stack_2 ( // @[stackmanage_35.scala 36:48]
    .clock(Stack_2_clock),
    .reset(Stack_2_reset),
    .io_push(Stack_2_io_push),
    .io_pop(Stack_2_io_pop),
    .io_dataIn(Stack_2_io_dataIn),
    .io_ray_id(Stack_2_io_ray_id),
    .io_dataOut(Stack_2_io_dataOut),
    .io_empty(Stack_2_io_empty),
    .io_hit_in(Stack_2_io_hit_in),
    .io_hit_out(Stack_2_io_hit_out),
    .io_ray_out(Stack_2_io_ray_out),
    .io_enable(Stack_2_io_enable)
  );
  Stack Stack_3 ( // @[stackmanage_35.scala 37:48]
    .clock(Stack_3_clock),
    .reset(Stack_3_reset),
    .io_push(Stack_3_io_push),
    .io_pop(Stack_3_io_pop),
    .io_dataIn(Stack_3_io_dataIn),
    .io_ray_id(Stack_3_io_ray_id),
    .io_dataOut(Stack_3_io_dataOut),
    .io_empty(Stack_3_io_empty),
    .io_hit_in(Stack_3_io_hit_in),
    .io_hit_out(Stack_3_io_hit_out),
    .io_ray_out(Stack_3_io_ray_out),
    .io_enable(Stack_3_io_enable)
  );
  Stack Stack_4 ( // @[stackmanage_35.scala 38:48]
    .clock(Stack_4_clock),
    .reset(Stack_4_reset),
    .io_push(Stack_4_io_push),
    .io_pop(Stack_4_io_pop),
    .io_dataIn(Stack_4_io_dataIn),
    .io_ray_id(Stack_4_io_ray_id),
    .io_dataOut(Stack_4_io_dataOut),
    .io_empty(Stack_4_io_empty),
    .io_hit_in(Stack_4_io_hit_in),
    .io_hit_out(Stack_4_io_hit_out),
    .io_ray_out(Stack_4_io_ray_out),
    .io_enable(Stack_4_io_enable)
  );
  Stack Stack_5 ( // @[stackmanage_35.scala 39:48]
    .clock(Stack_5_clock),
    .reset(Stack_5_reset),
    .io_push(Stack_5_io_push),
    .io_pop(Stack_5_io_pop),
    .io_dataIn(Stack_5_io_dataIn),
    .io_ray_id(Stack_5_io_ray_id),
    .io_dataOut(Stack_5_io_dataOut),
    .io_empty(Stack_5_io_empty),
    .io_hit_in(Stack_5_io_hit_in),
    .io_hit_out(Stack_5_io_hit_out),
    .io_ray_out(Stack_5_io_ray_out),
    .io_enable(Stack_5_io_enable)
  );
  Stack Stack_6 ( // @[stackmanage_35.scala 40:48]
    .clock(Stack_6_clock),
    .reset(Stack_6_reset),
    .io_push(Stack_6_io_push),
    .io_pop(Stack_6_io_pop),
    .io_dataIn(Stack_6_io_dataIn),
    .io_ray_id(Stack_6_io_ray_id),
    .io_dataOut(Stack_6_io_dataOut),
    .io_empty(Stack_6_io_empty),
    .io_hit_in(Stack_6_io_hit_in),
    .io_hit_out(Stack_6_io_hit_out),
    .io_ray_out(Stack_6_io_ray_out),
    .io_enable(Stack_6_io_enable)
  );
  Stack Stack_7 ( // @[stackmanage_35.scala 41:48]
    .clock(Stack_7_clock),
    .reset(Stack_7_reset),
    .io_push(Stack_7_io_push),
    .io_pop(Stack_7_io_pop),
    .io_dataIn(Stack_7_io_dataIn),
    .io_ray_id(Stack_7_io_ray_id),
    .io_dataOut(Stack_7_io_dataOut),
    .io_empty(Stack_7_io_empty),
    .io_hit_in(Stack_7_io_hit_in),
    .io_hit_out(Stack_7_io_hit_out),
    .io_ray_out(Stack_7_io_ray_out),
    .io_enable(Stack_7_io_enable)
  );
  Stack Stack_8 ( // @[stackmanage_35.scala 42:48]
    .clock(Stack_8_clock),
    .reset(Stack_8_reset),
    .io_push(Stack_8_io_push),
    .io_pop(Stack_8_io_pop),
    .io_dataIn(Stack_8_io_dataIn),
    .io_ray_id(Stack_8_io_ray_id),
    .io_dataOut(Stack_8_io_dataOut),
    .io_empty(Stack_8_io_empty),
    .io_hit_in(Stack_8_io_hit_in),
    .io_hit_out(Stack_8_io_hit_out),
    .io_ray_out(Stack_8_io_ray_out),
    .io_enable(Stack_8_io_enable)
  );
  Stack Stack_9 ( // @[stackmanage_35.scala 43:48]
    .clock(Stack_9_clock),
    .reset(Stack_9_reset),
    .io_push(Stack_9_io_push),
    .io_pop(Stack_9_io_pop),
    .io_dataIn(Stack_9_io_dataIn),
    .io_ray_id(Stack_9_io_ray_id),
    .io_dataOut(Stack_9_io_dataOut),
    .io_empty(Stack_9_io_empty),
    .io_hit_in(Stack_9_io_hit_in),
    .io_hit_out(Stack_9_io_hit_out),
    .io_ray_out(Stack_9_io_ray_out),
    .io_enable(Stack_9_io_enable)
  );
  Stack Stack_10 ( // @[stackmanage_35.scala 44:47]
    .clock(Stack_10_clock),
    .reset(Stack_10_reset),
    .io_push(Stack_10_io_push),
    .io_pop(Stack_10_io_pop),
    .io_dataIn(Stack_10_io_dataIn),
    .io_ray_id(Stack_10_io_ray_id),
    .io_dataOut(Stack_10_io_dataOut),
    .io_empty(Stack_10_io_empty),
    .io_hit_in(Stack_10_io_hit_in),
    .io_hit_out(Stack_10_io_hit_out),
    .io_ray_out(Stack_10_io_ray_out),
    .io_enable(Stack_10_io_enable)
  );
  Stack Stack_11 ( // @[stackmanage_35.scala 45:47]
    .clock(Stack_11_clock),
    .reset(Stack_11_reset),
    .io_push(Stack_11_io_push),
    .io_pop(Stack_11_io_pop),
    .io_dataIn(Stack_11_io_dataIn),
    .io_ray_id(Stack_11_io_ray_id),
    .io_dataOut(Stack_11_io_dataOut),
    .io_empty(Stack_11_io_empty),
    .io_hit_in(Stack_11_io_hit_in),
    .io_hit_out(Stack_11_io_hit_out),
    .io_ray_out(Stack_11_io_ray_out),
    .io_enable(Stack_11_io_enable)
  );
  Stack Stack_12 ( // @[stackmanage_35.scala 46:47]
    .clock(Stack_12_clock),
    .reset(Stack_12_reset),
    .io_push(Stack_12_io_push),
    .io_pop(Stack_12_io_pop),
    .io_dataIn(Stack_12_io_dataIn),
    .io_ray_id(Stack_12_io_ray_id),
    .io_dataOut(Stack_12_io_dataOut),
    .io_empty(Stack_12_io_empty),
    .io_hit_in(Stack_12_io_hit_in),
    .io_hit_out(Stack_12_io_hit_out),
    .io_ray_out(Stack_12_io_ray_out),
    .io_enable(Stack_12_io_enable)
  );
  Stack Stack_13 ( // @[stackmanage_35.scala 47:47]
    .clock(Stack_13_clock),
    .reset(Stack_13_reset),
    .io_push(Stack_13_io_push),
    .io_pop(Stack_13_io_pop),
    .io_dataIn(Stack_13_io_dataIn),
    .io_ray_id(Stack_13_io_ray_id),
    .io_dataOut(Stack_13_io_dataOut),
    .io_empty(Stack_13_io_empty),
    .io_hit_in(Stack_13_io_hit_in),
    .io_hit_out(Stack_13_io_hit_out),
    .io_ray_out(Stack_13_io_ray_out),
    .io_enable(Stack_13_io_enable)
  );
  Stack Stack_14 ( // @[stackmanage_35.scala 48:47]
    .clock(Stack_14_clock),
    .reset(Stack_14_reset),
    .io_push(Stack_14_io_push),
    .io_pop(Stack_14_io_pop),
    .io_dataIn(Stack_14_io_dataIn),
    .io_ray_id(Stack_14_io_ray_id),
    .io_dataOut(Stack_14_io_dataOut),
    .io_empty(Stack_14_io_empty),
    .io_hit_in(Stack_14_io_hit_in),
    .io_hit_out(Stack_14_io_hit_out),
    .io_ray_out(Stack_14_io_ray_out),
    .io_enable(Stack_14_io_enable)
  );
  Stack Stack_15 ( // @[stackmanage_35.scala 49:47]
    .clock(Stack_15_clock),
    .reset(Stack_15_reset),
    .io_push(Stack_15_io_push),
    .io_pop(Stack_15_io_pop),
    .io_dataIn(Stack_15_io_dataIn),
    .io_ray_id(Stack_15_io_ray_id),
    .io_dataOut(Stack_15_io_dataOut),
    .io_empty(Stack_15_io_empty),
    .io_hit_in(Stack_15_io_hit_in),
    .io_hit_out(Stack_15_io_hit_out),
    .io_ray_out(Stack_15_io_ray_out),
    .io_enable(Stack_15_io_enable)
  );
  Stack Stack_16 ( // @[stackmanage_35.scala 50:49]
    .clock(Stack_16_clock),
    .reset(Stack_16_reset),
    .io_push(Stack_16_io_push),
    .io_pop(Stack_16_io_pop),
    .io_dataIn(Stack_16_io_dataIn),
    .io_ray_id(Stack_16_io_ray_id),
    .io_dataOut(Stack_16_io_dataOut),
    .io_empty(Stack_16_io_empty),
    .io_hit_in(Stack_16_io_hit_in),
    .io_hit_out(Stack_16_io_hit_out),
    .io_ray_out(Stack_16_io_ray_out),
    .io_enable(Stack_16_io_enable)
  );
  Stack Stack_17 ( // @[stackmanage_35.scala 51:49]
    .clock(Stack_17_clock),
    .reset(Stack_17_reset),
    .io_push(Stack_17_io_push),
    .io_pop(Stack_17_io_pop),
    .io_dataIn(Stack_17_io_dataIn),
    .io_ray_id(Stack_17_io_ray_id),
    .io_dataOut(Stack_17_io_dataOut),
    .io_empty(Stack_17_io_empty),
    .io_hit_in(Stack_17_io_hit_in),
    .io_hit_out(Stack_17_io_hit_out),
    .io_ray_out(Stack_17_io_ray_out),
    .io_enable(Stack_17_io_enable)
  );
  Stack Stack_18 ( // @[stackmanage_35.scala 52:49]
    .clock(Stack_18_clock),
    .reset(Stack_18_reset),
    .io_push(Stack_18_io_push),
    .io_pop(Stack_18_io_pop),
    .io_dataIn(Stack_18_io_dataIn),
    .io_ray_id(Stack_18_io_ray_id),
    .io_dataOut(Stack_18_io_dataOut),
    .io_empty(Stack_18_io_empty),
    .io_hit_in(Stack_18_io_hit_in),
    .io_hit_out(Stack_18_io_hit_out),
    .io_ray_out(Stack_18_io_ray_out),
    .io_enable(Stack_18_io_enable)
  );
  Stack Stack_19 ( // @[stackmanage_35.scala 53:49]
    .clock(Stack_19_clock),
    .reset(Stack_19_reset),
    .io_push(Stack_19_io_push),
    .io_pop(Stack_19_io_pop),
    .io_dataIn(Stack_19_io_dataIn),
    .io_ray_id(Stack_19_io_ray_id),
    .io_dataOut(Stack_19_io_dataOut),
    .io_empty(Stack_19_io_empty),
    .io_hit_in(Stack_19_io_hit_in),
    .io_hit_out(Stack_19_io_hit_out),
    .io_ray_out(Stack_19_io_ray_out),
    .io_enable(Stack_19_io_enable)
  );
  Stack Stack_20 ( // @[stackmanage_35.scala 54:49]
    .clock(Stack_20_clock),
    .reset(Stack_20_reset),
    .io_push(Stack_20_io_push),
    .io_pop(Stack_20_io_pop),
    .io_dataIn(Stack_20_io_dataIn),
    .io_ray_id(Stack_20_io_ray_id),
    .io_dataOut(Stack_20_io_dataOut),
    .io_empty(Stack_20_io_empty),
    .io_hit_in(Stack_20_io_hit_in),
    .io_hit_out(Stack_20_io_hit_out),
    .io_ray_out(Stack_20_io_ray_out),
    .io_enable(Stack_20_io_enable)
  );
  Stack Stack_21 ( // @[stackmanage_35.scala 55:49]
    .clock(Stack_21_clock),
    .reset(Stack_21_reset),
    .io_push(Stack_21_io_push),
    .io_pop(Stack_21_io_pop),
    .io_dataIn(Stack_21_io_dataIn),
    .io_ray_id(Stack_21_io_ray_id),
    .io_dataOut(Stack_21_io_dataOut),
    .io_empty(Stack_21_io_empty),
    .io_hit_in(Stack_21_io_hit_in),
    .io_hit_out(Stack_21_io_hit_out),
    .io_ray_out(Stack_21_io_ray_out),
    .io_enable(Stack_21_io_enable)
  );
  Stack Stack_22 ( // @[stackmanage_35.scala 56:49]
    .clock(Stack_22_clock),
    .reset(Stack_22_reset),
    .io_push(Stack_22_io_push),
    .io_pop(Stack_22_io_pop),
    .io_dataIn(Stack_22_io_dataIn),
    .io_ray_id(Stack_22_io_ray_id),
    .io_dataOut(Stack_22_io_dataOut),
    .io_empty(Stack_22_io_empty),
    .io_hit_in(Stack_22_io_hit_in),
    .io_hit_out(Stack_22_io_hit_out),
    .io_ray_out(Stack_22_io_ray_out),
    .io_enable(Stack_22_io_enable)
  );
  Stack Stack_23 ( // @[stackmanage_35.scala 57:48]
    .clock(Stack_23_clock),
    .reset(Stack_23_reset),
    .io_push(Stack_23_io_push),
    .io_pop(Stack_23_io_pop),
    .io_dataIn(Stack_23_io_dataIn),
    .io_ray_id(Stack_23_io_ray_id),
    .io_dataOut(Stack_23_io_dataOut),
    .io_empty(Stack_23_io_empty),
    .io_hit_in(Stack_23_io_hit_in),
    .io_hit_out(Stack_23_io_hit_out),
    .io_ray_out(Stack_23_io_ray_out),
    .io_enable(Stack_23_io_enable)
  );
  Stack Stack_24 ( // @[stackmanage_35.scala 58:48]
    .clock(Stack_24_clock),
    .reset(Stack_24_reset),
    .io_push(Stack_24_io_push),
    .io_pop(Stack_24_io_pop),
    .io_dataIn(Stack_24_io_dataIn),
    .io_ray_id(Stack_24_io_ray_id),
    .io_dataOut(Stack_24_io_dataOut),
    .io_empty(Stack_24_io_empty),
    .io_hit_in(Stack_24_io_hit_in),
    .io_hit_out(Stack_24_io_hit_out),
    .io_ray_out(Stack_24_io_ray_out),
    .io_enable(Stack_24_io_enable)
  );
  Stack Stack_25 ( // @[stackmanage_35.scala 59:49]
    .clock(Stack_25_clock),
    .reset(Stack_25_reset),
    .io_push(Stack_25_io_push),
    .io_pop(Stack_25_io_pop),
    .io_dataIn(Stack_25_io_dataIn),
    .io_ray_id(Stack_25_io_ray_id),
    .io_dataOut(Stack_25_io_dataOut),
    .io_empty(Stack_25_io_empty),
    .io_hit_in(Stack_25_io_hit_in),
    .io_hit_out(Stack_25_io_hit_out),
    .io_ray_out(Stack_25_io_ray_out),
    .io_enable(Stack_25_io_enable)
  );
  Stack Stack_26 ( // @[stackmanage_35.scala 60:47]
    .clock(Stack_26_clock),
    .reset(Stack_26_reset),
    .io_push(Stack_26_io_push),
    .io_pop(Stack_26_io_pop),
    .io_dataIn(Stack_26_io_dataIn),
    .io_ray_id(Stack_26_io_ray_id),
    .io_dataOut(Stack_26_io_dataOut),
    .io_empty(Stack_26_io_empty),
    .io_hit_in(Stack_26_io_hit_in),
    .io_hit_out(Stack_26_io_hit_out),
    .io_ray_out(Stack_26_io_ray_out),
    .io_enable(Stack_26_io_enable)
  );
  Stack Stack_27 ( // @[stackmanage_35.scala 61:47]
    .clock(Stack_27_clock),
    .reset(Stack_27_reset),
    .io_push(Stack_27_io_push),
    .io_pop(Stack_27_io_pop),
    .io_dataIn(Stack_27_io_dataIn),
    .io_ray_id(Stack_27_io_ray_id),
    .io_dataOut(Stack_27_io_dataOut),
    .io_empty(Stack_27_io_empty),
    .io_hit_in(Stack_27_io_hit_in),
    .io_hit_out(Stack_27_io_hit_out),
    .io_ray_out(Stack_27_io_ray_out),
    .io_enable(Stack_27_io_enable)
  );
  Stack Stack_28 ( // @[stackmanage_35.scala 62:47]
    .clock(Stack_28_clock),
    .reset(Stack_28_reset),
    .io_push(Stack_28_io_push),
    .io_pop(Stack_28_io_pop),
    .io_dataIn(Stack_28_io_dataIn),
    .io_ray_id(Stack_28_io_ray_id),
    .io_dataOut(Stack_28_io_dataOut),
    .io_empty(Stack_28_io_empty),
    .io_hit_in(Stack_28_io_hit_in),
    .io_hit_out(Stack_28_io_hit_out),
    .io_ray_out(Stack_28_io_ray_out),
    .io_enable(Stack_28_io_enable)
  );
  Stack Stack_29 ( // @[stackmanage_35.scala 63:47]
    .clock(Stack_29_clock),
    .reset(Stack_29_reset),
    .io_push(Stack_29_io_push),
    .io_pop(Stack_29_io_pop),
    .io_dataIn(Stack_29_io_dataIn),
    .io_ray_id(Stack_29_io_ray_id),
    .io_dataOut(Stack_29_io_dataOut),
    .io_empty(Stack_29_io_empty),
    .io_hit_in(Stack_29_io_hit_in),
    .io_hit_out(Stack_29_io_hit_out),
    .io_ray_out(Stack_29_io_ray_out),
    .io_enable(Stack_29_io_enable)
  );
  Stack Stack_30 ( // @[stackmanage_35.scala 64:47]
    .clock(Stack_30_clock),
    .reset(Stack_30_reset),
    .io_push(Stack_30_io_push),
    .io_pop(Stack_30_io_pop),
    .io_dataIn(Stack_30_io_dataIn),
    .io_ray_id(Stack_30_io_ray_id),
    .io_dataOut(Stack_30_io_dataOut),
    .io_empty(Stack_30_io_empty),
    .io_hit_in(Stack_30_io_hit_in),
    .io_hit_out(Stack_30_io_hit_out),
    .io_ray_out(Stack_30_io_ray_out),
    .io_enable(Stack_30_io_enable)
  );
  Stack Stack_31 ( // @[stackmanage_35.scala 65:47]
    .clock(Stack_31_clock),
    .reset(Stack_31_reset),
    .io_push(Stack_31_io_push),
    .io_pop(Stack_31_io_pop),
    .io_dataIn(Stack_31_io_dataIn),
    .io_ray_id(Stack_31_io_ray_id),
    .io_dataOut(Stack_31_io_dataOut),
    .io_empty(Stack_31_io_empty),
    .io_hit_in(Stack_31_io_hit_in),
    .io_hit_out(Stack_31_io_hit_out),
    .io_ray_out(Stack_31_io_ray_out),
    .io_enable(Stack_31_io_enable)
  );
  Stack Stack_32 ( // @[stackmanage_35.scala 66:49]
    .clock(Stack_32_clock),
    .reset(Stack_32_reset),
    .io_push(Stack_32_io_push),
    .io_pop(Stack_32_io_pop),
    .io_dataIn(Stack_32_io_dataIn),
    .io_ray_id(Stack_32_io_ray_id),
    .io_dataOut(Stack_32_io_dataOut),
    .io_empty(Stack_32_io_empty),
    .io_hit_in(Stack_32_io_hit_in),
    .io_hit_out(Stack_32_io_hit_out),
    .io_ray_out(Stack_32_io_ray_out),
    .io_enable(Stack_32_io_enable)
  );
  Stack Stack_33 ( // @[stackmanage_35.scala 67:48]
    .clock(Stack_33_clock),
    .reset(Stack_33_reset),
    .io_push(Stack_33_io_push),
    .io_pop(Stack_33_io_pop),
    .io_dataIn(Stack_33_io_dataIn),
    .io_ray_id(Stack_33_io_ray_id),
    .io_dataOut(Stack_33_io_dataOut),
    .io_empty(Stack_33_io_empty),
    .io_hit_in(Stack_33_io_hit_in),
    .io_hit_out(Stack_33_io_hit_out),
    .io_ray_out(Stack_33_io_ray_out),
    .io_enable(Stack_33_io_enable)
  );
  Stack Stack_34 ( // @[stackmanage_35.scala 68:48]
    .clock(Stack_34_clock),
    .reset(Stack_34_reset),
    .io_push(Stack_34_io_push),
    .io_pop(Stack_34_io_pop),
    .io_dataIn(Stack_34_io_dataIn),
    .io_ray_id(Stack_34_io_ray_id),
    .io_dataOut(Stack_34_io_dataOut),
    .io_empty(Stack_34_io_empty),
    .io_hit_in(Stack_34_io_hit_in),
    .io_hit_out(Stack_34_io_hit_out),
    .io_ray_out(Stack_34_io_ray_out),
    .io_enable(Stack_34_io_enable)
  );
  assign io_hitT_out = hitT_out_temp; // @[stackmanage_35.scala 4471:33]
  assign io_node_id_out = node_out_temp; // @[stackmanage_35.scala 4472:27]
  assign io_ray_id_out = ray_out_temp; // @[stackmanage_35.scala 4473:30]
  assign io_pop_valid = pop_valid_1; // @[stackmanage_35.scala 4474:31]
  assign io_Dis_en = _T_468 | dispatch_25 | dispatch_26 | dispatch_27 | dispatch_28 | dispatch_29 | dispatch_30 |
    dispatch_31 | dispatch_32 | dispatch_33 | dispatch_34 | dispatch_no_match; // @[stackmanage_35.scala 5945:275]
  assign io_Finish = _T_514 & Stack_25_io_empty & Stack_26_io_empty & Stack_27_io_empty & Stack_28_io_empty &
    Stack_29_io_empty & Stack_30_io_empty & Stack_31_io_empty & Stack_32_io_empty & Stack_33_io_empty &
    Stack_34_io_empty; // @[stackmanage_35.scala 5947:237]
  assign LUT_stack_clock = clock;
  assign LUT_stack_reset = reset;
  assign LUT_stack_io_push = io_push; // @[stackmanage_35.scala 191:42]
  assign LUT_stack_io_push_valid = io_push_en; // @[stackmanage_35.scala 192:35]
  assign LUT_stack_io_pop = io_pop; // @[stackmanage_35.scala 193:42]
  assign LUT_stack_io_pop_valid = io_pop_en; // @[stackmanage_35.scala 194:36]
  assign LUT_stack_io_empty_0 = Stack_0_io_empty; // @[stackmanage_35.scala 70:29]
  assign LUT_stack_io_empty_1 = Stack_1_io_empty; // @[stackmanage_35.scala 71:29]
  assign LUT_stack_io_empty_2 = Stack_2_io_empty; // @[stackmanage_35.scala 72:29]
  assign LUT_stack_io_empty_3 = Stack_3_io_empty; // @[stackmanage_35.scala 73:29]
  assign LUT_stack_io_empty_4 = Stack_4_io_empty; // @[stackmanage_35.scala 74:29]
  assign LUT_stack_io_empty_5 = Stack_5_io_empty; // @[stackmanage_35.scala 75:29]
  assign LUT_stack_io_empty_6 = Stack_6_io_empty; // @[stackmanage_35.scala 76:29]
  assign LUT_stack_io_empty_7 = Stack_7_io_empty; // @[stackmanage_35.scala 77:29]
  assign LUT_stack_io_empty_8 = Stack_8_io_empty; // @[stackmanage_35.scala 78:29]
  assign LUT_stack_io_empty_9 = Stack_9_io_empty; // @[stackmanage_35.scala 79:29]
  assign LUT_stack_io_empty_10 = Stack_10_io_empty; // @[stackmanage_35.scala 81:30]
  assign LUT_stack_io_empty_11 = Stack_11_io_empty; // @[stackmanage_35.scala 82:30]
  assign LUT_stack_io_empty_12 = Stack_12_io_empty; // @[stackmanage_35.scala 83:30]
  assign LUT_stack_io_empty_13 = Stack_13_io_empty; // @[stackmanage_35.scala 84:30]
  assign LUT_stack_io_empty_14 = Stack_14_io_empty; // @[stackmanage_35.scala 85:30]
  assign LUT_stack_io_empty_15 = Stack_15_io_empty; // @[stackmanage_35.scala 86:30]
  assign LUT_stack_io_empty_16 = Stack_16_io_empty; // @[stackmanage_35.scala 87:30]
  assign LUT_stack_io_empty_17 = Stack_17_io_empty; // @[stackmanage_35.scala 88:30]
  assign LUT_stack_io_empty_18 = Stack_18_io_empty; // @[stackmanage_35.scala 89:30]
  assign LUT_stack_io_empty_19 = Stack_19_io_empty; // @[stackmanage_35.scala 90:30]
  assign LUT_stack_io_empty_20 = Stack_20_io_empty; // @[stackmanage_35.scala 92:30]
  assign LUT_stack_io_empty_21 = Stack_21_io_empty; // @[stackmanage_35.scala 93:30]
  assign LUT_stack_io_empty_22 = Stack_22_io_empty; // @[stackmanage_35.scala 94:30]
  assign LUT_stack_io_empty_23 = Stack_23_io_empty; // @[stackmanage_35.scala 95:30]
  assign LUT_stack_io_empty_24 = Stack_24_io_empty; // @[stackmanage_35.scala 96:30]
  assign LUT_stack_io_empty_25 = Stack_25_io_empty; // @[stackmanage_35.scala 97:30]
  assign LUT_stack_io_empty_26 = Stack_26_io_empty; // @[stackmanage_35.scala 98:30]
  assign LUT_stack_io_empty_27 = Stack_27_io_empty; // @[stackmanage_35.scala 99:30]
  assign LUT_stack_io_empty_28 = Stack_28_io_empty; // @[stackmanage_35.scala 100:30]
  assign LUT_stack_io_empty_29 = Stack_29_io_empty; // @[stackmanage_35.scala 101:30]
  assign LUT_stack_io_empty_30 = Stack_30_io_empty; // @[stackmanage_35.scala 103:30]
  assign LUT_stack_io_empty_31 = Stack_31_io_empty; // @[stackmanage_35.scala 104:30]
  assign LUT_stack_io_empty_32 = Stack_32_io_empty; // @[stackmanage_35.scala 105:30]
  assign LUT_stack_io_empty_33 = Stack_33_io_empty; // @[stackmanage_35.scala 106:30]
  assign LUT_stack_io_empty_34 = Stack_34_io_empty; // @[stackmanage_35.scala 107:30]
  assign LUT_stack_io_dispatch_0 = dispatch_0; // @[stackmanage_35.scala 5951:39]
  assign LUT_stack_io_dispatch_1 = dispatch_1; // @[stackmanage_35.scala 5952:39]
  assign LUT_stack_io_dispatch_2 = dispatch_2; // @[stackmanage_35.scala 5953:39]
  assign LUT_stack_io_dispatch_3 = dispatch_3; // @[stackmanage_35.scala 5954:39]
  assign LUT_stack_io_dispatch_4 = dispatch_4; // @[stackmanage_35.scala 5955:39]
  assign LUT_stack_io_dispatch_5 = dispatch_5; // @[stackmanage_35.scala 5956:39]
  assign LUT_stack_io_dispatch_6 = dispatch_6; // @[stackmanage_35.scala 5957:39]
  assign LUT_stack_io_dispatch_7 = dispatch_7; // @[stackmanage_35.scala 5958:39]
  assign LUT_stack_io_dispatch_8 = dispatch_8; // @[stackmanage_35.scala 5959:39]
  assign LUT_stack_io_dispatch_9 = dispatch_9; // @[stackmanage_35.scala 5960:39]
  assign LUT_stack_io_dispatch_10 = dispatch_10; // @[stackmanage_35.scala 5961:40]
  assign LUT_stack_io_dispatch_11 = dispatch_11; // @[stackmanage_35.scala 5962:40]
  assign LUT_stack_io_dispatch_12 = dispatch_12; // @[stackmanage_35.scala 5963:40]
  assign LUT_stack_io_dispatch_13 = dispatch_13; // @[stackmanage_35.scala 5964:40]
  assign LUT_stack_io_dispatch_14 = dispatch_14; // @[stackmanage_35.scala 5965:40]
  assign LUT_stack_io_dispatch_15 = dispatch_15; // @[stackmanage_35.scala 5966:40]
  assign LUT_stack_io_dispatch_16 = dispatch_16; // @[stackmanage_35.scala 5967:40]
  assign LUT_stack_io_dispatch_17 = dispatch_17; // @[stackmanage_35.scala 5968:40]
  assign LUT_stack_io_dispatch_18 = dispatch_18; // @[stackmanage_35.scala 5969:40]
  assign LUT_stack_io_dispatch_19 = dispatch_19; // @[stackmanage_35.scala 5970:40]
  assign LUT_stack_io_dispatch_20 = dispatch_20; // @[stackmanage_35.scala 5971:40]
  assign LUT_stack_io_dispatch_21 = dispatch_21; // @[stackmanage_35.scala 5972:40]
  assign LUT_stack_io_dispatch_22 = dispatch_22; // @[stackmanage_35.scala 5973:40]
  assign LUT_stack_io_dispatch_23 = dispatch_23; // @[stackmanage_35.scala 5974:40]
  assign LUT_stack_io_dispatch_24 = dispatch_24; // @[stackmanage_35.scala 5975:40]
  assign LUT_stack_io_dispatch_25 = dispatch_25; // @[stackmanage_35.scala 5976:40]
  assign LUT_stack_io_dispatch_26 = dispatch_26; // @[stackmanage_35.scala 5977:40]
  assign LUT_stack_io_dispatch_27 = dispatch_27; // @[stackmanage_35.scala 5978:40]
  assign LUT_stack_io_dispatch_28 = dispatch_28; // @[stackmanage_35.scala 5979:40]
  assign LUT_stack_io_dispatch_29 = dispatch_29; // @[stackmanage_35.scala 5980:40]
  assign LUT_stack_io_dispatch_30 = dispatch_30; // @[stackmanage_35.scala 5981:40]
  assign LUT_stack_io_dispatch_31 = dispatch_31; // @[stackmanage_35.scala 5982:40]
  assign LUT_stack_io_dispatch_32 = dispatch_32; // @[stackmanage_35.scala 5983:40]
  assign LUT_stack_io_dispatch_33 = dispatch_33; // @[stackmanage_35.scala 5984:40]
  assign LUT_stack_io_dispatch_34 = dispatch_34; // @[stackmanage_35.scala 5985:40]
  assign LUT_stack_io_ray_id_push = io_ray_id_push; // @[stackmanage_35.scala 195:33]
  assign LUT_stack_io_ray_id_pop = io_ray_id_pop; // @[stackmanage_35.scala 196:34]
  assign LUT_stack_io_node_id_push_in = io_node_id_push_in; // @[stackmanage_35.scala 197:37]
  assign LUT_stack_io_hitT_in = io_hitT_in; // @[stackmanage_35.scala 199:51]
  assign Stack_0_clock = clock;
  assign Stack_0_reset = reset;
  assign Stack_0_io_push = LUT_stack_io_push_0; // @[stackmanage_35.scala 149:37]
  assign Stack_0_io_pop = LUT_stack_io_pop_0; // @[stackmanage_35.scala 110:38]
  assign Stack_0_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(node_push_in_2) : $signed(32'sh0); // @[stackmanage_35.scala 339:64 stackmanage_35.scala 340:28]
  assign Stack_0_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? LUT_stack_io_ray_id_pop_out : 32'h0; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1644:28]
  assign Stack_0_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? LUT_stack_io_hitT_out : 32'h0; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1643:28]
  assign Stack_1_clock = clock;
  assign Stack_1_reset = reset;
  assign Stack_1_io_push = LUT_stack_io_push_1; // @[stackmanage_35.scala 150:37]
  assign Stack_1_io_pop = LUT_stack_io_pop_1; // @[stackmanage_35.scala 111:38]
  assign Stack_1_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_594); // @[stackmanage_35.scala 339:64 stackmanage_35.scala 341:30]
  assign Stack_1_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1820; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1646:27]
  assign Stack_1_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1819; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1645:28]
  assign Stack_2_clock = clock;
  assign Stack_2_reset = reset;
  assign Stack_2_io_push = LUT_stack_io_push_2; // @[stackmanage_35.scala 151:37]
  assign Stack_2_io_pop = LUT_stack_io_pop_2; // @[stackmanage_35.scala 112:38]
  assign Stack_2_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_596); // @[stackmanage_35.scala 339:64 stackmanage_35.scala 342:30]
  assign Stack_2_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1823; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1648:27]
  assign Stack_2_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1822; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1647:28]
  assign Stack_3_clock = clock;
  assign Stack_3_reset = reset;
  assign Stack_3_io_push = LUT_stack_io_push_3; // @[stackmanage_35.scala 152:37]
  assign Stack_3_io_pop = LUT_stack_io_pop_3; // @[stackmanage_35.scala 113:38]
  assign Stack_3_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_597); // @[stackmanage_35.scala 339:64 stackmanage_35.scala 343:30]
  assign Stack_3_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1825; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1650:27]
  assign Stack_3_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1824; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1649:28]
  assign Stack_4_clock = clock;
  assign Stack_4_reset = reset;
  assign Stack_4_io_push = LUT_stack_io_push_4; // @[stackmanage_35.scala 153:37]
  assign Stack_4_io_pop = LUT_stack_io_pop_4; // @[stackmanage_35.scala 114:38]
  assign Stack_4_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_598); // @[stackmanage_35.scala 339:64 stackmanage_35.scala 344:30]
  assign Stack_4_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1827; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1652:27]
  assign Stack_4_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1826; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1651:28]
  assign Stack_5_clock = clock;
  assign Stack_5_reset = reset;
  assign Stack_5_io_push = LUT_stack_io_push_5; // @[stackmanage_35.scala 154:37]
  assign Stack_5_io_pop = LUT_stack_io_pop_5; // @[stackmanage_35.scala 115:38]
  assign Stack_5_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_599); // @[stackmanage_35.scala 339:64 stackmanage_35.scala 345:30]
  assign Stack_5_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1829; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1654:27]
  assign Stack_5_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1828; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1653:28]
  assign Stack_6_clock = clock;
  assign Stack_6_reset = reset;
  assign Stack_6_io_push = LUT_stack_io_push_6; // @[stackmanage_35.scala 155:37]
  assign Stack_6_io_pop = LUT_stack_io_pop_6; // @[stackmanage_35.scala 116:38]
  assign Stack_6_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_600); // @[stackmanage_35.scala 339:64 stackmanage_35.scala 346:30]
  assign Stack_6_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1831; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1656:27]
  assign Stack_6_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1830; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1655:28]
  assign Stack_7_clock = clock;
  assign Stack_7_reset = reset;
  assign Stack_7_io_push = LUT_stack_io_push_7; // @[stackmanage_35.scala 156:37]
  assign Stack_7_io_pop = LUT_stack_io_pop_7; // @[stackmanage_35.scala 117:38]
  assign Stack_7_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_601); // @[stackmanage_35.scala 339:64 stackmanage_35.scala 347:30]
  assign Stack_7_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1833; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1658:27]
  assign Stack_7_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1832; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1657:28]
  assign Stack_8_clock = clock;
  assign Stack_8_reset = reset;
  assign Stack_8_io_push = LUT_stack_io_push_8; // @[stackmanage_35.scala 157:37]
  assign Stack_8_io_pop = LUT_stack_io_pop_8; // @[stackmanage_35.scala 118:38]
  assign Stack_8_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_602); // @[stackmanage_35.scala 339:64 stackmanage_35.scala 348:30]
  assign Stack_8_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1835; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1660:27]
  assign Stack_8_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1834; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1659:28]
  assign Stack_9_clock = clock;
  assign Stack_9_reset = reset;
  assign Stack_9_io_push = LUT_stack_io_push_9; // @[stackmanage_35.scala 158:37]
  assign Stack_9_io_pop = LUT_stack_io_pop_9; // @[stackmanage_35.scala 119:38]
  assign Stack_9_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_603); // @[stackmanage_35.scala 339:64 stackmanage_35.scala 349:30]
  assign Stack_9_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1837; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1662:27]
  assign Stack_9_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1836; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1661:28]
  assign Stack_10_clock = clock;
  assign Stack_10_reset = reset;
  assign Stack_10_io_push = LUT_stack_io_push_10; // @[stackmanage_35.scala 160:38]
  assign Stack_10_io_pop = LUT_stack_io_pop_10; // @[stackmanage_35.scala 121:39]
  assign Stack_10_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_604); // @[stackmanage_35.scala 339:64 stackmanage_35.scala 350:31]
  assign Stack_10_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1839; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1664:29]
  assign Stack_10_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1838; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1663:29]
  assign Stack_11_clock = clock;
  assign Stack_11_reset = reset;
  assign Stack_11_io_push = LUT_stack_io_push_11; // @[stackmanage_35.scala 161:38]
  assign Stack_11_io_pop = LUT_stack_io_pop_11; // @[stackmanage_35.scala 122:39]
  assign Stack_11_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_605); // @[stackmanage_35.scala 339:64 stackmanage_35.scala 351:31]
  assign Stack_11_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1841; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1666:28]
  assign Stack_11_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1840; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1665:29]
  assign Stack_12_clock = clock;
  assign Stack_12_reset = reset;
  assign Stack_12_io_push = LUT_stack_io_push_12; // @[stackmanage_35.scala 162:38]
  assign Stack_12_io_pop = LUT_stack_io_pop_12; // @[stackmanage_35.scala 123:39]
  assign Stack_12_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_606); // @[stackmanage_35.scala 339:64 stackmanage_35.scala 352:31]
  assign Stack_12_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1843; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1668:28]
  assign Stack_12_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1842; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1667:29]
  assign Stack_13_clock = clock;
  assign Stack_13_reset = reset;
  assign Stack_13_io_push = LUT_stack_io_push_13; // @[stackmanage_35.scala 163:38]
  assign Stack_13_io_pop = LUT_stack_io_pop_13; // @[stackmanage_35.scala 124:39]
  assign Stack_13_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_607); // @[stackmanage_35.scala 339:64 stackmanage_35.scala 353:31]
  assign Stack_13_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1845; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1670:28]
  assign Stack_13_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1844; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1669:29]
  assign Stack_14_clock = clock;
  assign Stack_14_reset = reset;
  assign Stack_14_io_push = LUT_stack_io_push_14; // @[stackmanage_35.scala 164:38]
  assign Stack_14_io_pop = LUT_stack_io_pop_14; // @[stackmanage_35.scala 125:39]
  assign Stack_14_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_608); // @[stackmanage_35.scala 339:64 stackmanage_35.scala 354:31]
  assign Stack_14_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1847; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1672:28]
  assign Stack_14_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1846; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1671:29]
  assign Stack_15_clock = clock;
  assign Stack_15_reset = reset;
  assign Stack_15_io_push = LUT_stack_io_push_15; // @[stackmanage_35.scala 165:38]
  assign Stack_15_io_pop = LUT_stack_io_pop_15; // @[stackmanage_35.scala 126:39]
  assign Stack_15_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_609); // @[stackmanage_35.scala 339:64 stackmanage_35.scala 355:31]
  assign Stack_15_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1849; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1674:28]
  assign Stack_15_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1848; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1673:29]
  assign Stack_16_clock = clock;
  assign Stack_16_reset = reset;
  assign Stack_16_io_push = LUT_stack_io_push_16; // @[stackmanage_35.scala 166:38]
  assign Stack_16_io_pop = LUT_stack_io_pop_16; // @[stackmanage_35.scala 127:39]
  assign Stack_16_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_610); // @[stackmanage_35.scala 339:64 stackmanage_35.scala 356:31]
  assign Stack_16_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1851; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1676:28]
  assign Stack_16_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1850; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1675:29]
  assign Stack_17_clock = clock;
  assign Stack_17_reset = reset;
  assign Stack_17_io_push = LUT_stack_io_push_17; // @[stackmanage_35.scala 167:38]
  assign Stack_17_io_pop = LUT_stack_io_pop_17; // @[stackmanage_35.scala 128:39]
  assign Stack_17_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_611); // @[stackmanage_35.scala 339:64 stackmanage_35.scala 357:31]
  assign Stack_17_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1853; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1678:28]
  assign Stack_17_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1852; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1677:29]
  assign Stack_18_clock = clock;
  assign Stack_18_reset = reset;
  assign Stack_18_io_push = LUT_stack_io_push_18; // @[stackmanage_35.scala 168:38]
  assign Stack_18_io_pop = LUT_stack_io_pop_18; // @[stackmanage_35.scala 129:39]
  assign Stack_18_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_612); // @[stackmanage_35.scala 339:64 stackmanage_35.scala 358:31]
  assign Stack_18_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1855; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1680:28]
  assign Stack_18_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1854; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1679:29]
  assign Stack_19_clock = clock;
  assign Stack_19_reset = reset;
  assign Stack_19_io_push = LUT_stack_io_push_19; // @[stackmanage_35.scala 169:38]
  assign Stack_19_io_pop = LUT_stack_io_pop_19; // @[stackmanage_35.scala 130:39]
  assign Stack_19_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_613); // @[stackmanage_35.scala 339:64 stackmanage_35.scala 359:31]
  assign Stack_19_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1857; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1682:28]
  assign Stack_19_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1856; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1681:29]
  assign Stack_20_clock = clock;
  assign Stack_20_reset = reset;
  assign Stack_20_io_push = LUT_stack_io_push_20; // @[stackmanage_35.scala 171:38]
  assign Stack_20_io_pop = LUT_stack_io_pop_20; // @[stackmanage_35.scala 132:39]
  assign Stack_20_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_614); // @[stackmanage_35.scala 339:64 stackmanage_35.scala 360:31]
  assign Stack_20_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1859; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1684:29]
  assign Stack_20_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1858; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1683:29]
  assign Stack_21_clock = clock;
  assign Stack_21_reset = reset;
  assign Stack_21_io_push = LUT_stack_io_push_21; // @[stackmanage_35.scala 172:38]
  assign Stack_21_io_pop = LUT_stack_io_pop_21; // @[stackmanage_35.scala 133:39]
  assign Stack_21_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_615); // @[stackmanage_35.scala 339:64 stackmanage_35.scala 361:31]
  assign Stack_21_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1861; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1686:28]
  assign Stack_21_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1860; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1685:29]
  assign Stack_22_clock = clock;
  assign Stack_22_reset = reset;
  assign Stack_22_io_push = LUT_stack_io_push_22; // @[stackmanage_35.scala 173:38]
  assign Stack_22_io_pop = LUT_stack_io_pop_22; // @[stackmanage_35.scala 134:39]
  assign Stack_22_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_616); // @[stackmanage_35.scala 339:64 stackmanage_35.scala 362:31]
  assign Stack_22_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1863; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1688:28]
  assign Stack_22_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1862; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1687:29]
  assign Stack_23_clock = clock;
  assign Stack_23_reset = reset;
  assign Stack_23_io_push = LUT_stack_io_push_23; // @[stackmanage_35.scala 174:38]
  assign Stack_23_io_pop = LUT_stack_io_pop_23; // @[stackmanage_35.scala 135:39]
  assign Stack_23_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_617); // @[stackmanage_35.scala 339:64 stackmanage_35.scala 363:31]
  assign Stack_23_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1865; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1690:28]
  assign Stack_23_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1864; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1689:29]
  assign Stack_24_clock = clock;
  assign Stack_24_reset = reset;
  assign Stack_24_io_push = LUT_stack_io_push_24; // @[stackmanage_35.scala 175:38]
  assign Stack_24_io_pop = LUT_stack_io_pop_24; // @[stackmanage_35.scala 136:39]
  assign Stack_24_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_618); // @[stackmanage_35.scala 339:64 stackmanage_35.scala 364:31]
  assign Stack_24_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1867; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1692:28]
  assign Stack_24_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1866; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1691:29]
  assign Stack_25_clock = clock;
  assign Stack_25_reset = reset;
  assign Stack_25_io_push = LUT_stack_io_push_25; // @[stackmanage_35.scala 176:38]
  assign Stack_25_io_pop = LUT_stack_io_pop_25; // @[stackmanage_35.scala 137:39]
  assign Stack_25_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_619); // @[stackmanage_35.scala 339:64 stackmanage_35.scala 365:31]
  assign Stack_25_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1869; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1694:28]
  assign Stack_25_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1868; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1693:29]
  assign Stack_26_clock = clock;
  assign Stack_26_reset = reset;
  assign Stack_26_io_push = LUT_stack_io_push_26; // @[stackmanage_35.scala 177:38]
  assign Stack_26_io_pop = LUT_stack_io_pop_26; // @[stackmanage_35.scala 138:39]
  assign Stack_26_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_620); // @[stackmanage_35.scala 339:64 stackmanage_35.scala 366:31]
  assign Stack_26_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1871; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1696:28]
  assign Stack_26_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1870; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1695:29]
  assign Stack_27_clock = clock;
  assign Stack_27_reset = reset;
  assign Stack_27_io_push = LUT_stack_io_push_27; // @[stackmanage_35.scala 178:38]
  assign Stack_27_io_pop = LUT_stack_io_pop_27; // @[stackmanage_35.scala 139:39]
  assign Stack_27_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_621); // @[stackmanage_35.scala 339:64 stackmanage_35.scala 367:31]
  assign Stack_27_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1873; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1698:28]
  assign Stack_27_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1872; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1697:29]
  assign Stack_28_clock = clock;
  assign Stack_28_reset = reset;
  assign Stack_28_io_push = LUT_stack_io_push_28; // @[stackmanage_35.scala 179:38]
  assign Stack_28_io_pop = LUT_stack_io_pop_28; // @[stackmanage_35.scala 140:39]
  assign Stack_28_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_622); // @[stackmanage_35.scala 339:64 stackmanage_35.scala 368:31]
  assign Stack_28_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1875; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1700:28]
  assign Stack_28_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1874; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1699:29]
  assign Stack_29_clock = clock;
  assign Stack_29_reset = reset;
  assign Stack_29_io_push = LUT_stack_io_push_29; // @[stackmanage_35.scala 180:38]
  assign Stack_29_io_pop = LUT_stack_io_pop_29; // @[stackmanage_35.scala 141:39]
  assign Stack_29_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_623); // @[stackmanage_35.scala 339:64 stackmanage_35.scala 369:31]
  assign Stack_29_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1877; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1702:28]
  assign Stack_29_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1876; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1701:29]
  assign Stack_30_clock = clock;
  assign Stack_30_reset = reset;
  assign Stack_30_io_push = LUT_stack_io_push_30; // @[stackmanage_35.scala 182:38]
  assign Stack_30_io_pop = LUT_stack_io_pop_30; // @[stackmanage_35.scala 143:39]
  assign Stack_30_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_624); // @[stackmanage_35.scala 339:64 stackmanage_35.scala 370:31]
  assign Stack_30_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1879; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1704:29]
  assign Stack_30_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1878; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1703:29]
  assign Stack_31_clock = clock;
  assign Stack_31_reset = reset;
  assign Stack_31_io_push = LUT_stack_io_push_31; // @[stackmanage_35.scala 183:38]
  assign Stack_31_io_pop = LUT_stack_io_pop_31; // @[stackmanage_35.scala 144:39]
  assign Stack_31_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_625); // @[stackmanage_35.scala 339:64 stackmanage_35.scala 371:31]
  assign Stack_31_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1881; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1706:28]
  assign Stack_31_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1880; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1705:29]
  assign Stack_32_clock = clock;
  assign Stack_32_reset = reset;
  assign Stack_32_io_push = LUT_stack_io_push_32; // @[stackmanage_35.scala 184:38]
  assign Stack_32_io_pop = LUT_stack_io_pop_32; // @[stackmanage_35.scala 145:39]
  assign Stack_32_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_626); // @[stackmanage_35.scala 339:64 stackmanage_35.scala 372:31]
  assign Stack_32_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1883; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1708:28]
  assign Stack_32_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1882; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1707:29]
  assign Stack_33_clock = clock;
  assign Stack_33_reset = reset;
  assign Stack_33_io_push = LUT_stack_io_push_33; // @[stackmanage_35.scala 185:38]
  assign Stack_33_io_pop = LUT_stack_io_pop_33; // @[stackmanage_35.scala 146:39]
  assign Stack_33_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_627); // @[stackmanage_35.scala 339:64 stackmanage_35.scala 373:31]
  assign Stack_33_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1885; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1710:28]
  assign Stack_33_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1884; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1709:29]
  assign Stack_34_clock = clock;
  assign Stack_34_reset = reset;
  assign Stack_34_io_push = LUT_stack_io_push_34; // @[stackmanage_35.scala 186:38]
  assign Stack_34_io_pop = LUT_stack_io_pop_34; // @[stackmanage_35.scala 147:39]
  assign Stack_34_io_dataIn = LUT_stack_io_push_0 & LUT_stack_io_push_en ? $signed(32'sh0) : $signed(_GEN_628); // @[stackmanage_35.scala 339:64 stackmanage_35.scala 374:31]
  assign Stack_34_io_ray_id = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1887; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1712:28]
  assign Stack_34_io_hit_in = LUT_stack_io_pop_en & LUT_stack_io_pop_0 ? 32'h0 : _GEN_1886; // @[stackmanage_35.scala 1642:63 stackmanage_35.scala 1711:29]
  always @(posedge clock) begin
    if (reset) begin // @[stackmanage_35.scala 331:34]
      node_push_in_1 <= 32'sh0; // @[stackmanage_35.scala 331:34]
    end else begin
      node_push_in_1 <= LUT_stack_io_node_id_push_in; // @[stackmanage_35.scala 335:29]
    end
    if (reset) begin // @[stackmanage_35.scala 332:34]
      node_push_in_2 <= 32'sh0; // @[stackmanage_35.scala 332:34]
    end else begin
      node_push_in_2 <= node_push_in_1; // @[stackmanage_35.scala 336:29]
    end
    if (reset) begin // @[stackmanage_35.scala 1638:34]
      hitT_out_temp <= 32'h0; // @[stackmanage_35.scala 1638:34]
    end else if (pop_0 & Stack_0_io_enable) begin // @[stackmanage_35.scala 4288:48]
      hitT_out_temp <= Stack_0_io_hit_out; // @[stackmanage_35.scala 4290:27]
    end else if (pop_1 & Stack_1_io_enable) begin // @[stackmanage_35.scala 4294:53]
      hitT_out_temp <= Stack_1_io_hit_out; // @[stackmanage_35.scala 4295:27]
    end else if (pop_2 & Stack_2_io_enable) begin // @[stackmanage_35.scala 4299:53]
      hitT_out_temp <= Stack_2_io_hit_out; // @[stackmanage_35.scala 4300:27]
    end else begin
      hitT_out_temp <= _GEN_2082;
    end
    if (reset) begin // @[stackmanage_35.scala 1639:35]
      ray_out_temp <= 32'h0; // @[stackmanage_35.scala 1639:35]
    end else if (pop_0 & Stack_0_io_enable) begin // @[stackmanage_35.scala 4288:48]
      ray_out_temp <= Stack_0_io_ray_out; // @[stackmanage_35.scala 4291:28]
    end else if (pop_1 & Stack_1_io_enable) begin // @[stackmanage_35.scala 4294:53]
      ray_out_temp <= Stack_1_io_ray_out; // @[stackmanage_35.scala 4296:28]
    end else if (pop_2 & Stack_2_io_enable) begin // @[stackmanage_35.scala 4299:53]
      ray_out_temp <= Stack_2_io_ray_out; // @[stackmanage_35.scala 4301:28]
    end else begin
      ray_out_temp <= _GEN_2083;
    end
    if (reset) begin // @[stackmanage_35.scala 1640:32]
      node_out_temp <= 32'sh0; // @[stackmanage_35.scala 1640:32]
    end else if (pop_0 & Stack_0_io_enable) begin // @[stackmanage_35.scala 4288:48]
      node_out_temp <= Stack_0_io_dataOut; // @[stackmanage_35.scala 4292:25]
    end else if (pop_1 & Stack_1_io_enable) begin // @[stackmanage_35.scala 4294:53]
      node_out_temp <= Stack_1_io_dataOut; // @[stackmanage_35.scala 4297:25]
    end else if (pop_2 & Stack_2_io_enable) begin // @[stackmanage_35.scala 4299:53]
      node_out_temp <= Stack_2_io_dataOut; // @[stackmanage_35.scala 4302:25]
    end else begin
      node_out_temp <= _GEN_2084;
    end
    if (reset) begin // @[stackmanage_35.scala 1641:38]
      pop_valid_1 <= 1'h0; // @[stackmanage_35.scala 1641:38]
    end else begin
      pop_valid_1 <= _GEN_2097;
    end
    if (reset) begin // @[stackmanage_35.scala 4201:46]
      pop_0 <= 1'h0; // @[stackmanage_35.scala 4201:46]
    end else begin
      pop_0 <= LUT_stack_io_pop_0; // @[stackmanage_35.scala 4251:40]
    end
    if (reset) begin // @[stackmanage_35.scala 4202:46]
      pop_1 <= 1'h0; // @[stackmanage_35.scala 4202:46]
    end else begin
      pop_1 <= LUT_stack_io_pop_1; // @[stackmanage_35.scala 4252:40]
    end
    if (reset) begin // @[stackmanage_35.scala 4203:46]
      pop_2 <= 1'h0; // @[stackmanage_35.scala 4203:46]
    end else begin
      pop_2 <= LUT_stack_io_pop_2; // @[stackmanage_35.scala 4253:40]
    end
    if (reset) begin // @[stackmanage_35.scala 4204:46]
      pop_3 <= 1'h0; // @[stackmanage_35.scala 4204:46]
    end else begin
      pop_3 <= LUT_stack_io_pop_3; // @[stackmanage_35.scala 4254:40]
    end
    if (reset) begin // @[stackmanage_35.scala 4205:46]
      pop_4 <= 1'h0; // @[stackmanage_35.scala 4205:46]
    end else begin
      pop_4 <= LUT_stack_io_pop_4; // @[stackmanage_35.scala 4255:40]
    end
    if (reset) begin // @[stackmanage_35.scala 4206:46]
      pop_5 <= 1'h0; // @[stackmanage_35.scala 4206:46]
    end else begin
      pop_5 <= LUT_stack_io_pop_5; // @[stackmanage_35.scala 4256:40]
    end
    if (reset) begin // @[stackmanage_35.scala 4207:46]
      pop_6 <= 1'h0; // @[stackmanage_35.scala 4207:46]
    end else begin
      pop_6 <= LUT_stack_io_pop_6; // @[stackmanage_35.scala 4257:40]
    end
    if (reset) begin // @[stackmanage_35.scala 4208:46]
      pop_7 <= 1'h0; // @[stackmanage_35.scala 4208:46]
    end else begin
      pop_7 <= LUT_stack_io_pop_7; // @[stackmanage_35.scala 4258:40]
    end
    if (reset) begin // @[stackmanage_35.scala 4209:46]
      pop_8 <= 1'h0; // @[stackmanage_35.scala 4209:46]
    end else begin
      pop_8 <= LUT_stack_io_pop_8; // @[stackmanage_35.scala 4259:40]
    end
    if (reset) begin // @[stackmanage_35.scala 4210:46]
      pop_9 <= 1'h0; // @[stackmanage_35.scala 4210:46]
    end else begin
      pop_9 <= LUT_stack_io_pop_9; // @[stackmanage_35.scala 4260:40]
    end
    if (reset) begin // @[stackmanage_35.scala 4212:47]
      pop_10 <= 1'h0; // @[stackmanage_35.scala 4212:47]
    end else begin
      pop_10 <= LUT_stack_io_pop_10; // @[stackmanage_35.scala 4261:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4213:47]
      pop_11 <= 1'h0; // @[stackmanage_35.scala 4213:47]
    end else begin
      pop_11 <= LUT_stack_io_pop_11; // @[stackmanage_35.scala 4262:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4214:47]
      pop_12 <= 1'h0; // @[stackmanage_35.scala 4214:47]
    end else begin
      pop_12 <= LUT_stack_io_pop_12; // @[stackmanage_35.scala 4263:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4215:47]
      pop_13 <= 1'h0; // @[stackmanage_35.scala 4215:47]
    end else begin
      pop_13 <= LUT_stack_io_pop_13; // @[stackmanage_35.scala 4264:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4216:47]
      pop_14 <= 1'h0; // @[stackmanage_35.scala 4216:47]
    end else begin
      pop_14 <= LUT_stack_io_pop_14; // @[stackmanage_35.scala 4265:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4217:47]
      pop_15 <= 1'h0; // @[stackmanage_35.scala 4217:47]
    end else begin
      pop_15 <= LUT_stack_io_pop_15; // @[stackmanage_35.scala 4266:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4218:47]
      pop_16 <= 1'h0; // @[stackmanage_35.scala 4218:47]
    end else begin
      pop_16 <= LUT_stack_io_pop_16; // @[stackmanage_35.scala 4267:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4219:47]
      pop_17 <= 1'h0; // @[stackmanage_35.scala 4219:47]
    end else begin
      pop_17 <= LUT_stack_io_pop_17; // @[stackmanage_35.scala 4268:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4220:47]
      pop_18 <= 1'h0; // @[stackmanage_35.scala 4220:47]
    end else begin
      pop_18 <= LUT_stack_io_pop_18; // @[stackmanage_35.scala 4269:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4221:47]
      pop_19 <= 1'h0; // @[stackmanage_35.scala 4221:47]
    end else begin
      pop_19 <= LUT_stack_io_pop_19; // @[stackmanage_35.scala 4270:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4223:47]
      pop_20 <= 1'h0; // @[stackmanage_35.scala 4223:47]
    end else begin
      pop_20 <= LUT_stack_io_pop_20; // @[stackmanage_35.scala 4271:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4224:47]
      pop_21 <= 1'h0; // @[stackmanage_35.scala 4224:47]
    end else begin
      pop_21 <= LUT_stack_io_pop_21; // @[stackmanage_35.scala 4272:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4225:47]
      pop_22 <= 1'h0; // @[stackmanage_35.scala 4225:47]
    end else begin
      pop_22 <= LUT_stack_io_pop_22; // @[stackmanage_35.scala 4273:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4226:47]
      pop_23 <= 1'h0; // @[stackmanage_35.scala 4226:47]
    end else begin
      pop_23 <= LUT_stack_io_pop_23; // @[stackmanage_35.scala 4274:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4227:47]
      pop_24 <= 1'h0; // @[stackmanage_35.scala 4227:47]
    end else begin
      pop_24 <= LUT_stack_io_pop_24; // @[stackmanage_35.scala 4275:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4228:47]
      pop_25 <= 1'h0; // @[stackmanage_35.scala 4228:47]
    end else begin
      pop_25 <= LUT_stack_io_pop_25; // @[stackmanage_35.scala 4276:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4229:47]
      pop_26 <= 1'h0; // @[stackmanage_35.scala 4229:47]
    end else begin
      pop_26 <= LUT_stack_io_pop_26; // @[stackmanage_35.scala 4277:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4230:47]
      pop_27 <= 1'h0; // @[stackmanage_35.scala 4230:47]
    end else begin
      pop_27 <= LUT_stack_io_pop_27; // @[stackmanage_35.scala 4278:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4231:47]
      pop_28 <= 1'h0; // @[stackmanage_35.scala 4231:47]
    end else begin
      pop_28 <= LUT_stack_io_pop_28; // @[stackmanage_35.scala 4279:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4232:47]
      pop_29 <= 1'h0; // @[stackmanage_35.scala 4232:47]
    end else begin
      pop_29 <= LUT_stack_io_pop_29; // @[stackmanage_35.scala 4280:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4234:47]
      pop_30 <= 1'h0; // @[stackmanage_35.scala 4234:47]
    end else begin
      pop_30 <= LUT_stack_io_pop_30; // @[stackmanage_35.scala 4281:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4235:47]
      pop_31 <= 1'h0; // @[stackmanage_35.scala 4235:47]
    end else begin
      pop_31 <= LUT_stack_io_pop_31; // @[stackmanage_35.scala 4282:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4236:47]
      pop_32 <= 1'h0; // @[stackmanage_35.scala 4236:47]
    end else begin
      pop_32 <= LUT_stack_io_pop_32; // @[stackmanage_35.scala 4283:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4237:47]
      pop_33 <= 1'h0; // @[stackmanage_35.scala 4237:47]
    end else begin
      pop_33 <= LUT_stack_io_pop_33; // @[stackmanage_35.scala 4284:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4238:47]
      pop_34 <= 1'h0; // @[stackmanage_35.scala 4238:47]
    end else begin
      pop_34 <= LUT_stack_io_pop_34; // @[stackmanage_35.scala 4285:41]
    end
    if (reset) begin // @[stackmanage_35.scala 4476:41]
      dispatch_0 <= 1'h0; // @[stackmanage_35.scala 4476:41]
    end else begin
      dispatch_0 <= _T_317;
    end
    if (reset) begin // @[stackmanage_35.scala 4477:41]
      dispatch_1 <= 1'h0; // @[stackmanage_35.scala 4477:41]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4599:38]
      dispatch_1 <= 1'h0; // @[stackmanage_35.scala 4601:33]
    end else begin
      dispatch_1 <= _T_320;
    end
    if (reset) begin // @[stackmanage_35.scala 4478:41]
      dispatch_2 <= 1'h0; // @[stackmanage_35.scala 4478:41]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4599:38]
      dispatch_2 <= 1'h0; // @[stackmanage_35.scala 4602:33]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4635:43]
      dispatch_2 <= 1'h0; // @[stackmanage_35.scala 4638:33]
    end else begin
      dispatch_2 <= _T_323;
    end
    if (reset) begin // @[stackmanage_35.scala 4479:41]
      dispatch_3 <= 1'h0; // @[stackmanage_35.scala 4479:41]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4599:38]
      dispatch_3 <= 1'h0; // @[stackmanage_35.scala 4603:33]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4635:43]
      dispatch_3 <= 1'h0; // @[stackmanage_35.scala 4639:33]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4672:43]
      dispatch_3 <= 1'h0; // @[stackmanage_35.scala 4676:33]
    end else begin
      dispatch_3 <= _T_326;
    end
    if (reset) begin // @[stackmanage_35.scala 4480:41]
      dispatch_4 <= 1'h0; // @[stackmanage_35.scala 4480:41]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4599:38]
      dispatch_4 <= 1'h0; // @[stackmanage_35.scala 4604:33]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4635:43]
      dispatch_4 <= 1'h0; // @[stackmanage_35.scala 4640:33]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4672:43]
      dispatch_4 <= 1'h0; // @[stackmanage_35.scala 4678:33]
    end else begin
      dispatch_4 <= _GEN_2627;
    end
    if (reset) begin // @[stackmanage_35.scala 4481:41]
      dispatch_5 <= 1'h0; // @[stackmanage_35.scala 4481:41]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4599:38]
      dispatch_5 <= 1'h0; // @[stackmanage_35.scala 4605:33]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4635:43]
      dispatch_5 <= 1'h0; // @[stackmanage_35.scala 4641:33]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4672:43]
      dispatch_5 <= 1'h0; // @[stackmanage_35.scala 4679:33]
    end else begin
      dispatch_5 <= _GEN_2628;
    end
    if (reset) begin // @[stackmanage_35.scala 4482:41]
      dispatch_6 <= 1'h0; // @[stackmanage_35.scala 4482:41]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4599:38]
      dispatch_6 <= 1'h0; // @[stackmanage_35.scala 4606:33]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4635:43]
      dispatch_6 <= 1'h0; // @[stackmanage_35.scala 4642:33]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4672:43]
      dispatch_6 <= 1'h0; // @[stackmanage_35.scala 4680:33]
    end else begin
      dispatch_6 <= _GEN_2629;
    end
    if (reset) begin // @[stackmanage_35.scala 4483:41]
      dispatch_7 <= 1'h0; // @[stackmanage_35.scala 4483:41]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4599:38]
      dispatch_7 <= 1'h0; // @[stackmanage_35.scala 4607:33]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4635:43]
      dispatch_7 <= 1'h0; // @[stackmanage_35.scala 4643:33]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4672:43]
      dispatch_7 <= 1'h0; // @[stackmanage_35.scala 4681:33]
    end else begin
      dispatch_7 <= _GEN_2630;
    end
    if (reset) begin // @[stackmanage_35.scala 4484:41]
      dispatch_8 <= 1'h0; // @[stackmanage_35.scala 4484:41]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4599:38]
      dispatch_8 <= 1'h0; // @[stackmanage_35.scala 4608:33]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4635:43]
      dispatch_8 <= 1'h0; // @[stackmanage_35.scala 4644:33]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4672:43]
      dispatch_8 <= 1'h0; // @[stackmanage_35.scala 4682:33]
    end else begin
      dispatch_8 <= _GEN_2631;
    end
    if (reset) begin // @[stackmanage_35.scala 4485:41]
      dispatch_9 <= 1'h0; // @[stackmanage_35.scala 4485:41]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4599:38]
      dispatch_9 <= 1'h0; // @[stackmanage_35.scala 4609:33]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4635:43]
      dispatch_9 <= 1'h0; // @[stackmanage_35.scala 4645:33]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4672:43]
      dispatch_9 <= 1'h0; // @[stackmanage_35.scala 4683:33]
    end else begin
      dispatch_9 <= _GEN_2632;
    end
    if (reset) begin // @[stackmanage_35.scala 4487:42]
      dispatch_10 <= 1'h0; // @[stackmanage_35.scala 4487:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4599:38]
      dispatch_10 <= 1'h0; // @[stackmanage_35.scala 4610:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4635:43]
      dispatch_10 <= 1'h0; // @[stackmanage_35.scala 4646:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4672:43]
      dispatch_10 <= 1'h0; // @[stackmanage_35.scala 4684:34]
    end else begin
      dispatch_10 <= _GEN_2633;
    end
    if (reset) begin // @[stackmanage_35.scala 4488:42]
      dispatch_11 <= 1'h0; // @[stackmanage_35.scala 4488:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4599:38]
      dispatch_11 <= 1'h0; // @[stackmanage_35.scala 4611:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4635:43]
      dispatch_11 <= 1'h0; // @[stackmanage_35.scala 4647:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4672:43]
      dispatch_11 <= 1'h0; // @[stackmanage_35.scala 4685:34]
    end else begin
      dispatch_11 <= _GEN_2634;
    end
    if (reset) begin // @[stackmanage_35.scala 4489:42]
      dispatch_12 <= 1'h0; // @[stackmanage_35.scala 4489:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4599:38]
      dispatch_12 <= 1'h0; // @[stackmanage_35.scala 4612:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4635:43]
      dispatch_12 <= 1'h0; // @[stackmanage_35.scala 4648:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4672:43]
      dispatch_12 <= 1'h0; // @[stackmanage_35.scala 4686:34]
    end else begin
      dispatch_12 <= _GEN_2635;
    end
    if (reset) begin // @[stackmanage_35.scala 4490:42]
      dispatch_13 <= 1'h0; // @[stackmanage_35.scala 4490:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4599:38]
      dispatch_13 <= 1'h0; // @[stackmanage_35.scala 4613:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4635:43]
      dispatch_13 <= 1'h0; // @[stackmanage_35.scala 4649:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4672:43]
      dispatch_13 <= 1'h0; // @[stackmanage_35.scala 4687:34]
    end else begin
      dispatch_13 <= _GEN_2636;
    end
    if (reset) begin // @[stackmanage_35.scala 4491:42]
      dispatch_14 <= 1'h0; // @[stackmanage_35.scala 4491:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4599:38]
      dispatch_14 <= 1'h0; // @[stackmanage_35.scala 4614:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4635:43]
      dispatch_14 <= 1'h0; // @[stackmanage_35.scala 4650:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4672:43]
      dispatch_14 <= 1'h0; // @[stackmanage_35.scala 4688:34]
    end else begin
      dispatch_14 <= _GEN_2637;
    end
    if (reset) begin // @[stackmanage_35.scala 4492:42]
      dispatch_15 <= 1'h0; // @[stackmanage_35.scala 4492:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4599:38]
      dispatch_15 <= 1'h0; // @[stackmanage_35.scala 4615:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4635:43]
      dispatch_15 <= 1'h0; // @[stackmanage_35.scala 4651:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4672:43]
      dispatch_15 <= 1'h0; // @[stackmanage_35.scala 4689:34]
    end else begin
      dispatch_15 <= _GEN_2638;
    end
    if (reset) begin // @[stackmanage_35.scala 4493:42]
      dispatch_16 <= 1'h0; // @[stackmanage_35.scala 4493:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4599:38]
      dispatch_16 <= 1'h0; // @[stackmanage_35.scala 4616:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4635:43]
      dispatch_16 <= 1'h0; // @[stackmanage_35.scala 4652:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4672:43]
      dispatch_16 <= 1'h0; // @[stackmanage_35.scala 4690:34]
    end else begin
      dispatch_16 <= _GEN_2639;
    end
    if (reset) begin // @[stackmanage_35.scala 4494:42]
      dispatch_17 <= 1'h0; // @[stackmanage_35.scala 4494:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4599:38]
      dispatch_17 <= 1'h0; // @[stackmanage_35.scala 4617:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4635:43]
      dispatch_17 <= 1'h0; // @[stackmanage_35.scala 4653:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4672:43]
      dispatch_17 <= 1'h0; // @[stackmanage_35.scala 4691:34]
    end else begin
      dispatch_17 <= _GEN_2640;
    end
    if (reset) begin // @[stackmanage_35.scala 4495:42]
      dispatch_18 <= 1'h0; // @[stackmanage_35.scala 4495:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4599:38]
      dispatch_18 <= 1'h0; // @[stackmanage_35.scala 4618:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4635:43]
      dispatch_18 <= 1'h0; // @[stackmanage_35.scala 4654:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4672:43]
      dispatch_18 <= 1'h0; // @[stackmanage_35.scala 4692:34]
    end else begin
      dispatch_18 <= _GEN_2641;
    end
    if (reset) begin // @[stackmanage_35.scala 4496:42]
      dispatch_19 <= 1'h0; // @[stackmanage_35.scala 4496:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4599:38]
      dispatch_19 <= 1'h0; // @[stackmanage_35.scala 4619:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4635:43]
      dispatch_19 <= 1'h0; // @[stackmanage_35.scala 4655:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4672:43]
      dispatch_19 <= 1'h0; // @[stackmanage_35.scala 4693:34]
    end else begin
      dispatch_19 <= _GEN_2642;
    end
    if (reset) begin // @[stackmanage_35.scala 4498:42]
      dispatch_20 <= 1'h0; // @[stackmanage_35.scala 4498:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4599:38]
      dispatch_20 <= 1'h0; // @[stackmanage_35.scala 4620:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4635:43]
      dispatch_20 <= 1'h0; // @[stackmanage_35.scala 4656:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4672:43]
      dispatch_20 <= 1'h0; // @[stackmanage_35.scala 4694:34]
    end else begin
      dispatch_20 <= _GEN_2643;
    end
    if (reset) begin // @[stackmanage_35.scala 4499:42]
      dispatch_21 <= 1'h0; // @[stackmanage_35.scala 4499:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4599:38]
      dispatch_21 <= 1'h0; // @[stackmanage_35.scala 4621:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4635:43]
      dispatch_21 <= 1'h0; // @[stackmanage_35.scala 4657:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4672:43]
      dispatch_21 <= 1'h0; // @[stackmanage_35.scala 4695:34]
    end else begin
      dispatch_21 <= _GEN_2644;
    end
    if (reset) begin // @[stackmanage_35.scala 4500:42]
      dispatch_22 <= 1'h0; // @[stackmanage_35.scala 4500:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4599:38]
      dispatch_22 <= 1'h0; // @[stackmanage_35.scala 4622:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4635:43]
      dispatch_22 <= 1'h0; // @[stackmanage_35.scala 4658:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4672:43]
      dispatch_22 <= 1'h0; // @[stackmanage_35.scala 4696:34]
    end else begin
      dispatch_22 <= _GEN_2645;
    end
    if (reset) begin // @[stackmanage_35.scala 4501:42]
      dispatch_23 <= 1'h0; // @[stackmanage_35.scala 4501:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4599:38]
      dispatch_23 <= 1'h0; // @[stackmanage_35.scala 4623:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4635:43]
      dispatch_23 <= 1'h0; // @[stackmanage_35.scala 4659:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4672:43]
      dispatch_23 <= 1'h0; // @[stackmanage_35.scala 4697:34]
    end else begin
      dispatch_23 <= _GEN_2646;
    end
    if (reset) begin // @[stackmanage_35.scala 4502:42]
      dispatch_24 <= 1'h0; // @[stackmanage_35.scala 4502:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4599:38]
      dispatch_24 <= 1'h0; // @[stackmanage_35.scala 4624:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4635:43]
      dispatch_24 <= 1'h0; // @[stackmanage_35.scala 4660:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4672:43]
      dispatch_24 <= 1'h0; // @[stackmanage_35.scala 4698:34]
    end else begin
      dispatch_24 <= _GEN_2647;
    end
    if (reset) begin // @[stackmanage_35.scala 4503:42]
      dispatch_25 <= 1'h0; // @[stackmanage_35.scala 4503:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4599:38]
      dispatch_25 <= 1'h0; // @[stackmanage_35.scala 4625:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4635:43]
      dispatch_25 <= 1'h0; // @[stackmanage_35.scala 4661:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4672:43]
      dispatch_25 <= 1'h0; // @[stackmanage_35.scala 4699:34]
    end else begin
      dispatch_25 <= _GEN_2648;
    end
    if (reset) begin // @[stackmanage_35.scala 4504:42]
      dispatch_26 <= 1'h0; // @[stackmanage_35.scala 4504:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4599:38]
      dispatch_26 <= 1'h0; // @[stackmanage_35.scala 4626:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4635:43]
      dispatch_26 <= 1'h0; // @[stackmanage_35.scala 4662:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4672:43]
      dispatch_26 <= 1'h0; // @[stackmanage_35.scala 4700:34]
    end else begin
      dispatch_26 <= _GEN_2649;
    end
    if (reset) begin // @[stackmanage_35.scala 4505:42]
      dispatch_27 <= 1'h0; // @[stackmanage_35.scala 4505:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4599:38]
      dispatch_27 <= 1'h0; // @[stackmanage_35.scala 4627:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4635:43]
      dispatch_27 <= 1'h0; // @[stackmanage_35.scala 4663:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4672:43]
      dispatch_27 <= 1'h0; // @[stackmanage_35.scala 4701:34]
    end else begin
      dispatch_27 <= _GEN_2650;
    end
    if (reset) begin // @[stackmanage_35.scala 4506:42]
      dispatch_28 <= 1'h0; // @[stackmanage_35.scala 4506:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4599:38]
      dispatch_28 <= 1'h0; // @[stackmanage_35.scala 4628:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4635:43]
      dispatch_28 <= 1'h0; // @[stackmanage_35.scala 4664:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4672:43]
      dispatch_28 <= 1'h0; // @[stackmanage_35.scala 4702:34]
    end else begin
      dispatch_28 <= _GEN_2651;
    end
    if (reset) begin // @[stackmanage_35.scala 4507:42]
      dispatch_29 <= 1'h0; // @[stackmanage_35.scala 4507:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4599:38]
      dispatch_29 <= 1'h0; // @[stackmanage_35.scala 4629:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4635:43]
      dispatch_29 <= 1'h0; // @[stackmanage_35.scala 4665:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4672:43]
      dispatch_29 <= 1'h0; // @[stackmanage_35.scala 4703:34]
    end else begin
      dispatch_29 <= _GEN_2652;
    end
    if (reset) begin // @[stackmanage_35.scala 4509:42]
      dispatch_30 <= 1'h0; // @[stackmanage_35.scala 4509:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4599:38]
      dispatch_30 <= 1'h0; // @[stackmanage_35.scala 4630:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4635:43]
      dispatch_30 <= 1'h0; // @[stackmanage_35.scala 4666:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4672:43]
      dispatch_30 <= 1'h0; // @[stackmanage_35.scala 4704:34]
    end else begin
      dispatch_30 <= _GEN_2653;
    end
    if (reset) begin // @[stackmanage_35.scala 4510:42]
      dispatch_31 <= 1'h0; // @[stackmanage_35.scala 4510:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4599:38]
      dispatch_31 <= 1'h0; // @[stackmanage_35.scala 4631:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4635:43]
      dispatch_31 <= 1'h0; // @[stackmanage_35.scala 4667:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4672:43]
      dispatch_31 <= 1'h0; // @[stackmanage_35.scala 4705:34]
    end else begin
      dispatch_31 <= _GEN_2654;
    end
    if (reset) begin // @[stackmanage_35.scala 4511:42]
      dispatch_32 <= 1'h0; // @[stackmanage_35.scala 4511:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4599:38]
      dispatch_32 <= 1'h0; // @[stackmanage_35.scala 4632:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4635:43]
      dispatch_32 <= 1'h0; // @[stackmanage_35.scala 4668:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4672:43]
      dispatch_32 <= 1'h0; // @[stackmanage_35.scala 4706:34]
    end else begin
      dispatch_32 <= _GEN_2655;
    end
    if (reset) begin // @[stackmanage_35.scala 4512:42]
      dispatch_33 <= 1'h0; // @[stackmanage_35.scala 4512:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4599:38]
      dispatch_33 <= 1'h0; // @[stackmanage_35.scala 4633:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4635:43]
      dispatch_33 <= 1'h0; // @[stackmanage_35.scala 4669:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4672:43]
      dispatch_33 <= 1'h0; // @[stackmanage_35.scala 4707:34]
    end else begin
      dispatch_33 <= _GEN_2656;
    end
    if (reset) begin // @[stackmanage_35.scala 4513:42]
      dispatch_34 <= 1'h0; // @[stackmanage_35.scala 4513:42]
    end else if (pop_0 & empty_0) begin // @[stackmanage_35.scala 4599:38]
      dispatch_34 <= 1'h0; // @[stackmanage_35.scala 4634:34]
    end else if (pop_1 & empty_1) begin // @[stackmanage_35.scala 4635:43]
      dispatch_34 <= 1'h0; // @[stackmanage_35.scala 4670:34]
    end else if (pop_2 & empty_2) begin // @[stackmanage_35.scala 4672:43]
      dispatch_34 <= 1'h0; // @[stackmanage_35.scala 4708:34]
    end else begin
      dispatch_34 <= _GEN_2657;
    end
    if (reset) begin // @[stackmanage_35.scala 4514:42]
      dispatch_no_match <= 1'h0; // @[stackmanage_35.scala 4514:42]
    end else begin
      dispatch_no_match <= LUT_stack_io_no_match; // @[stackmanage_35.scala 5940:25]
    end
    if (reset) begin // @[stackmanage_35.scala 4518:42]
      empty_0 <= 1'h0; // @[stackmanage_35.scala 4518:42]
    end else begin
      empty_0 <= Stack_0_io_empty; // @[stackmanage_35.scala 4557:35]
    end
    if (reset) begin // @[stackmanage_35.scala 4519:42]
      empty_1 <= 1'h0; // @[stackmanage_35.scala 4519:42]
    end else begin
      empty_1 <= Stack_1_io_empty; // @[stackmanage_35.scala 4558:35]
    end
    if (reset) begin // @[stackmanage_35.scala 4520:42]
      empty_2 <= 1'h0; // @[stackmanage_35.scala 4520:42]
    end else begin
      empty_2 <= Stack_2_io_empty; // @[stackmanage_35.scala 4559:35]
    end
    if (reset) begin // @[stackmanage_35.scala 4521:42]
      empty_3 <= 1'h0; // @[stackmanage_35.scala 4521:42]
    end else begin
      empty_3 <= Stack_3_io_empty; // @[stackmanage_35.scala 4560:35]
    end
    if (reset) begin // @[stackmanage_35.scala 4522:42]
      empty_4 <= 1'h0; // @[stackmanage_35.scala 4522:42]
    end else begin
      empty_4 <= Stack_4_io_empty; // @[stackmanage_35.scala 4561:35]
    end
    if (reset) begin // @[stackmanage_35.scala 4523:42]
      empty_5 <= 1'h0; // @[stackmanage_35.scala 4523:42]
    end else begin
      empty_5 <= Stack_5_io_empty; // @[stackmanage_35.scala 4562:35]
    end
    if (reset) begin // @[stackmanage_35.scala 4524:42]
      empty_6 <= 1'h0; // @[stackmanage_35.scala 4524:42]
    end else begin
      empty_6 <= Stack_6_io_empty; // @[stackmanage_35.scala 4563:35]
    end
    if (reset) begin // @[stackmanage_35.scala 4525:42]
      empty_7 <= 1'h0; // @[stackmanage_35.scala 4525:42]
    end else begin
      empty_7 <= Stack_7_io_empty; // @[stackmanage_35.scala 4564:35]
    end
    if (reset) begin // @[stackmanage_35.scala 4526:42]
      empty_8 <= 1'h0; // @[stackmanage_35.scala 4526:42]
    end else begin
      empty_8 <= Stack_8_io_empty; // @[stackmanage_35.scala 4565:35]
    end
    if (reset) begin // @[stackmanage_35.scala 4527:42]
      empty_9 <= 1'h0; // @[stackmanage_35.scala 4527:42]
    end else begin
      empty_9 <= Stack_9_io_empty; // @[stackmanage_35.scala 4566:35]
    end
    if (reset) begin // @[stackmanage_35.scala 4529:43]
      empty_10 <= 1'h0; // @[stackmanage_35.scala 4529:43]
    end else begin
      empty_10 <= Stack_10_io_empty; // @[stackmanage_35.scala 4568:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4530:43]
      empty_11 <= 1'h0; // @[stackmanage_35.scala 4530:43]
    end else begin
      empty_11 <= Stack_11_io_empty; // @[stackmanage_35.scala 4569:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4531:43]
      empty_12 <= 1'h0; // @[stackmanage_35.scala 4531:43]
    end else begin
      empty_12 <= Stack_12_io_empty; // @[stackmanage_35.scala 4570:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4532:43]
      empty_13 <= 1'h0; // @[stackmanage_35.scala 4532:43]
    end else begin
      empty_13 <= Stack_13_io_empty; // @[stackmanage_35.scala 4571:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4533:43]
      empty_14 <= 1'h0; // @[stackmanage_35.scala 4533:43]
    end else begin
      empty_14 <= Stack_14_io_empty; // @[stackmanage_35.scala 4572:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4534:43]
      empty_15 <= 1'h0; // @[stackmanage_35.scala 4534:43]
    end else begin
      empty_15 <= Stack_15_io_empty; // @[stackmanage_35.scala 4573:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4535:43]
      empty_16 <= 1'h0; // @[stackmanage_35.scala 4535:43]
    end else begin
      empty_16 <= Stack_16_io_empty; // @[stackmanage_35.scala 4574:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4536:43]
      empty_17 <= 1'h0; // @[stackmanage_35.scala 4536:43]
    end else begin
      empty_17 <= Stack_17_io_empty; // @[stackmanage_35.scala 4575:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4537:43]
      empty_18 <= 1'h0; // @[stackmanage_35.scala 4537:43]
    end else begin
      empty_18 <= Stack_18_io_empty; // @[stackmanage_35.scala 4576:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4538:43]
      empty_19 <= 1'h0; // @[stackmanage_35.scala 4538:43]
    end else begin
      empty_19 <= Stack_19_io_empty; // @[stackmanage_35.scala 4577:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4540:43]
      empty_20 <= 1'h0; // @[stackmanage_35.scala 4540:43]
    end else begin
      empty_20 <= Stack_20_io_empty; // @[stackmanage_35.scala 4579:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4541:43]
      empty_21 <= 1'h0; // @[stackmanage_35.scala 4541:43]
    end else begin
      empty_21 <= Stack_21_io_empty; // @[stackmanage_35.scala 4580:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4542:43]
      empty_22 <= 1'h0; // @[stackmanage_35.scala 4542:43]
    end else begin
      empty_22 <= Stack_22_io_empty; // @[stackmanage_35.scala 4581:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4543:43]
      empty_23 <= 1'h0; // @[stackmanage_35.scala 4543:43]
    end else begin
      empty_23 <= Stack_23_io_empty; // @[stackmanage_35.scala 4582:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4544:43]
      empty_24 <= 1'h0; // @[stackmanage_35.scala 4544:43]
    end else begin
      empty_24 <= Stack_24_io_empty; // @[stackmanage_35.scala 4583:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4545:43]
      empty_25 <= 1'h0; // @[stackmanage_35.scala 4545:43]
    end else begin
      empty_25 <= Stack_25_io_empty; // @[stackmanage_35.scala 4584:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4546:43]
      empty_26 <= 1'h0; // @[stackmanage_35.scala 4546:43]
    end else begin
      empty_26 <= Stack_26_io_empty; // @[stackmanage_35.scala 4585:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4547:43]
      empty_27 <= 1'h0; // @[stackmanage_35.scala 4547:43]
    end else begin
      empty_27 <= Stack_27_io_empty; // @[stackmanage_35.scala 4586:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4548:43]
      empty_28 <= 1'h0; // @[stackmanage_35.scala 4548:43]
    end else begin
      empty_28 <= Stack_28_io_empty; // @[stackmanage_35.scala 4587:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4549:43]
      empty_29 <= 1'h0; // @[stackmanage_35.scala 4549:43]
    end else begin
      empty_29 <= Stack_29_io_empty; // @[stackmanage_35.scala 4588:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4551:43]
      empty_30 <= 1'h0; // @[stackmanage_35.scala 4551:43]
    end else begin
      empty_30 <= Stack_30_io_empty; // @[stackmanage_35.scala 4590:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4552:43]
      empty_31 <= 1'h0; // @[stackmanage_35.scala 4552:43]
    end else begin
      empty_31 <= Stack_31_io_empty; // @[stackmanage_35.scala 4591:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4553:43]
      empty_32 <= 1'h0; // @[stackmanage_35.scala 4553:43]
    end else begin
      empty_32 <= Stack_32_io_empty; // @[stackmanage_35.scala 4592:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4554:43]
      empty_33 <= 1'h0; // @[stackmanage_35.scala 4554:43]
    end else begin
      empty_33 <= Stack_33_io_empty; // @[stackmanage_35.scala 4593:36]
    end
    if (reset) begin // @[stackmanage_35.scala 4555:43]
      empty_34 <= 1'h0; // @[stackmanage_35.scala 4555:43]
    end else begin
      empty_34 <= Stack_34_io_empty; // @[stackmanage_35.scala 4594:36]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  node_push_in_1 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  node_push_in_2 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  hitT_out_temp = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  ray_out_temp = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  node_out_temp = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  pop_valid_1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  pop_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  pop_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  pop_2 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  pop_3 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  pop_4 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  pop_5 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  pop_6 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  pop_7 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  pop_8 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  pop_9 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  pop_10 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  pop_11 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  pop_12 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  pop_13 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  pop_14 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  pop_15 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  pop_16 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  pop_17 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  pop_18 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  pop_19 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  pop_20 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  pop_21 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  pop_22 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  pop_23 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  pop_24 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  pop_25 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  pop_26 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  pop_27 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  pop_28 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  pop_29 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  pop_30 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  pop_31 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  pop_32 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  pop_33 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  pop_34 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  dispatch_0 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  dispatch_1 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  dispatch_2 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  dispatch_3 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  dispatch_4 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  dispatch_5 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  dispatch_6 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  dispatch_7 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  dispatch_8 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  dispatch_9 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  dispatch_10 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  dispatch_11 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  dispatch_12 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  dispatch_13 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  dispatch_14 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  dispatch_15 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  dispatch_16 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  dispatch_17 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  dispatch_18 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  dispatch_19 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  dispatch_20 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  dispatch_21 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  dispatch_22 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  dispatch_23 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  dispatch_24 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  dispatch_25 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  dispatch_26 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  dispatch_27 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  dispatch_28 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  dispatch_29 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  dispatch_30 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  dispatch_31 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  dispatch_32 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  dispatch_33 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  dispatch_34 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  dispatch_no_match = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  empty_0 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  empty_1 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  empty_2 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  empty_3 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  empty_4 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  empty_5 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  empty_6 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  empty_7 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  empty_8 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  empty_9 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  empty_10 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  empty_11 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  empty_12 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  empty_13 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  empty_14 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  empty_15 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  empty_16 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  empty_17 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  empty_18 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  empty_19 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  empty_20 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  empty_21 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  empty_22 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  empty_23 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  empty_24 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  empty_25 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  empty_26 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  empty_27 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  empty_28 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  empty_29 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  empty_30 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  empty_31 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  empty_32 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  empty_33 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  empty_34 = _RAND_111[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MY_MUL(
  input         clock,
  input         reset,
  input  [31:0] io_a,
  input  [31:0] io_b,
  output [31:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_REG_INIT
  wire [32:0] mulAddRecFNToRaw_preMul_io_a; // @[FMUL_1.scala 36:15]
  wire [32:0] mulAddRecFNToRaw_preMul_io_b; // @[FMUL_1.scala 36:15]
  wire [32:0] mulAddRecFNToRaw_preMul_io_c; // @[FMUL_1.scala 36:15]
  wire [23:0] mulAddRecFNToRaw_preMul_io_mulAddA; // @[FMUL_1.scala 36:15]
  wire [23:0] mulAddRecFNToRaw_preMul_io_mulAddB; // @[FMUL_1.scala 36:15]
  wire [47:0] mulAddRecFNToRaw_preMul_io_mulAddC; // @[FMUL_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny; // @[FMUL_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB; // @[FMUL_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfA; // @[FMUL_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA; // @[FMUL_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfB; // @[FMUL_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB; // @[FMUL_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_signProd; // @[FMUL_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC; // @[FMUL_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfC; // @[FMUL_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC; // @[FMUL_1.scala 36:15]
  wire [9:0] mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum; // @[FMUL_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags; // @[FMUL_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant; // @[FMUL_1.scala 36:15]
  wire [4:0] mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist; // @[FMUL_1.scala 36:15]
  wire [25:0] mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC; // @[FMUL_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC; // @[FMUL_1.scala 36:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny; // @[FMUL_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB; // @[FMUL_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA; // @[FMUL_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA; // @[FMUL_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB; // @[FMUL_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB; // @[FMUL_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_signProd; // @[FMUL_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC; // @[FMUL_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC; // @[FMUL_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC; // @[FMUL_1.scala 116:15]
  wire [9:0] mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum; // @[FMUL_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags; // @[FMUL_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant; // @[FMUL_1.scala 116:15]
  wire [4:0] mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist; // @[FMUL_1.scala 116:15]
  wire [25:0] mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC; // @[FMUL_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC; // @[FMUL_1.scala 116:15]
  wire [48:0] mulAddRecFNToRaw_postMul_io_mulAddResult; // @[FMUL_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_invalidExc; // @[FMUL_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isNaN; // @[FMUL_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isInf; // @[FMUL_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isZero; // @[FMUL_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_sign; // @[FMUL_1.scala 116:15]
  wire [9:0] mulAddRecFNToRaw_postMul_io_rawOut_sExp; // @[FMUL_1.scala 116:15]
  wire [26:0] mulAddRecFNToRaw_postMul_io_rawOut_sig; // @[FMUL_1.scala 116:15]
  wire  roundRawFNToRecFN_io_invalidExc; // @[FMUL_1.scala 137:15]
  wire  roundRawFNToRecFN_io_in_isNaN; // @[FMUL_1.scala 137:15]
  wire  roundRawFNToRecFN_io_in_isInf; // @[FMUL_1.scala 137:15]
  wire  roundRawFNToRecFN_io_in_isZero; // @[FMUL_1.scala 137:15]
  wire  roundRawFNToRecFN_io_in_sign; // @[FMUL_1.scala 137:15]
  wire [9:0] roundRawFNToRecFN_io_in_sExp; // @[FMUL_1.scala 137:15]
  wire [26:0] roundRawFNToRecFN_io_in_sig; // @[FMUL_1.scala 137:15]
  wire [32:0] roundRawFNToRecFN_io_out; // @[FMUL_1.scala 137:15]
  reg [23:0] premul_a; // @[FMUL_1.scala 15:37]
  reg [23:0] premul_b; // @[FMUL_1.scala 16:37]
  reg [47:0] premul_c; // @[FMUL_1.scala 17:37]
  reg  isSigNaNAny; // @[FMUL_1.scala 18:33]
  reg  isNaNAOrB; // @[FMUL_1.scala 19:34]
  reg  isInfA; // @[FMUL_1.scala 20:43]
  reg  isZeroA; // @[FMUL_1.scala 21:40]
  reg  isInfB; // @[FMUL_1.scala 22:43]
  reg  isZeroB; // @[FMUL_1.scala 23:40]
  reg  signProd; // @[FMUL_1.scala 24:38]
  reg  isNaNC; // @[FMUL_1.scala 25:39]
  reg  isInfC; // @[FMUL_1.scala 26:42]
  reg  isZeroC; // @[FMUL_1.scala 27:39]
  reg [9:0] sExpSum; // @[FMUL_1.scala 28:36]
  reg  doSubMags; // @[FMUL_1.scala 29:33]
  reg  CIsDominant; // @[FMUL_1.scala 30:33]
  reg [4:0] CDom_CAlignDist; // @[FMUL_1.scala 31:34]
  reg [25:0] highAlignedSigC; // @[FMUL_1.scala 32:37]
  reg  bit0AlignedSigC; // @[FMUL_1.scala 33:38]
  wire  _T_3 = io_a[30:23] == 8'h0; // @[rawFloatFromFN.scala 50:34]
  wire  _T_4 = io_a[22:0] == 23'h0; // @[rawFloatFromFN.scala 51:38]
  wire [4:0] _T_28 = io_a[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:69]
  wire [4:0] _T_29 = io_a[2] ? 5'h14 : _T_28; // @[Mux.scala 47:69]
  wire [4:0] _T_30 = io_a[3] ? 5'h13 : _T_29; // @[Mux.scala 47:69]
  wire [4:0] _T_31 = io_a[4] ? 5'h12 : _T_30; // @[Mux.scala 47:69]
  wire [4:0] _T_32 = io_a[5] ? 5'h11 : _T_31; // @[Mux.scala 47:69]
  wire [4:0] _T_33 = io_a[6] ? 5'h10 : _T_32; // @[Mux.scala 47:69]
  wire [4:0] _T_34 = io_a[7] ? 5'hf : _T_33; // @[Mux.scala 47:69]
  wire [4:0] _T_35 = io_a[8] ? 5'he : _T_34; // @[Mux.scala 47:69]
  wire [4:0] _T_36 = io_a[9] ? 5'hd : _T_35; // @[Mux.scala 47:69]
  wire [4:0] _T_37 = io_a[10] ? 5'hc : _T_36; // @[Mux.scala 47:69]
  wire [4:0] _T_38 = io_a[11] ? 5'hb : _T_37; // @[Mux.scala 47:69]
  wire [4:0] _T_39 = io_a[12] ? 5'ha : _T_38; // @[Mux.scala 47:69]
  wire [4:0] _T_40 = io_a[13] ? 5'h9 : _T_39; // @[Mux.scala 47:69]
  wire [4:0] _T_41 = io_a[14] ? 5'h8 : _T_40; // @[Mux.scala 47:69]
  wire [4:0] _T_42 = io_a[15] ? 5'h7 : _T_41; // @[Mux.scala 47:69]
  wire [4:0] _T_43 = io_a[16] ? 5'h6 : _T_42; // @[Mux.scala 47:69]
  wire [4:0] _T_44 = io_a[17] ? 5'h5 : _T_43; // @[Mux.scala 47:69]
  wire [4:0] _T_45 = io_a[18] ? 5'h4 : _T_44; // @[Mux.scala 47:69]
  wire [4:0] _T_46 = io_a[19] ? 5'h3 : _T_45; // @[Mux.scala 47:69]
  wire [4:0] _T_47 = io_a[20] ? 5'h2 : _T_46; // @[Mux.scala 47:69]
  wire [4:0] _T_48 = io_a[21] ? 5'h1 : _T_47; // @[Mux.scala 47:69]
  wire [4:0] _T_49 = io_a[22] ? 5'h0 : _T_48; // @[Mux.scala 47:69]
  wire [53:0] _GEN_0 = {{31'd0}, io_a[22:0]}; // @[rawFloatFromFN.scala 54:36]
  wire [53:0] _T_50 = _GEN_0 << _T_49; // @[rawFloatFromFN.scala 54:36]
  wire [22:0] _T_52 = {_T_50[21:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  wire [8:0] _GEN_1 = {{4'd0}, _T_49}; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_53 = _GEN_1 ^ 9'h1ff; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_54 = _T_3 ? _T_53 : {{1'd0}, io_a[30:23]}; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_55 = _T_3 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  wire [7:0] _GEN_2 = {{6'd0}, _T_55}; // @[rawFloatFromFN.scala 60:22]
  wire [7:0] _T_56 = 8'h80 | _GEN_2; // @[rawFloatFromFN.scala 60:22]
  wire [8:0] _GEN_3 = {{1'd0}, _T_56}; // @[rawFloatFromFN.scala 59:15]
  wire [8:0] _T_58 = _T_54 + _GEN_3; // @[rawFloatFromFN.scala 59:15]
  wire  _T_59 = _T_3 & _T_4; // @[rawFloatFromFN.scala 62:34]
  wire  _T_61 = _T_58[8:7] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  wire  _T_63 = _T_61 & ~_T_4; // @[rawFloatFromFN.scala 66:33]
  wire [9:0] _T_66 = {1'b0,$signed(_T_58)}; // @[rawFloatFromFN.scala 70:48]
  wire  hi_lo = ~_T_59; // @[rawFloatFromFN.scala 72:29]
  wire [22:0] lo = _T_3 ? _T_52 : io_a[22:0]; // @[rawFloatFromFN.scala 72:42]
  wire [24:0] _T_67 = {1'h0,hi_lo,lo}; // @[Cat.scala 30:58]
  wire [2:0] _T_69 = _T_59 ? 3'h0 : _T_66[8:6]; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_4 = {{2'd0}, _T_63}; // @[recFNFromFN.scala 48:79]
  wire [2:0] hi_lo_1 = _T_69 | _GEN_4; // @[recFNFromFN.scala 48:79]
  wire [5:0] lo_hi = _T_66[5:0]; // @[recFNFromFN.scala 50:23]
  wire [22:0] lo_lo = _T_67[22:0]; // @[recFNFromFN.scala 51:22]
  wire [28:0] lo_1 = {lo_hi,lo_lo}; // @[Cat.scala 30:58]
  wire [3:0] hi_1 = {io_a[31],hi_lo_1}; // @[Cat.scala 30:58]
  wire  _T_75 = io_b[30:23] == 8'h0; // @[rawFloatFromFN.scala 50:34]
  wire  _T_76 = io_b[22:0] == 23'h0; // @[rawFloatFromFN.scala 51:38]
  wire [4:0] _T_100 = io_b[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:69]
  wire [4:0] _T_101 = io_b[2] ? 5'h14 : _T_100; // @[Mux.scala 47:69]
  wire [4:0] _T_102 = io_b[3] ? 5'h13 : _T_101; // @[Mux.scala 47:69]
  wire [4:0] _T_103 = io_b[4] ? 5'h12 : _T_102; // @[Mux.scala 47:69]
  wire [4:0] _T_104 = io_b[5] ? 5'h11 : _T_103; // @[Mux.scala 47:69]
  wire [4:0] _T_105 = io_b[6] ? 5'h10 : _T_104; // @[Mux.scala 47:69]
  wire [4:0] _T_106 = io_b[7] ? 5'hf : _T_105; // @[Mux.scala 47:69]
  wire [4:0] _T_107 = io_b[8] ? 5'he : _T_106; // @[Mux.scala 47:69]
  wire [4:0] _T_108 = io_b[9] ? 5'hd : _T_107; // @[Mux.scala 47:69]
  wire [4:0] _T_109 = io_b[10] ? 5'hc : _T_108; // @[Mux.scala 47:69]
  wire [4:0] _T_110 = io_b[11] ? 5'hb : _T_109; // @[Mux.scala 47:69]
  wire [4:0] _T_111 = io_b[12] ? 5'ha : _T_110; // @[Mux.scala 47:69]
  wire [4:0] _T_112 = io_b[13] ? 5'h9 : _T_111; // @[Mux.scala 47:69]
  wire [4:0] _T_113 = io_b[14] ? 5'h8 : _T_112; // @[Mux.scala 47:69]
  wire [4:0] _T_114 = io_b[15] ? 5'h7 : _T_113; // @[Mux.scala 47:69]
  wire [4:0] _T_115 = io_b[16] ? 5'h6 : _T_114; // @[Mux.scala 47:69]
  wire [4:0] _T_116 = io_b[17] ? 5'h5 : _T_115; // @[Mux.scala 47:69]
  wire [4:0] _T_117 = io_b[18] ? 5'h4 : _T_116; // @[Mux.scala 47:69]
  wire [4:0] _T_118 = io_b[19] ? 5'h3 : _T_117; // @[Mux.scala 47:69]
  wire [4:0] _T_119 = io_b[20] ? 5'h2 : _T_118; // @[Mux.scala 47:69]
  wire [4:0] _T_120 = io_b[21] ? 5'h1 : _T_119; // @[Mux.scala 47:69]
  wire [4:0] _T_121 = io_b[22] ? 5'h0 : _T_120; // @[Mux.scala 47:69]
  wire [53:0] _GEN_5 = {{31'd0}, io_b[22:0]}; // @[rawFloatFromFN.scala 54:36]
  wire [53:0] _T_122 = _GEN_5 << _T_121; // @[rawFloatFromFN.scala 54:36]
  wire [22:0] _T_124 = {_T_122[21:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  wire [8:0] _GEN_6 = {{4'd0}, _T_121}; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_125 = _GEN_6 ^ 9'h1ff; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_126 = _T_75 ? _T_125 : {{1'd0}, io_b[30:23]}; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_127 = _T_75 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  wire [7:0] _GEN_7 = {{6'd0}, _T_127}; // @[rawFloatFromFN.scala 60:22]
  wire [7:0] _T_128 = 8'h80 | _GEN_7; // @[rawFloatFromFN.scala 60:22]
  wire [8:0] _GEN_8 = {{1'd0}, _T_128}; // @[rawFloatFromFN.scala 59:15]
  wire [8:0] _T_130 = _T_126 + _GEN_8; // @[rawFloatFromFN.scala 59:15]
  wire  _T_131 = _T_75 & _T_76; // @[rawFloatFromFN.scala 62:34]
  wire  _T_133 = _T_130[8:7] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  wire  _T_135 = _T_133 & ~_T_76; // @[rawFloatFromFN.scala 66:33]
  wire [9:0] _T_138 = {1'b0,$signed(_T_130)}; // @[rawFloatFromFN.scala 70:48]
  wire  hi_lo_2 = ~_T_131; // @[rawFloatFromFN.scala 72:29]
  wire [22:0] lo_2 = _T_75 ? _T_124 : io_b[22:0]; // @[rawFloatFromFN.scala 72:42]
  wire [24:0] _T_139 = {1'h0,hi_lo_2,lo_2}; // @[Cat.scala 30:58]
  wire [2:0] _T_141 = _T_131 ? 3'h0 : _T_138[8:6]; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_9 = {{2'd0}, _T_135}; // @[recFNFromFN.scala 48:79]
  wire [2:0] hi_lo_3 = _T_141 | _GEN_9; // @[recFNFromFN.scala 48:79]
  wire [5:0] lo_hi_1 = _T_138[5:0]; // @[recFNFromFN.scala 50:23]
  wire [22:0] lo_lo_1 = _T_139[22:0]; // @[recFNFromFN.scala 51:22]
  wire [28:0] lo_3 = {lo_hi_1,lo_lo_1}; // @[Cat.scala 30:58]
  wire [3:0] hi_3 = {io_b[31],hi_lo_3}; // @[Cat.scala 30:58]
  wire [31:0] _T_144 = io_a ^ io_b; // @[FMUL_1.scala 41:45]
  wire [31:0] _T_145 = _T_144 & 32'h80000000; // @[FMUL_1.scala 41:53]
  wire [47:0] _T_147 = premul_a * premul_b; // @[FMUL_1.scala 113:19]
  wire  _T_150 = roundRawFNToRecFN_io_out[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_152 = roundRawFNToRecFN_io_out[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  wire  _T_154 = _T_152 & roundRawFNToRecFN_io_out[29]; // @[rawFloatFromRecFN.scala 55:33]
  wire  _T_157 = _T_152 & ~roundRawFNToRecFN_io_out[29]; // @[rawFloatFromRecFN.scala 56:33]
  wire [9:0] _T_159 = {1'b0,$signed(roundRawFNToRecFN_io_out[31:23])}; // @[rawFloatFromRecFN.scala 59:27]
  wire  hi_lo_4 = ~_T_150; // @[rawFloatFromRecFN.scala 60:39]
  wire [22:0] lo_4 = roundRawFNToRecFN_io_out[22:0]; // @[rawFloatFromRecFN.scala 60:51]
  wire [24:0] _T_160 = {1'h0,hi_lo_4,lo_4}; // @[Cat.scala 30:58]
  wire  _T_161 = $signed(_T_159) < 10'sh82; // @[fNFromRecFN.scala 50:39]
  wire [4:0] _T_164 = 5'h1 - _T_159[4:0]; // @[fNFromRecFN.scala 51:39]
  wire [23:0] _T_166 = _T_160[24:1] >> _T_164; // @[fNFromRecFN.scala 52:42]
  wire [7:0] _T_170 = _T_159[7:0] - 8'h81; // @[fNFromRecFN.scala 57:45]
  wire [7:0] _T_171 = _T_161 ? 8'h0 : _T_170; // @[fNFromRecFN.scala 55:16]
  wire  _T_172 = _T_154 | _T_157; // @[fNFromRecFN.scala 59:44]
  wire [7:0] _T_174 = _T_172 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] hi_lo_5 = _T_171 | _T_174; // @[fNFromRecFN.scala 59:15]
  wire [22:0] _T_176 = _T_157 ? 23'h0 : _T_160[22:0]; // @[fNFromRecFN.scala 63:20]
  wire [22:0] lo_5 = _T_161 ? _T_166[22:0] : _T_176; // @[fNFromRecFN.scala 61:16]
  wire [8:0] hi_5 = {roundRawFNToRecFN_io_out[32],hi_lo_5}; // @[Cat.scala 30:58]
  MulAddRecFNToRaw_preMul mulAddRecFNToRaw_preMul ( // @[FMUL_1.scala 36:15]
    .io_a(mulAddRecFNToRaw_preMul_io_a),
    .io_b(mulAddRecFNToRaw_preMul_io_b),
    .io_c(mulAddRecFNToRaw_preMul_io_c),
    .io_mulAddA(mulAddRecFNToRaw_preMul_io_mulAddA),
    .io_mulAddB(mulAddRecFNToRaw_preMul_io_mulAddB),
    .io_mulAddC(mulAddRecFNToRaw_preMul_io_mulAddC),
    .io_toPostMul_isSigNaNAny(mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny),
    .io_toPostMul_isNaNAOrB(mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB),
    .io_toPostMul_isInfA(mulAddRecFNToRaw_preMul_io_toPostMul_isInfA),
    .io_toPostMul_isZeroA(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA),
    .io_toPostMul_isInfB(mulAddRecFNToRaw_preMul_io_toPostMul_isInfB),
    .io_toPostMul_isZeroB(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB),
    .io_toPostMul_signProd(mulAddRecFNToRaw_preMul_io_toPostMul_signProd),
    .io_toPostMul_isNaNC(mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC),
    .io_toPostMul_isInfC(mulAddRecFNToRaw_preMul_io_toPostMul_isInfC),
    .io_toPostMul_isZeroC(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC),
    .io_toPostMul_sExpSum(mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum),
    .io_toPostMul_doSubMags(mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags),
    .io_toPostMul_CIsDominant(mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant),
    .io_toPostMul_CDom_CAlignDist(mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist),
    .io_toPostMul_highAlignedSigC(mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC),
    .io_toPostMul_bit0AlignedSigC(mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC)
  );
  MulAddRecFNToRaw_postMul mulAddRecFNToRaw_postMul ( // @[FMUL_1.scala 116:15]
    .io_fromPreMul_isSigNaNAny(mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny),
    .io_fromPreMul_isNaNAOrB(mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB),
    .io_fromPreMul_isInfA(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA),
    .io_fromPreMul_isZeroA(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA),
    .io_fromPreMul_isInfB(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB),
    .io_fromPreMul_isZeroB(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB),
    .io_fromPreMul_signProd(mulAddRecFNToRaw_postMul_io_fromPreMul_signProd),
    .io_fromPreMul_isNaNC(mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC),
    .io_fromPreMul_isInfC(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC),
    .io_fromPreMul_isZeroC(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC),
    .io_fromPreMul_sExpSum(mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum),
    .io_fromPreMul_doSubMags(mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags),
    .io_fromPreMul_CIsDominant(mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant),
    .io_fromPreMul_CDom_CAlignDist(mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist),
    .io_fromPreMul_highAlignedSigC(mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC),
    .io_fromPreMul_bit0AlignedSigC(mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC),
    .io_mulAddResult(mulAddRecFNToRaw_postMul_io_mulAddResult),
    .io_invalidExc(mulAddRecFNToRaw_postMul_io_invalidExc),
    .io_rawOut_isNaN(mulAddRecFNToRaw_postMul_io_rawOut_isNaN),
    .io_rawOut_isInf(mulAddRecFNToRaw_postMul_io_rawOut_isInf),
    .io_rawOut_isZero(mulAddRecFNToRaw_postMul_io_rawOut_isZero),
    .io_rawOut_sign(mulAddRecFNToRaw_postMul_io_rawOut_sign),
    .io_rawOut_sExp(mulAddRecFNToRaw_postMul_io_rawOut_sExp),
    .io_rawOut_sig(mulAddRecFNToRaw_postMul_io_rawOut_sig)
  );
  RoundRawFNToRecFN roundRawFNToRecFN ( // @[FMUL_1.scala 137:15]
    .io_invalidExc(roundRawFNToRecFN_io_invalidExc),
    .io_in_isNaN(roundRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundRawFNToRecFN_io_in_sig),
    .io_out(roundRawFNToRecFN_io_out)
  );
  assign io_out = {hi_5,lo_5}; // @[Cat.scala 30:58]
  assign mulAddRecFNToRaw_preMul_io_a = {hi_1,lo_1}; // @[Cat.scala 30:58]
  assign mulAddRecFNToRaw_preMul_io_b = {hi_3,lo_3}; // @[Cat.scala 30:58]
  assign mulAddRecFNToRaw_preMul_io_c = {_T_145, 1'h0}; // @[FMUL_1.scala 41:75]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny = isSigNaNAny; // @[FMUL_1.scala 119:84]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB = isNaNAOrB; // @[FMUL_1.scala 120:86]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA = isInfA; // @[FMUL_1.scala 121:94]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA = isZeroA; // @[FMUL_1.scala 122:91]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB = isInfB; // @[FMUL_1.scala 123:94]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB = isZeroB; // @[FMUL_1.scala 124:91]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_signProd = signProd; // @[FMUL_1.scala 125:89]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC = isNaNC; // @[FMUL_1.scala 126:90]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC = isInfC; // @[FMUL_1.scala 127:94]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC = isZeroC; // @[FMUL_1.scala 128:91]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum = sExpSum; // @[FMUL_1.scala 129:88]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags = doSubMags; // @[FMUL_1.scala 130:85]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant = CIsDominant; // @[FMUL_1.scala 131:84]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist = CDom_CAlignDist; // @[FMUL_1.scala 132:78]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC = highAlignedSigC; // @[FMUL_1.scala 133:80]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC = bit0AlignedSigC; // @[FMUL_1.scala 134:82]
  assign mulAddRecFNToRaw_postMul_io_mulAddResult = _T_147 + premul_c; // @[FMUL_1.scala 113:31]
  assign roundRawFNToRecFN_io_invalidExc = mulAddRecFNToRaw_postMul_io_invalidExc; // @[FMUL_1.scala 138:39]
  assign roundRawFNToRecFN_io_in_isNaN = mulAddRecFNToRaw_postMul_io_rawOut_isNaN; // @[FMUL_1.scala 140:39]
  assign roundRawFNToRecFN_io_in_isInf = mulAddRecFNToRaw_postMul_io_rawOut_isInf; // @[FMUL_1.scala 140:39]
  assign roundRawFNToRecFN_io_in_isZero = mulAddRecFNToRaw_postMul_io_rawOut_isZero; // @[FMUL_1.scala 140:39]
  assign roundRawFNToRecFN_io_in_sign = mulAddRecFNToRaw_postMul_io_rawOut_sign; // @[FMUL_1.scala 140:39]
  assign roundRawFNToRecFN_io_in_sExp = mulAddRecFNToRaw_postMul_io_rawOut_sExp; // @[FMUL_1.scala 140:39]
  assign roundRawFNToRecFN_io_in_sig = mulAddRecFNToRaw_postMul_io_rawOut_sig; // @[FMUL_1.scala 140:39]
  always @(posedge clock) begin
    if (reset) begin // @[FMUL_1.scala 15:37]
      premul_a <= 24'h0; // @[FMUL_1.scala 15:37]
    end else begin
      premul_a <= mulAddRecFNToRaw_preMul_io_mulAddA; // @[FMUL_1.scala 103:63]
    end
    if (reset) begin // @[FMUL_1.scala 16:37]
      premul_b <= 24'h0; // @[FMUL_1.scala 16:37]
    end else begin
      premul_b <= mulAddRecFNToRaw_preMul_io_mulAddB; // @[FMUL_1.scala 104:63]
    end
    if (reset) begin // @[FMUL_1.scala 17:37]
      premul_c <= 48'h0; // @[FMUL_1.scala 17:37]
    end else begin
      premul_c <= mulAddRecFNToRaw_preMul_io_mulAddC; // @[FMUL_1.scala 105:63]
    end
    if (reset) begin // @[FMUL_1.scala 18:33]
      isSigNaNAny <= 1'h0; // @[FMUL_1.scala 18:33]
    end else begin
      isSigNaNAny <= mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny; // @[FMUL_1.scala 43:61]
    end
    if (reset) begin // @[FMUL_1.scala 19:34]
      isNaNAOrB <= 1'h0; // @[FMUL_1.scala 19:34]
    end else begin
      isNaNAOrB <= mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB; // @[FMUL_1.scala 44:62]
    end
    if (reset) begin // @[FMUL_1.scala 20:43]
      isInfA <= 1'h0; // @[FMUL_1.scala 20:43]
    end else begin
      isInfA <= mulAddRecFNToRaw_preMul_io_toPostMul_isInfA; // @[FMUL_1.scala 45:70]
    end
    if (reset) begin // @[FMUL_1.scala 21:40]
      isZeroA <= 1'h0; // @[FMUL_1.scala 21:40]
    end else begin
      isZeroA <= mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA; // @[FMUL_1.scala 46:67]
    end
    if (reset) begin // @[FMUL_1.scala 22:43]
      isInfB <= 1'h0; // @[FMUL_1.scala 22:43]
    end else begin
      isInfB <= mulAddRecFNToRaw_preMul_io_toPostMul_isInfB; // @[FMUL_1.scala 47:70]
    end
    if (reset) begin // @[FMUL_1.scala 23:40]
      isZeroB <= 1'h0; // @[FMUL_1.scala 23:40]
    end else begin
      isZeroB <= mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB; // @[FMUL_1.scala 48:67]
    end
    if (reset) begin // @[FMUL_1.scala 24:38]
      signProd <= 1'h0; // @[FMUL_1.scala 24:38]
    end else begin
      signProd <= mulAddRecFNToRaw_preMul_io_toPostMul_signProd; // @[FMUL_1.scala 49:65]
    end
    if (reset) begin // @[FMUL_1.scala 25:39]
      isNaNC <= 1'h0; // @[FMUL_1.scala 25:39]
    end else begin
      isNaNC <= mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC; // @[FMUL_1.scala 50:66]
    end
    if (reset) begin // @[FMUL_1.scala 26:42]
      isInfC <= 1'h0; // @[FMUL_1.scala 26:42]
    end else begin
      isInfC <= mulAddRecFNToRaw_preMul_io_toPostMul_isInfC; // @[FMUL_1.scala 51:69]
    end
    if (reset) begin // @[FMUL_1.scala 27:39]
      isZeroC <= 1'h0; // @[FMUL_1.scala 27:39]
    end else begin
      isZeroC <= mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC; // @[FMUL_1.scala 52:66]
    end
    if (reset) begin // @[FMUL_1.scala 28:36]
      sExpSum <= 10'sh0; // @[FMUL_1.scala 28:36]
    end else begin
      sExpSum <= mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum; // @[FMUL_1.scala 53:63]
    end
    if (reset) begin // @[FMUL_1.scala 29:33]
      doSubMags <= 1'h0; // @[FMUL_1.scala 29:33]
    end else begin
      doSubMags <= mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags; // @[FMUL_1.scala 54:60]
    end
    if (reset) begin // @[FMUL_1.scala 30:33]
      CIsDominant <= 1'h0; // @[FMUL_1.scala 30:33]
    end else begin
      CIsDominant <= mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant; // @[FMUL_1.scala 55:59]
    end
    if (reset) begin // @[FMUL_1.scala 31:34]
      CDom_CAlignDist <= 5'h0; // @[FMUL_1.scala 31:34]
    end else begin
      CDom_CAlignDist <= mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist; // @[FMUL_1.scala 56:54]
    end
    if (reset) begin // @[FMUL_1.scala 32:37]
      highAlignedSigC <= 26'h0; // @[FMUL_1.scala 32:37]
    end else begin
      highAlignedSigC <= mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC; // @[FMUL_1.scala 57:56]
    end
    if (reset) begin // @[FMUL_1.scala 33:38]
      bit0AlignedSigC <= 1'h0; // @[FMUL_1.scala 33:38]
    end else begin
      bit0AlignedSigC <= mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC; // @[FMUL_1.scala 58:57]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  premul_a = _RAND_0[23:0];
  _RAND_1 = {1{`RANDOM}};
  premul_b = _RAND_1[23:0];
  _RAND_2 = {2{`RANDOM}};
  premul_c = _RAND_2[47:0];
  _RAND_3 = {1{`RANDOM}};
  isSigNaNAny = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  isNaNAOrB = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  isInfA = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  isZeroA = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  isInfB = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  isZeroB = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  signProd = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  isNaNC = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  isInfC = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  isZeroC = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  sExpSum = _RAND_13[9:0];
  _RAND_14 = {1{`RANDOM}};
  doSubMags = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  CIsDominant = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  CDom_CAlignDist = _RAND_16[4:0];
  _RAND_17 = {1{`RANDOM}};
  highAlignedSigC = _RAND_17[25:0];
  _RAND_18 = {1{`RANDOM}};
  bit0AlignedSigC = _RAND_18[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MY_ADD(
  input         clock,
  input         reset,
  input  [31:0] io_a,
  input  [31:0] io_b,
  output [31:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_REG_INIT
  wire [32:0] mulAddRecFNToRaw_preMul_io_a; // @[FADD_1.scala 36:15]
  wire [32:0] mulAddRecFNToRaw_preMul_io_b; // @[FADD_1.scala 36:15]
  wire [32:0] mulAddRecFNToRaw_preMul_io_c; // @[FADD_1.scala 36:15]
  wire [23:0] mulAddRecFNToRaw_preMul_io_mulAddA; // @[FADD_1.scala 36:15]
  wire [23:0] mulAddRecFNToRaw_preMul_io_mulAddB; // @[FADD_1.scala 36:15]
  wire [47:0] mulAddRecFNToRaw_preMul_io_mulAddC; // @[FADD_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny; // @[FADD_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB; // @[FADD_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfA; // @[FADD_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA; // @[FADD_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfB; // @[FADD_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB; // @[FADD_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_signProd; // @[FADD_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC; // @[FADD_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfC; // @[FADD_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC; // @[FADD_1.scala 36:15]
  wire [9:0] mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum; // @[FADD_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags; // @[FADD_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant; // @[FADD_1.scala 36:15]
  wire [4:0] mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist; // @[FADD_1.scala 36:15]
  wire [25:0] mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC; // @[FADD_1.scala 36:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC; // @[FADD_1.scala 36:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny; // @[FADD_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB; // @[FADD_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA; // @[FADD_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA; // @[FADD_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB; // @[FADD_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB; // @[FADD_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_signProd; // @[FADD_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC; // @[FADD_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC; // @[FADD_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC; // @[FADD_1.scala 116:15]
  wire [9:0] mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum; // @[FADD_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags; // @[FADD_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant; // @[FADD_1.scala 116:15]
  wire [4:0] mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist; // @[FADD_1.scala 116:15]
  wire [25:0] mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC; // @[FADD_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC; // @[FADD_1.scala 116:15]
  wire [48:0] mulAddRecFNToRaw_postMul_io_mulAddResult; // @[FADD_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_invalidExc; // @[FADD_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isNaN; // @[FADD_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isInf; // @[FADD_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isZero; // @[FADD_1.scala 116:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_sign; // @[FADD_1.scala 116:15]
  wire [9:0] mulAddRecFNToRaw_postMul_io_rawOut_sExp; // @[FADD_1.scala 116:15]
  wire [26:0] mulAddRecFNToRaw_postMul_io_rawOut_sig; // @[FADD_1.scala 116:15]
  wire  roundRawFNToRecFN_io_invalidExc; // @[FADD_1.scala 137:15]
  wire  roundRawFNToRecFN_io_in_isNaN; // @[FADD_1.scala 137:15]
  wire  roundRawFNToRecFN_io_in_isInf; // @[FADD_1.scala 137:15]
  wire  roundRawFNToRecFN_io_in_isZero; // @[FADD_1.scala 137:15]
  wire  roundRawFNToRecFN_io_in_sign; // @[FADD_1.scala 137:15]
  wire [9:0] roundRawFNToRecFN_io_in_sExp; // @[FADD_1.scala 137:15]
  wire [26:0] roundRawFNToRecFN_io_in_sig; // @[FADD_1.scala 137:15]
  wire [32:0] roundRawFNToRecFN_io_out; // @[FADD_1.scala 137:15]
  reg [23:0] premul_a; // @[FADD_1.scala 15:37]
  reg [23:0] premul_b; // @[FADD_1.scala 16:37]
  reg [47:0] premul_c; // @[FADD_1.scala 17:37]
  reg  isSigNaNAny; // @[FADD_1.scala 18:33]
  reg  isNaNAOrB; // @[FADD_1.scala 19:34]
  reg  isInfA; // @[FADD_1.scala 20:43]
  reg  isZeroA; // @[FADD_1.scala 21:40]
  reg  isInfB; // @[FADD_1.scala 22:43]
  reg  isZeroB; // @[FADD_1.scala 23:40]
  reg  signProd; // @[FADD_1.scala 24:38]
  reg  isNaNC; // @[FADD_1.scala 25:39]
  reg  isInfC; // @[FADD_1.scala 26:42]
  reg  isZeroC; // @[FADD_1.scala 27:39]
  reg [9:0] sExpSum; // @[FADD_1.scala 28:36]
  reg  doSubMags; // @[FADD_1.scala 29:33]
  reg  CIsDominant; // @[FADD_1.scala 30:33]
  reg [4:0] CDom_CAlignDist; // @[FADD_1.scala 31:34]
  reg [25:0] highAlignedSigC; // @[FADD_1.scala 32:37]
  reg  bit0AlignedSigC; // @[FADD_1.scala 33:38]
  wire  _T_3 = io_a[30:23] == 8'h0; // @[rawFloatFromFN.scala 50:34]
  wire  _T_4 = io_a[22:0] == 23'h0; // @[rawFloatFromFN.scala 51:38]
  wire [4:0] _T_28 = io_a[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:69]
  wire [4:0] _T_29 = io_a[2] ? 5'h14 : _T_28; // @[Mux.scala 47:69]
  wire [4:0] _T_30 = io_a[3] ? 5'h13 : _T_29; // @[Mux.scala 47:69]
  wire [4:0] _T_31 = io_a[4] ? 5'h12 : _T_30; // @[Mux.scala 47:69]
  wire [4:0] _T_32 = io_a[5] ? 5'h11 : _T_31; // @[Mux.scala 47:69]
  wire [4:0] _T_33 = io_a[6] ? 5'h10 : _T_32; // @[Mux.scala 47:69]
  wire [4:0] _T_34 = io_a[7] ? 5'hf : _T_33; // @[Mux.scala 47:69]
  wire [4:0] _T_35 = io_a[8] ? 5'he : _T_34; // @[Mux.scala 47:69]
  wire [4:0] _T_36 = io_a[9] ? 5'hd : _T_35; // @[Mux.scala 47:69]
  wire [4:0] _T_37 = io_a[10] ? 5'hc : _T_36; // @[Mux.scala 47:69]
  wire [4:0] _T_38 = io_a[11] ? 5'hb : _T_37; // @[Mux.scala 47:69]
  wire [4:0] _T_39 = io_a[12] ? 5'ha : _T_38; // @[Mux.scala 47:69]
  wire [4:0] _T_40 = io_a[13] ? 5'h9 : _T_39; // @[Mux.scala 47:69]
  wire [4:0] _T_41 = io_a[14] ? 5'h8 : _T_40; // @[Mux.scala 47:69]
  wire [4:0] _T_42 = io_a[15] ? 5'h7 : _T_41; // @[Mux.scala 47:69]
  wire [4:0] _T_43 = io_a[16] ? 5'h6 : _T_42; // @[Mux.scala 47:69]
  wire [4:0] _T_44 = io_a[17] ? 5'h5 : _T_43; // @[Mux.scala 47:69]
  wire [4:0] _T_45 = io_a[18] ? 5'h4 : _T_44; // @[Mux.scala 47:69]
  wire [4:0] _T_46 = io_a[19] ? 5'h3 : _T_45; // @[Mux.scala 47:69]
  wire [4:0] _T_47 = io_a[20] ? 5'h2 : _T_46; // @[Mux.scala 47:69]
  wire [4:0] _T_48 = io_a[21] ? 5'h1 : _T_47; // @[Mux.scala 47:69]
  wire [4:0] _T_49 = io_a[22] ? 5'h0 : _T_48; // @[Mux.scala 47:69]
  wire [53:0] _GEN_0 = {{31'd0}, io_a[22:0]}; // @[rawFloatFromFN.scala 54:36]
  wire [53:0] _T_50 = _GEN_0 << _T_49; // @[rawFloatFromFN.scala 54:36]
  wire [22:0] _T_52 = {_T_50[21:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  wire [8:0] _GEN_1 = {{4'd0}, _T_49}; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_53 = _GEN_1 ^ 9'h1ff; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_54 = _T_3 ? _T_53 : {{1'd0}, io_a[30:23]}; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_55 = _T_3 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  wire [7:0] _GEN_2 = {{6'd0}, _T_55}; // @[rawFloatFromFN.scala 60:22]
  wire [7:0] _T_56 = 8'h80 | _GEN_2; // @[rawFloatFromFN.scala 60:22]
  wire [8:0] _GEN_3 = {{1'd0}, _T_56}; // @[rawFloatFromFN.scala 59:15]
  wire [8:0] _T_58 = _T_54 + _GEN_3; // @[rawFloatFromFN.scala 59:15]
  wire  _T_59 = _T_3 & _T_4; // @[rawFloatFromFN.scala 62:34]
  wire  _T_61 = _T_58[8:7] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  wire  _T_63 = _T_61 & ~_T_4; // @[rawFloatFromFN.scala 66:33]
  wire [9:0] _T_66 = {1'b0,$signed(_T_58)}; // @[rawFloatFromFN.scala 70:48]
  wire  hi_lo = ~_T_59; // @[rawFloatFromFN.scala 72:29]
  wire [22:0] lo = _T_3 ? _T_52 : io_a[22:0]; // @[rawFloatFromFN.scala 72:42]
  wire [24:0] _T_67 = {1'h0,hi_lo,lo}; // @[Cat.scala 30:58]
  wire [2:0] _T_69 = _T_59 ? 3'h0 : _T_66[8:6]; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_4 = {{2'd0}, _T_63}; // @[recFNFromFN.scala 48:79]
  wire [2:0] hi_lo_1 = _T_69 | _GEN_4; // @[recFNFromFN.scala 48:79]
  wire [5:0] lo_hi = _T_66[5:0]; // @[recFNFromFN.scala 50:23]
  wire [22:0] lo_lo = _T_67[22:0]; // @[recFNFromFN.scala 51:22]
  wire [28:0] lo_1 = {lo_hi,lo_lo}; // @[Cat.scala 30:58]
  wire [3:0] hi_1 = {io_a[31],hi_lo_1}; // @[Cat.scala 30:58]
  wire  _T_75 = io_b[30:23] == 8'h0; // @[rawFloatFromFN.scala 50:34]
  wire  _T_76 = io_b[22:0] == 23'h0; // @[rawFloatFromFN.scala 51:38]
  wire [4:0] _T_100 = io_b[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:69]
  wire [4:0] _T_101 = io_b[2] ? 5'h14 : _T_100; // @[Mux.scala 47:69]
  wire [4:0] _T_102 = io_b[3] ? 5'h13 : _T_101; // @[Mux.scala 47:69]
  wire [4:0] _T_103 = io_b[4] ? 5'h12 : _T_102; // @[Mux.scala 47:69]
  wire [4:0] _T_104 = io_b[5] ? 5'h11 : _T_103; // @[Mux.scala 47:69]
  wire [4:0] _T_105 = io_b[6] ? 5'h10 : _T_104; // @[Mux.scala 47:69]
  wire [4:0] _T_106 = io_b[7] ? 5'hf : _T_105; // @[Mux.scala 47:69]
  wire [4:0] _T_107 = io_b[8] ? 5'he : _T_106; // @[Mux.scala 47:69]
  wire [4:0] _T_108 = io_b[9] ? 5'hd : _T_107; // @[Mux.scala 47:69]
  wire [4:0] _T_109 = io_b[10] ? 5'hc : _T_108; // @[Mux.scala 47:69]
  wire [4:0] _T_110 = io_b[11] ? 5'hb : _T_109; // @[Mux.scala 47:69]
  wire [4:0] _T_111 = io_b[12] ? 5'ha : _T_110; // @[Mux.scala 47:69]
  wire [4:0] _T_112 = io_b[13] ? 5'h9 : _T_111; // @[Mux.scala 47:69]
  wire [4:0] _T_113 = io_b[14] ? 5'h8 : _T_112; // @[Mux.scala 47:69]
  wire [4:0] _T_114 = io_b[15] ? 5'h7 : _T_113; // @[Mux.scala 47:69]
  wire [4:0] _T_115 = io_b[16] ? 5'h6 : _T_114; // @[Mux.scala 47:69]
  wire [4:0] _T_116 = io_b[17] ? 5'h5 : _T_115; // @[Mux.scala 47:69]
  wire [4:0] _T_117 = io_b[18] ? 5'h4 : _T_116; // @[Mux.scala 47:69]
  wire [4:0] _T_118 = io_b[19] ? 5'h3 : _T_117; // @[Mux.scala 47:69]
  wire [4:0] _T_119 = io_b[20] ? 5'h2 : _T_118; // @[Mux.scala 47:69]
  wire [4:0] _T_120 = io_b[21] ? 5'h1 : _T_119; // @[Mux.scala 47:69]
  wire [4:0] _T_121 = io_b[22] ? 5'h0 : _T_120; // @[Mux.scala 47:69]
  wire [53:0] _GEN_5 = {{31'd0}, io_b[22:0]}; // @[rawFloatFromFN.scala 54:36]
  wire [53:0] _T_122 = _GEN_5 << _T_121; // @[rawFloatFromFN.scala 54:36]
  wire [22:0] _T_124 = {_T_122[21:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  wire [8:0] _GEN_6 = {{4'd0}, _T_121}; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_125 = _GEN_6 ^ 9'h1ff; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_126 = _T_75 ? _T_125 : {{1'd0}, io_b[30:23]}; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_127 = _T_75 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  wire [7:0] _GEN_7 = {{6'd0}, _T_127}; // @[rawFloatFromFN.scala 60:22]
  wire [7:0] _T_128 = 8'h80 | _GEN_7; // @[rawFloatFromFN.scala 60:22]
  wire [8:0] _GEN_8 = {{1'd0}, _T_128}; // @[rawFloatFromFN.scala 59:15]
  wire [8:0] _T_130 = _T_126 + _GEN_8; // @[rawFloatFromFN.scala 59:15]
  wire  _T_131 = _T_75 & _T_76; // @[rawFloatFromFN.scala 62:34]
  wire  _T_133 = _T_130[8:7] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  wire  _T_135 = _T_133 & ~_T_76; // @[rawFloatFromFN.scala 66:33]
  wire [9:0] _T_138 = {1'b0,$signed(_T_130)}; // @[rawFloatFromFN.scala 70:48]
  wire  hi_lo_2 = ~_T_131; // @[rawFloatFromFN.scala 72:29]
  wire [22:0] lo_2 = _T_75 ? _T_124 : io_b[22:0]; // @[rawFloatFromFN.scala 72:42]
  wire [24:0] _T_139 = {1'h0,hi_lo_2,lo_2}; // @[Cat.scala 30:58]
  wire [2:0] _T_141 = _T_131 ? 3'h0 : _T_138[8:6]; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_9 = {{2'd0}, _T_135}; // @[recFNFromFN.scala 48:79]
  wire [2:0] hi_lo_3 = _T_141 | _GEN_9; // @[recFNFromFN.scala 48:79]
  wire [5:0] lo_hi_1 = _T_138[5:0]; // @[recFNFromFN.scala 50:23]
  wire [22:0] lo_lo_1 = _T_139[22:0]; // @[recFNFromFN.scala 51:22]
  wire [28:0] lo_3 = {lo_hi_1,lo_lo_1}; // @[Cat.scala 30:58]
  wire [3:0] hi_3 = {io_b[31],hi_lo_3}; // @[Cat.scala 30:58]
  wire [47:0] _T_144 = premul_a * premul_b; // @[FADD_1.scala 113:19]
  wire  _T_147 = roundRawFNToRecFN_io_out[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_149 = roundRawFNToRecFN_io_out[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  wire  _T_151 = _T_149 & roundRawFNToRecFN_io_out[29]; // @[rawFloatFromRecFN.scala 55:33]
  wire  _T_154 = _T_149 & ~roundRawFNToRecFN_io_out[29]; // @[rawFloatFromRecFN.scala 56:33]
  wire [9:0] _T_156 = {1'b0,$signed(roundRawFNToRecFN_io_out[31:23])}; // @[rawFloatFromRecFN.scala 59:27]
  wire  hi_lo_4 = ~_T_147; // @[rawFloatFromRecFN.scala 60:39]
  wire [22:0] lo_4 = roundRawFNToRecFN_io_out[22:0]; // @[rawFloatFromRecFN.scala 60:51]
  wire [24:0] _T_157 = {1'h0,hi_lo_4,lo_4}; // @[Cat.scala 30:58]
  wire  _T_158 = $signed(_T_156) < 10'sh82; // @[fNFromRecFN.scala 50:39]
  wire [4:0] _T_161 = 5'h1 - _T_156[4:0]; // @[fNFromRecFN.scala 51:39]
  wire [23:0] _T_163 = _T_157[24:1] >> _T_161; // @[fNFromRecFN.scala 52:42]
  wire [7:0] _T_167 = _T_156[7:0] - 8'h81; // @[fNFromRecFN.scala 57:45]
  wire [7:0] _T_168 = _T_158 ? 8'h0 : _T_167; // @[fNFromRecFN.scala 55:16]
  wire  _T_169 = _T_151 | _T_154; // @[fNFromRecFN.scala 59:44]
  wire [7:0] _T_171 = _T_169 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] hi_lo_5 = _T_168 | _T_171; // @[fNFromRecFN.scala 59:15]
  wire [22:0] _T_173 = _T_154 ? 23'h0 : _T_157[22:0]; // @[fNFromRecFN.scala 63:20]
  wire [22:0] lo_5 = _T_158 ? _T_163[22:0] : _T_173; // @[fNFromRecFN.scala 61:16]
  wire [8:0] hi_5 = {roundRawFNToRecFN_io_out[32],hi_lo_5}; // @[Cat.scala 30:58]
  MulAddRecFNToRaw_preMul mulAddRecFNToRaw_preMul ( // @[FADD_1.scala 36:15]
    .io_a(mulAddRecFNToRaw_preMul_io_a),
    .io_b(mulAddRecFNToRaw_preMul_io_b),
    .io_c(mulAddRecFNToRaw_preMul_io_c),
    .io_mulAddA(mulAddRecFNToRaw_preMul_io_mulAddA),
    .io_mulAddB(mulAddRecFNToRaw_preMul_io_mulAddB),
    .io_mulAddC(mulAddRecFNToRaw_preMul_io_mulAddC),
    .io_toPostMul_isSigNaNAny(mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny),
    .io_toPostMul_isNaNAOrB(mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB),
    .io_toPostMul_isInfA(mulAddRecFNToRaw_preMul_io_toPostMul_isInfA),
    .io_toPostMul_isZeroA(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA),
    .io_toPostMul_isInfB(mulAddRecFNToRaw_preMul_io_toPostMul_isInfB),
    .io_toPostMul_isZeroB(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB),
    .io_toPostMul_signProd(mulAddRecFNToRaw_preMul_io_toPostMul_signProd),
    .io_toPostMul_isNaNC(mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC),
    .io_toPostMul_isInfC(mulAddRecFNToRaw_preMul_io_toPostMul_isInfC),
    .io_toPostMul_isZeroC(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC),
    .io_toPostMul_sExpSum(mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum),
    .io_toPostMul_doSubMags(mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags),
    .io_toPostMul_CIsDominant(mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant),
    .io_toPostMul_CDom_CAlignDist(mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist),
    .io_toPostMul_highAlignedSigC(mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC),
    .io_toPostMul_bit0AlignedSigC(mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC)
  );
  MulAddRecFNToRaw_postMul mulAddRecFNToRaw_postMul ( // @[FADD_1.scala 116:15]
    .io_fromPreMul_isSigNaNAny(mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny),
    .io_fromPreMul_isNaNAOrB(mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB),
    .io_fromPreMul_isInfA(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA),
    .io_fromPreMul_isZeroA(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA),
    .io_fromPreMul_isInfB(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB),
    .io_fromPreMul_isZeroB(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB),
    .io_fromPreMul_signProd(mulAddRecFNToRaw_postMul_io_fromPreMul_signProd),
    .io_fromPreMul_isNaNC(mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC),
    .io_fromPreMul_isInfC(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC),
    .io_fromPreMul_isZeroC(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC),
    .io_fromPreMul_sExpSum(mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum),
    .io_fromPreMul_doSubMags(mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags),
    .io_fromPreMul_CIsDominant(mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant),
    .io_fromPreMul_CDom_CAlignDist(mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist),
    .io_fromPreMul_highAlignedSigC(mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC),
    .io_fromPreMul_bit0AlignedSigC(mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC),
    .io_mulAddResult(mulAddRecFNToRaw_postMul_io_mulAddResult),
    .io_invalidExc(mulAddRecFNToRaw_postMul_io_invalidExc),
    .io_rawOut_isNaN(mulAddRecFNToRaw_postMul_io_rawOut_isNaN),
    .io_rawOut_isInf(mulAddRecFNToRaw_postMul_io_rawOut_isInf),
    .io_rawOut_isZero(mulAddRecFNToRaw_postMul_io_rawOut_isZero),
    .io_rawOut_sign(mulAddRecFNToRaw_postMul_io_rawOut_sign),
    .io_rawOut_sExp(mulAddRecFNToRaw_postMul_io_rawOut_sExp),
    .io_rawOut_sig(mulAddRecFNToRaw_postMul_io_rawOut_sig)
  );
  RoundRawFNToRecFN roundRawFNToRecFN ( // @[FADD_1.scala 137:15]
    .io_invalidExc(roundRawFNToRecFN_io_invalidExc),
    .io_in_isNaN(roundRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundRawFNToRecFN_io_in_sig),
    .io_out(roundRawFNToRecFN_io_out)
  );
  assign io_out = {hi_5,lo_5}; // @[Cat.scala 30:58]
  assign mulAddRecFNToRaw_preMul_io_a = {hi_1,lo_1}; // @[Cat.scala 30:58]
  assign mulAddRecFNToRaw_preMul_io_b = 33'h80000000; // @[FADD_1.scala 40:35]
  assign mulAddRecFNToRaw_preMul_io_c = {hi_3,lo_3}; // @[Cat.scala 30:58]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny = isSigNaNAny; // @[FADD_1.scala 119:84]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB = isNaNAOrB; // @[FADD_1.scala 120:86]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA = isInfA; // @[FADD_1.scala 121:94]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA = isZeroA; // @[FADD_1.scala 122:91]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB = isInfB; // @[FADD_1.scala 123:94]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB = isZeroB; // @[FADD_1.scala 124:91]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_signProd = signProd; // @[FADD_1.scala 125:89]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC = isNaNC; // @[FADD_1.scala 126:90]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC = isInfC; // @[FADD_1.scala 127:94]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC = isZeroC; // @[FADD_1.scala 128:91]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum = sExpSum; // @[FADD_1.scala 129:88]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags = doSubMags; // @[FADD_1.scala 130:85]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant = CIsDominant; // @[FADD_1.scala 131:84]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist = CDom_CAlignDist; // @[FADD_1.scala 132:78]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC = highAlignedSigC; // @[FADD_1.scala 133:80]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC = bit0AlignedSigC; // @[FADD_1.scala 134:82]
  assign mulAddRecFNToRaw_postMul_io_mulAddResult = _T_144 + premul_c; // @[FADD_1.scala 113:31]
  assign roundRawFNToRecFN_io_invalidExc = mulAddRecFNToRaw_postMul_io_invalidExc; // @[FADD_1.scala 138:39]
  assign roundRawFNToRecFN_io_in_isNaN = mulAddRecFNToRaw_postMul_io_rawOut_isNaN; // @[FADD_1.scala 140:39]
  assign roundRawFNToRecFN_io_in_isInf = mulAddRecFNToRaw_postMul_io_rawOut_isInf; // @[FADD_1.scala 140:39]
  assign roundRawFNToRecFN_io_in_isZero = mulAddRecFNToRaw_postMul_io_rawOut_isZero; // @[FADD_1.scala 140:39]
  assign roundRawFNToRecFN_io_in_sign = mulAddRecFNToRaw_postMul_io_rawOut_sign; // @[FADD_1.scala 140:39]
  assign roundRawFNToRecFN_io_in_sExp = mulAddRecFNToRaw_postMul_io_rawOut_sExp; // @[FADD_1.scala 140:39]
  assign roundRawFNToRecFN_io_in_sig = mulAddRecFNToRaw_postMul_io_rawOut_sig; // @[FADD_1.scala 140:39]
  always @(posedge clock) begin
    if (reset) begin // @[FADD_1.scala 15:37]
      premul_a <= 24'h0; // @[FADD_1.scala 15:37]
    end else begin
      premul_a <= mulAddRecFNToRaw_preMul_io_mulAddA; // @[FADD_1.scala 103:63]
    end
    if (reset) begin // @[FADD_1.scala 16:37]
      premul_b <= 24'h0; // @[FADD_1.scala 16:37]
    end else begin
      premul_b <= mulAddRecFNToRaw_preMul_io_mulAddB; // @[FADD_1.scala 104:63]
    end
    if (reset) begin // @[FADD_1.scala 17:37]
      premul_c <= 48'h0; // @[FADD_1.scala 17:37]
    end else begin
      premul_c <= mulAddRecFNToRaw_preMul_io_mulAddC; // @[FADD_1.scala 105:63]
    end
    if (reset) begin // @[FADD_1.scala 18:33]
      isSigNaNAny <= 1'h0; // @[FADD_1.scala 18:33]
    end else begin
      isSigNaNAny <= mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny; // @[FADD_1.scala 43:61]
    end
    if (reset) begin // @[FADD_1.scala 19:34]
      isNaNAOrB <= 1'h0; // @[FADD_1.scala 19:34]
    end else begin
      isNaNAOrB <= mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB; // @[FADD_1.scala 44:62]
    end
    if (reset) begin // @[FADD_1.scala 20:43]
      isInfA <= 1'h0; // @[FADD_1.scala 20:43]
    end else begin
      isInfA <= mulAddRecFNToRaw_preMul_io_toPostMul_isInfA; // @[FADD_1.scala 45:70]
    end
    if (reset) begin // @[FADD_1.scala 21:40]
      isZeroA <= 1'h0; // @[FADD_1.scala 21:40]
    end else begin
      isZeroA <= mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA; // @[FADD_1.scala 46:67]
    end
    if (reset) begin // @[FADD_1.scala 22:43]
      isInfB <= 1'h0; // @[FADD_1.scala 22:43]
    end else begin
      isInfB <= mulAddRecFNToRaw_preMul_io_toPostMul_isInfB; // @[FADD_1.scala 47:70]
    end
    if (reset) begin // @[FADD_1.scala 23:40]
      isZeroB <= 1'h0; // @[FADD_1.scala 23:40]
    end else begin
      isZeroB <= mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB; // @[FADD_1.scala 48:67]
    end
    if (reset) begin // @[FADD_1.scala 24:38]
      signProd <= 1'h0; // @[FADD_1.scala 24:38]
    end else begin
      signProd <= mulAddRecFNToRaw_preMul_io_toPostMul_signProd; // @[FADD_1.scala 49:65]
    end
    if (reset) begin // @[FADD_1.scala 25:39]
      isNaNC <= 1'h0; // @[FADD_1.scala 25:39]
    end else begin
      isNaNC <= mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC; // @[FADD_1.scala 50:66]
    end
    if (reset) begin // @[FADD_1.scala 26:42]
      isInfC <= 1'h0; // @[FADD_1.scala 26:42]
    end else begin
      isInfC <= mulAddRecFNToRaw_preMul_io_toPostMul_isInfC; // @[FADD_1.scala 51:69]
    end
    if (reset) begin // @[FADD_1.scala 27:39]
      isZeroC <= 1'h0; // @[FADD_1.scala 27:39]
    end else begin
      isZeroC <= mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC; // @[FADD_1.scala 52:66]
    end
    if (reset) begin // @[FADD_1.scala 28:36]
      sExpSum <= 10'sh0; // @[FADD_1.scala 28:36]
    end else begin
      sExpSum <= mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum; // @[FADD_1.scala 53:63]
    end
    if (reset) begin // @[FADD_1.scala 29:33]
      doSubMags <= 1'h0; // @[FADD_1.scala 29:33]
    end else begin
      doSubMags <= mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags; // @[FADD_1.scala 54:60]
    end
    if (reset) begin // @[FADD_1.scala 30:33]
      CIsDominant <= 1'h0; // @[FADD_1.scala 30:33]
    end else begin
      CIsDominant <= mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant; // @[FADD_1.scala 55:59]
    end
    if (reset) begin // @[FADD_1.scala 31:34]
      CDom_CAlignDist <= 5'h0; // @[FADD_1.scala 31:34]
    end else begin
      CDom_CAlignDist <= mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist; // @[FADD_1.scala 56:54]
    end
    if (reset) begin // @[FADD_1.scala 32:37]
      highAlignedSigC <= 26'h0; // @[FADD_1.scala 32:37]
    end else begin
      highAlignedSigC <= mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC; // @[FADD_1.scala 57:56]
    end
    if (reset) begin // @[FADD_1.scala 33:38]
      bit0AlignedSigC <= 1'h0; // @[FADD_1.scala 33:38]
    end else begin
      bit0AlignedSigC <= mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC; // @[FADD_1.scala 58:57]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  premul_a = _RAND_0[23:0];
  _RAND_1 = {1{`RANDOM}};
  premul_b = _RAND_1[23:0];
  _RAND_2 = {2{`RANDOM}};
  premul_c = _RAND_2[47:0];
  _RAND_3 = {1{`RANDOM}};
  isSigNaNAny = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  isNaNAOrB = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  isInfA = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  isZeroA = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  isInfB = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  isZeroB = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  signProd = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  isNaNC = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  isInfC = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  isZeroC = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  sExpSum = _RAND_13[9:0];
  _RAND_14 = {1{`RANDOM}};
  doSubMags = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  CIsDominant = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  CDom_CAlignDist = _RAND_16[4:0];
  _RAND_17 = {1{`RANDOM}};
  highAlignedSigC = _RAND_17[25:0];
  _RAND_18 = {1{`RANDOM}};
  bit0AlignedSigC = _RAND_18[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IST0(
  input         clock,
  input         reset,
  input         io_enable_IST0,
  input  [31:0] io_nodeid_leaf,
  input  [31:0] io_rayid_leaf,
  input  [31:0] io_hiT_in,
  input  [31:0] io_v00_x,
  input  [31:0] io_v00_y,
  input  [31:0] io_v00_z,
  input  [31:0] io_v00_w,
  input  [31:0] io_v11_in_x,
  input  [31:0] io_v11_in_y,
  input  [31:0] io_v11_in_z,
  input  [31:0] io_v11_in_w,
  input  [31:0] io_v22_in_x,
  input  [31:0] io_v22_in_y,
  input  [31:0] io_v22_in_z,
  input  [31:0] io_v22_in_w,
  input  [31:0] io_ray_o_in_x,
  input  [31:0] io_ray_o_in_y,
  input  [31:0] io_ray_o_in_z,
  input  [31:0] io_ray_d_in_x,
  input  [31:0] io_ray_d_in_y,
  input  [31:0] io_ray_d_in_z,
  input         io_RAY_AABB_1,
  input         io_RAY_AABB_2,
  input         io_break_in,
  output [31:0] io_Oz,
  output [31:0] io_invDz_div,
  output [31:0] io_nodeid_ist0_out,
  output [31:0] io_rayid_ist0_out,
  output [31:0] io_hiT_out,
  output [31:0] io_v11_out_x,
  output [31:0] io_v11_out_y,
  output [31:0] io_v11_out_z,
  output [31:0] io_v11_out_w,
  output [31:0] io_v22_out_x,
  output [31:0] io_v22_out_y,
  output [31:0] io_v22_out_z,
  output [31:0] io_v22_out_w,
  output [31:0] io_ray_o_out_x,
  output [31:0] io_ray_o_out_y,
  output [31:0] io_ray_o_out_z,
  output [31:0] io_ray_d_out_x,
  output [31:0] io_ray_d_out_y,
  output [31:0] io_ray_d_out_z,
  output        io_enable_SU_out,
  output        io_break_out,
  output        io_RAY_AABB_1_out,
  output        io_RAY_AABB_2_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [127:0] _RAND_10;
  reg [127:0] _RAND_11;
  reg [95:0] _RAND_12;
  reg [95:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [127:0] _RAND_20;
  reg [127:0] _RAND_21;
  reg [95:0] _RAND_22;
  reg [95:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [127:0] _RAND_31;
  reg [127:0] _RAND_32;
  reg [95:0] _RAND_33;
  reg [95:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [127:0] _RAND_46;
  reg [127:0] _RAND_47;
  reg [95:0] _RAND_48;
  reg [95:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [127:0] _RAND_59;
  reg [127:0] _RAND_60;
  reg [95:0] _RAND_61;
  reg [95:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
`endif // RANDOMIZE_REG_INIT
  wire  FADD_MUL_13_clock; // @[IST0.scala 73:33]
  wire  FADD_MUL_13_reset; // @[IST0.scala 73:33]
  wire [31:0] FADD_MUL_13_io_a; // @[IST0.scala 73:33]
  wire [31:0] FADD_MUL_13_io_b; // @[IST0.scala 73:33]
  wire [31:0] FADD_MUL_13_io_c; // @[IST0.scala 73:33]
  wire [31:0] FADD_MUL_13_io_out; // @[IST0.scala 73:33]
  wire  FMUL_1_clock; // @[IST0.scala 79:24]
  wire  FMUL_1_reset; // @[IST0.scala 79:24]
  wire [31:0] FMUL_1_io_a; // @[IST0.scala 79:24]
  wire [31:0] FMUL_1_io_b; // @[IST0.scala 79:24]
  wire [31:0] FMUL_1_io_out; // @[IST0.scala 79:24]
  wire  FMUL_2_clock; // @[IST0.scala 84:24]
  wire  FMUL_2_reset; // @[IST0.scala 84:24]
  wire [31:0] FMUL_2_io_a; // @[IST0.scala 84:24]
  wire [31:0] FMUL_2_io_b; // @[IST0.scala 84:24]
  wire [31:0] FMUL_2_io_out; // @[IST0.scala 84:24]
  wire  FMUL_3_clock; // @[IST0.scala 89:24]
  wire  FMUL_3_reset; // @[IST0.scala 89:24]
  wire [31:0] FMUL_3_io_a; // @[IST0.scala 89:24]
  wire [31:0] FMUL_3_io_b; // @[IST0.scala 89:24]
  wire [31:0] FMUL_3_io_out; // @[IST0.scala 89:24]
  wire  FMUL_4_clock; // @[IST0.scala 94:24]
  wire  FMUL_4_reset; // @[IST0.scala 94:24]
  wire [31:0] FMUL_4_io_a; // @[IST0.scala 94:24]
  wire [31:0] FMUL_4_io_b; // @[IST0.scala 94:24]
  wire [31:0] FMUL_4_io_out; // @[IST0.scala 94:24]
  wire  FMUL_5_clock; // @[IST0.scala 99:24]
  wire  FMUL_5_reset; // @[IST0.scala 99:24]
  wire [31:0] FMUL_5_io_a; // @[IST0.scala 99:24]
  wire [31:0] FMUL_5_io_b; // @[IST0.scala 99:24]
  wire [31:0] FMUL_5_io_out; // @[IST0.scala 99:24]
  wire  FADD_1_clock; // @[IST0.scala 164:24]
  wire  FADD_1_reset; // @[IST0.scala 164:24]
  wire [31:0] FADD_1_io_a; // @[IST0.scala 164:24]
  wire [31:0] FADD_1_io_b; // @[IST0.scala 164:24]
  wire [31:0] FADD_1_io_out; // @[IST0.scala 164:24]
  wire  FADD_2_clock; // @[IST0.scala 173:24]
  wire  FADD_2_reset; // @[IST0.scala 173:24]
  wire [31:0] FADD_2_io_a; // @[IST0.scala 173:24]
  wire [31:0] FADD_2_io_b; // @[IST0.scala 173:24]
  wire [31:0] FADD_2_io_out; // @[IST0.scala 173:24]
  wire  FADD_3_clock; // @[IST0.scala 262:24]
  wire  FADD_3_reset; // @[IST0.scala 262:24]
  wire [31:0] FADD_3_io_a; // @[IST0.scala 262:24]
  wire [31:0] FADD_3_io_b; // @[IST0.scala 262:24]
  wire [31:0] FADD_3_io_out; // @[IST0.scala 262:24]
  wire  FADD_4_clock; // @[IST0.scala 271:24]
  wire  FADD_4_reset; // @[IST0.scala 271:24]
  wire [31:0] FADD_4_io_a; // @[IST0.scala 271:24]
  wire [31:0] FADD_4_io_b; // @[IST0.scala 271:24]
  wire [31:0] FADD_4_io_out; // @[IST0.scala 271:24]
  reg [31:0] temp_0; // @[IST0.scala 42:33]
  reg [31:0] temp_1; // @[IST0.scala 43:33]
  reg [31:0] temp_2; // @[IST0.scala 44:33]
  reg [31:0] temp_3; // @[IST0.scala 45:33]
  reg [31:0] temp_4; // @[IST0.scala 46:33]
  reg [31:0] temp_5; // @[IST0.scala 47:33]
  reg  enable_1; // @[IST0.scala 49:51]
  reg [31:0] nodeid_ist0_temp_1; // @[IST0.scala 50:38]
  reg [31:0] rayid_ist0_temp_1; // @[IST0.scala 51:41]
  reg [31:0] hitT_temp_1; // @[IST0.scala 52:47]
  reg [127:0] v11_1; // @[IST0.scala 53:56]
  reg [127:0] v22_1; // @[IST0.scala 54:56]
  reg [95:0] ray_o_in_1; // @[IST0.scala 55:50]
  reg [95:0] ray_d_in_1; // @[IST0.scala 56:50]
  reg  break_1; // @[IST0.scala 57:51]
  reg  ray_aabb_1; // @[IST0.scala 58:46]
  reg  ray_aabb_2; // @[IST0.scala 59:46]
  wire [127:0] _T = {io_v11_in_w,io_v11_in_z,io_v11_in_y,io_v11_in_x}; // @[Cat.scala 30:58]
  wire [127:0] _T_1 = {io_v22_in_w,io_v22_in_z,io_v22_in_y,io_v22_in_x}; // @[Cat.scala 30:58]
  wire [95:0] _T_2 = {io_ray_o_in_z,io_ray_o_in_y,io_ray_o_in_x}; // @[Cat.scala 30:58]
  wire [95:0] _T_3 = {io_ray_d_in_z,io_ray_d_in_y,io_ray_d_in_x}; // @[Cat.scala 30:58]
  wire  hi_4 = ~io_ray_o_in_x[31]; // @[common.scala 90:20]
  wire [30:0] lo_2 = io_ray_o_in_x[30:0]; // @[common.scala 90:30]
  reg [31:0] nodeid_ist0_temp_temp; // @[IST0.scala 104:41]
  reg [31:0] rayid_ist0_temp_temp; // @[IST0.scala 105:44]
  reg [31:0] hitT_temp_temp; // @[IST0.scala 106:50]
  reg [127:0] v11_temp; // @[IST0.scala 107:59]
  reg [127:0] v22_temp; // @[IST0.scala 108:59]
  reg [95:0] ray_o_in_temp; // @[IST0.scala 109:53]
  reg [95:0] ray_d_in_temp; // @[IST0.scala 110:53]
  reg  enable_temp; // @[IST0.scala 111:54]
  reg  break_temp; // @[IST0.scala 112:54]
  reg  ray_aabb_1_temp; // @[IST0.scala 113:46]
  reg  ray_aabb_2_temp; // @[IST0.scala 114:46]
  reg [31:0] nodeid_ist0_temp_2; // @[IST0.scala 131:38]
  reg [31:0] rayid_ist0_temp_2; // @[IST0.scala 132:41]
  reg [31:0] hitT_temp_2; // @[IST0.scala 133:47]
  reg [127:0] v11_2; // @[IST0.scala 134:56]
  reg [127:0] v22_2; // @[IST0.scala 135:56]
  reg [95:0] ray_o_in_2; // @[IST0.scala 136:50]
  reg [95:0] ray_d_in_2; // @[IST0.scala 137:50]
  reg  enable_2; // @[IST0.scala 138:51]
  reg  break_2; // @[IST0.scala 139:51]
  reg  ray_aabb_1_2; // @[IST0.scala 140:43]
  reg  ray_aabb_2_2; // @[IST0.scala 141:44]
  reg [31:0] temp_6; // @[IST0.scala 156:50]
  reg [31:0] temp_7; // @[IST0.scala 157:50]
  reg [31:0] temp_0_2; // @[IST0.scala 158:47]
  reg [31:0] temp_5_2; // @[IST0.scala 159:46]
  reg [31:0] add_nodeid_ist0_temp_2; // @[IST0.scala 182:42]
  reg [31:0] add_rayid_ist0_temp_2; // @[IST0.scala 183:45]
  reg [31:0] add_hitT_temp_2; // @[IST0.scala 184:51]
  reg [127:0] add_v11_2; // @[IST0.scala 185:60]
  reg [127:0] add_v22_2; // @[IST0.scala 186:60]
  reg [95:0] add_ray_o_in_2; // @[IST0.scala 187:54]
  reg [95:0] add_ray_d_in_2; // @[IST0.scala 188:54]
  reg  add_enable_2; // @[IST0.scala 189:55]
  reg  add_break_2; // @[IST0.scala 190:55]
  reg  add_ray_aabb_1_2; // @[IST0.scala 191:47]
  reg  add_ray_aabb_2_2; // @[IST0.scala 192:48]
  reg [31:0] add_temp_0_2; // @[IST0.scala 206:51]
  reg [31:0] add_temp_5_2; // @[IST0.scala 207:50]
  reg [31:0] add2_nodeid_ist0_temp_2; // @[IST0.scala 214:43]
  reg [31:0] add2_rayid_ist0_temp_2; // @[IST0.scala 215:46]
  reg [31:0] add2_hitT_temp_2; // @[IST0.scala 216:52]
  reg [127:0] add2_v11_2; // @[IST0.scala 217:61]
  reg [127:0] add2_v22_2; // @[IST0.scala 218:61]
  reg [95:0] add2_ray_o_in_2; // @[IST0.scala 219:55]
  reg [95:0] add2_ray_d_in_2; // @[IST0.scala 220:55]
  reg  add2_enable_2; // @[IST0.scala 221:56]
  reg  add2_break_2; // @[IST0.scala 222:56]
  reg  add2_ray_aabb_1_2; // @[IST0.scala 223:48]
  reg  add2_ray_aabb_2_2; // @[IST0.scala 224:49]
  wire  hi_5 = ~temp_6[31]; // @[common.scala 90:20]
  wire [30:0] lo_3 = temp_6[30:0]; // @[common.scala 90:30]
  MY_MULADD FADD_MUL_13 ( // @[IST0.scala 73:33]
    .clock(FADD_MUL_13_clock),
    .reset(FADD_MUL_13_reset),
    .io_a(FADD_MUL_13_io_a),
    .io_b(FADD_MUL_13_io_b),
    .io_c(FADD_MUL_13_io_c),
    .io_out(FADD_MUL_13_io_out)
  );
  MY_MUL FMUL_1 ( // @[IST0.scala 79:24]
    .clock(FMUL_1_clock),
    .reset(FMUL_1_reset),
    .io_a(FMUL_1_io_a),
    .io_b(FMUL_1_io_b),
    .io_out(FMUL_1_io_out)
  );
  MY_MUL FMUL_2 ( // @[IST0.scala 84:24]
    .clock(FMUL_2_clock),
    .reset(FMUL_2_reset),
    .io_a(FMUL_2_io_a),
    .io_b(FMUL_2_io_b),
    .io_out(FMUL_2_io_out)
  );
  MY_MUL FMUL_3 ( // @[IST0.scala 89:24]
    .clock(FMUL_3_clock),
    .reset(FMUL_3_reset),
    .io_a(FMUL_3_io_a),
    .io_b(FMUL_3_io_b),
    .io_out(FMUL_3_io_out)
  );
  MY_MUL FMUL_4 ( // @[IST0.scala 94:24]
    .clock(FMUL_4_clock),
    .reset(FMUL_4_reset),
    .io_a(FMUL_4_io_a),
    .io_b(FMUL_4_io_b),
    .io_out(FMUL_4_io_out)
  );
  MY_MUL FMUL_5 ( // @[IST0.scala 99:24]
    .clock(FMUL_5_clock),
    .reset(FMUL_5_reset),
    .io_a(FMUL_5_io_a),
    .io_b(FMUL_5_io_b),
    .io_out(FMUL_5_io_out)
  );
  MY_ADD FADD_1 ( // @[IST0.scala 164:24]
    .clock(FADD_1_clock),
    .reset(FADD_1_reset),
    .io_a(FADD_1_io_a),
    .io_b(FADD_1_io_b),
    .io_out(FADD_1_io_out)
  );
  MY_ADD FADD_2 ( // @[IST0.scala 173:24]
    .clock(FADD_2_clock),
    .reset(FADD_2_reset),
    .io_a(FADD_2_io_a),
    .io_b(FADD_2_io_b),
    .io_out(FADD_2_io_out)
  );
  MY_ADD FADD_3 ( // @[IST0.scala 262:24]
    .clock(FADD_3_clock),
    .reset(FADD_3_reset),
    .io_a(FADD_3_io_a),
    .io_b(FADD_3_io_b),
    .io_out(FADD_3_io_out)
  );
  MY_ADD FADD_4 ( // @[IST0.scala 271:24]
    .clock(FADD_4_clock),
    .reset(FADD_4_reset),
    .io_a(FADD_4_io_a),
    .io_b(FADD_4_io_b),
    .io_out(FADD_4_io_out)
  );
  assign io_Oz = FADD_3_io_out; // @[IST0.scala 269:29]
  assign io_invDz_div = FADD_4_io_out; // @[IST0.scala 278:22]
  assign io_nodeid_ist0_out = add2_nodeid_ist0_temp_2; // @[IST0.scala 238:32]
  assign io_rayid_ist0_out = add2_rayid_ist0_temp_2; // @[IST0.scala 239:35]
  assign io_hiT_out = add2_hitT_temp_2; // @[IST0.scala 240:42]
  assign io_v11_out_x = add2_v11_2[31:0]; // @[IST0.scala 241:53]
  assign io_v11_out_y = add2_v11_2[63:32]; // @[IST0.scala 242:53]
  assign io_v11_out_z = add2_v11_2[95:64]; // @[IST0.scala 243:53]
  assign io_v11_out_w = add2_v11_2[127:96]; // @[IST0.scala 244:52]
  assign io_v22_out_x = add2_v22_2[31:0]; // @[IST0.scala 246:57]
  assign io_v22_out_y = add2_v22_2[63:32]; // @[IST0.scala 247:57]
  assign io_v22_out_z = add2_v22_2[95:64]; // @[IST0.scala 248:57]
  assign io_v22_out_w = add2_v22_2[127:96]; // @[IST0.scala 249:55]
  assign io_ray_o_out_x = add2_ray_o_in_2[31:0]; // @[IST0.scala 252:59]
  assign io_ray_o_out_y = add2_ray_o_in_2[63:32]; // @[IST0.scala 253:59]
  assign io_ray_o_out_z = add2_ray_o_in_2[95:64]; // @[IST0.scala 254:59]
  assign io_ray_d_out_x = add2_ray_d_in_2[31:0]; // @[IST0.scala 255:59]
  assign io_ray_d_out_y = add2_ray_d_in_2[63:32]; // @[IST0.scala 256:59]
  assign io_ray_d_out_z = add2_ray_d_in_2[95:64]; // @[IST0.scala 257:59]
  assign io_enable_SU_out = add2_enable_2; // @[IST0.scala 258:36]
  assign io_break_out = add2_break_2; // @[IST0.scala 259:42]
  assign io_RAY_AABB_1_out = add2_ray_aabb_1_2; // @[IST0.scala 260:33]
  assign io_RAY_AABB_2_out = add2_ray_aabb_2_2; // @[IST0.scala 261:33]
  assign FADD_MUL_13_clock = clock;
  assign FADD_MUL_13_reset = reset;
  assign FADD_MUL_13_io_a = {hi_4,lo_2}; // @[Cat.scala 30:58]
  assign FADD_MUL_13_io_b = io_v00_x; // @[IST0.scala 75:26]
  assign FADD_MUL_13_io_c = io_v00_w; // @[IST0.scala 76:26]
  assign FMUL_1_clock = clock;
  assign FMUL_1_reset = reset;
  assign FMUL_1_io_a = io_ray_o_in_y; // @[IST0.scala 80:21]
  assign FMUL_1_io_b = io_v00_y; // @[IST0.scala 81:21]
  assign FMUL_2_clock = clock;
  assign FMUL_2_reset = reset;
  assign FMUL_2_io_a = io_ray_o_in_z; // @[IST0.scala 85:21]
  assign FMUL_2_io_b = io_v00_z; // @[IST0.scala 86:21]
  assign FMUL_3_clock = clock;
  assign FMUL_3_reset = reset;
  assign FMUL_3_io_a = io_ray_d_in_x; // @[IST0.scala 90:21]
  assign FMUL_3_io_b = io_v00_x; // @[IST0.scala 91:21]
  assign FMUL_4_clock = clock;
  assign FMUL_4_reset = reset;
  assign FMUL_4_io_a = io_ray_d_in_y; // @[IST0.scala 95:21]
  assign FMUL_4_io_b = io_v00_y; // @[IST0.scala 96:21]
  assign FMUL_5_clock = clock;
  assign FMUL_5_reset = reset;
  assign FMUL_5_io_a = io_ray_d_in_z; // @[IST0.scala 100:21]
  assign FMUL_5_io_b = io_v00_z; // @[IST0.scala 101:21]
  assign FADD_1_clock = clock;
  assign FADD_1_reset = reset;
  assign FADD_1_io_a = temp_1; // @[IST0.scala 165:21]
  assign FADD_1_io_b = temp_2; // @[IST0.scala 166:21]
  assign FADD_2_clock = clock;
  assign FADD_2_reset = reset;
  assign FADD_2_io_a = temp_3; // @[IST0.scala 174:21]
  assign FADD_2_io_b = temp_4; // @[IST0.scala 175:21]
  assign FADD_3_clock = clock;
  assign FADD_3_reset = reset;
  assign FADD_3_io_a = add_temp_0_2; // @[IST0.scala 263:21]
  assign FADD_3_io_b = {hi_5,lo_3}; // @[Cat.scala 30:58]
  assign FADD_4_clock = clock;
  assign FADD_4_reset = reset;
  assign FADD_4_io_a = add_temp_5_2; // @[IST0.scala 272:21]
  assign FADD_4_io_b = temp_7; // @[IST0.scala 273:21]
  always @(posedge clock) begin
    if (reset) begin // @[IST0.scala 42:33]
      temp_0 <= 32'h0; // @[IST0.scala 42:33]
    end else begin
      temp_0 <= FADD_MUL_13_io_out; // @[IST0.scala 77:42]
    end
    if (reset) begin // @[IST0.scala 43:33]
      temp_1 <= 32'h0; // @[IST0.scala 43:33]
    end else begin
      temp_1 <= FMUL_1_io_out; // @[IST0.scala 82:42]
    end
    if (reset) begin // @[IST0.scala 44:33]
      temp_2 <= 32'h0; // @[IST0.scala 44:33]
    end else begin
      temp_2 <= FMUL_2_io_out; // @[IST0.scala 87:42]
    end
    if (reset) begin // @[IST0.scala 45:33]
      temp_3 <= 32'h0; // @[IST0.scala 45:33]
    end else begin
      temp_3 <= FMUL_3_io_out; // @[IST0.scala 92:42]
    end
    if (reset) begin // @[IST0.scala 46:33]
      temp_4 <= 32'h0; // @[IST0.scala 46:33]
    end else begin
      temp_4 <= FMUL_4_io_out; // @[IST0.scala 97:42]
    end
    if (reset) begin // @[IST0.scala 47:33]
      temp_5 <= 32'h0; // @[IST0.scala 47:33]
    end else begin
      temp_5 <= FMUL_5_io_out; // @[IST0.scala 102:42]
    end
    if (reset) begin // @[IST0.scala 49:51]
      enable_1 <= 1'h0; // @[IST0.scala 49:51]
    end else begin
      enable_1 <= io_enable_IST0; // @[IST0.scala 68:42]
    end
    if (reset) begin // @[IST0.scala 50:38]
      nodeid_ist0_temp_1 <= 32'sh0; // @[IST0.scala 50:38]
    end else begin
      nodeid_ist0_temp_1 <= io_nodeid_leaf; // @[IST0.scala 61:29]
    end
    if (reset) begin // @[IST0.scala 51:41]
      rayid_ist0_temp_1 <= 32'h0; // @[IST0.scala 51:41]
    end else begin
      rayid_ist0_temp_1 <= io_rayid_leaf; // @[IST0.scala 62:32]
    end
    if (reset) begin // @[IST0.scala 52:47]
      hitT_temp_1 <= 32'h0; // @[IST0.scala 52:47]
    end else begin
      hitT_temp_1 <= io_hiT_in; // @[IST0.scala 63:38]
    end
    if (reset) begin // @[IST0.scala 53:56]
      v11_1 <= 128'h0; // @[IST0.scala 53:56]
    end else begin
      v11_1 <= _T; // @[IST0.scala 64:46]
    end
    if (reset) begin // @[IST0.scala 54:56]
      v22_1 <= 128'h0; // @[IST0.scala 54:56]
    end else begin
      v22_1 <= _T_1; // @[IST0.scala 65:46]
    end
    if (reset) begin // @[IST0.scala 55:50]
      ray_o_in_1 <= 96'h0; // @[IST0.scala 55:50]
    end else begin
      ray_o_in_1 <= _T_2; // @[IST0.scala 66:40]
    end
    if (reset) begin // @[IST0.scala 56:50]
      ray_d_in_1 <= 96'h0; // @[IST0.scala 56:50]
    end else begin
      ray_d_in_1 <= _T_3; // @[IST0.scala 67:40]
    end
    if (reset) begin // @[IST0.scala 57:51]
      break_1 <= 1'h0; // @[IST0.scala 57:51]
    end else begin
      break_1 <= io_break_in; // @[IST0.scala 69:44]
    end
    if (reset) begin // @[IST0.scala 58:46]
      ray_aabb_1 <= 1'h0; // @[IST0.scala 58:46]
    end else begin
      ray_aabb_1 <= io_RAY_AABB_1; // @[IST0.scala 70:40]
    end
    if (reset) begin // @[IST0.scala 59:46]
      ray_aabb_2 <= 1'h0; // @[IST0.scala 59:46]
    end else begin
      ray_aabb_2 <= io_RAY_AABB_2; // @[IST0.scala 71:40]
    end
    if (reset) begin // @[IST0.scala 104:41]
      nodeid_ist0_temp_temp <= 32'sh0; // @[IST0.scala 104:41]
    end else begin
      nodeid_ist0_temp_temp <= nodeid_ist0_temp_1; // @[IST0.scala 116:32]
    end
    if (reset) begin // @[IST0.scala 105:44]
      rayid_ist0_temp_temp <= 32'h0; // @[IST0.scala 105:44]
    end else begin
      rayid_ist0_temp_temp <= rayid_ist0_temp_1; // @[IST0.scala 117:35]
    end
    if (reset) begin // @[IST0.scala 106:50]
      hitT_temp_temp <= 32'h0; // @[IST0.scala 106:50]
    end else begin
      hitT_temp_temp <= hitT_temp_1; // @[IST0.scala 118:41]
    end
    if (reset) begin // @[IST0.scala 107:59]
      v11_temp <= 128'h0; // @[IST0.scala 107:59]
    end else begin
      v11_temp <= v11_1; // @[IST0.scala 119:49]
    end
    if (reset) begin // @[IST0.scala 108:59]
      v22_temp <= 128'h0; // @[IST0.scala 108:59]
    end else begin
      v22_temp <= v22_1; // @[IST0.scala 120:49]
    end
    if (reset) begin // @[IST0.scala 109:53]
      ray_o_in_temp <= 96'h0; // @[IST0.scala 109:53]
    end else begin
      ray_o_in_temp <= ray_o_in_1; // @[IST0.scala 121:43]
    end
    if (reset) begin // @[IST0.scala 110:53]
      ray_d_in_temp <= 96'h0; // @[IST0.scala 110:53]
    end else begin
      ray_d_in_temp <= ray_d_in_1; // @[IST0.scala 122:43]
    end
    if (reset) begin // @[IST0.scala 111:54]
      enable_temp <= 1'h0; // @[IST0.scala 111:54]
    end else begin
      enable_temp <= enable_1; // @[IST0.scala 123:45]
    end
    if (reset) begin // @[IST0.scala 112:54]
      break_temp <= 1'h0; // @[IST0.scala 112:54]
    end else begin
      break_temp <= break_1; // @[IST0.scala 124:47]
    end
    if (reset) begin // @[IST0.scala 113:46]
      ray_aabb_1_temp <= 1'h0; // @[IST0.scala 113:46]
    end else begin
      ray_aabb_1_temp <= ray_aabb_1; // @[IST0.scala 125:39]
    end
    if (reset) begin // @[IST0.scala 114:46]
      ray_aabb_2_temp <= 1'h0; // @[IST0.scala 114:46]
    end else begin
      ray_aabb_2_temp <= ray_aabb_2; // @[IST0.scala 126:39]
    end
    if (reset) begin // @[IST0.scala 131:38]
      nodeid_ist0_temp_2 <= 32'sh0; // @[IST0.scala 131:38]
    end else begin
      nodeid_ist0_temp_2 <= nodeid_ist0_temp_temp; // @[IST0.scala 143:29]
    end
    if (reset) begin // @[IST0.scala 132:41]
      rayid_ist0_temp_2 <= 32'h0; // @[IST0.scala 132:41]
    end else begin
      rayid_ist0_temp_2 <= rayid_ist0_temp_temp; // @[IST0.scala 144:32]
    end
    if (reset) begin // @[IST0.scala 133:47]
      hitT_temp_2 <= 32'h0; // @[IST0.scala 133:47]
    end else begin
      hitT_temp_2 <= hitT_temp_temp; // @[IST0.scala 145:38]
    end
    if (reset) begin // @[IST0.scala 134:56]
      v11_2 <= 128'h0; // @[IST0.scala 134:56]
    end else begin
      v11_2 <= v11_temp; // @[IST0.scala 146:46]
    end
    if (reset) begin // @[IST0.scala 135:56]
      v22_2 <= 128'h0; // @[IST0.scala 135:56]
    end else begin
      v22_2 <= v22_temp; // @[IST0.scala 147:46]
    end
    if (reset) begin // @[IST0.scala 136:50]
      ray_o_in_2 <= 96'h0; // @[IST0.scala 136:50]
    end else begin
      ray_o_in_2 <= ray_o_in_temp; // @[IST0.scala 148:40]
    end
    if (reset) begin // @[IST0.scala 137:50]
      ray_d_in_2 <= 96'h0; // @[IST0.scala 137:50]
    end else begin
      ray_d_in_2 <= ray_d_in_temp; // @[IST0.scala 149:40]
    end
    if (reset) begin // @[IST0.scala 138:51]
      enable_2 <= 1'h0; // @[IST0.scala 138:51]
    end else begin
      enable_2 <= enable_temp; // @[IST0.scala 152:42]
    end
    if (reset) begin // @[IST0.scala 139:51]
      break_2 <= 1'h0; // @[IST0.scala 139:51]
    end else begin
      break_2 <= break_temp; // @[IST0.scala 153:44]
    end
    if (reset) begin // @[IST0.scala 140:43]
      ray_aabb_1_2 <= 1'h0; // @[IST0.scala 140:43]
    end else begin
      ray_aabb_1_2 <= ray_aabb_1_temp; // @[IST0.scala 154:37]
    end
    if (reset) begin // @[IST0.scala 141:44]
      ray_aabb_2_2 <= 1'h0; // @[IST0.scala 141:44]
    end else begin
      ray_aabb_2_2 <= ray_aabb_2_temp; // @[IST0.scala 155:37]
    end
    if (reset) begin // @[IST0.scala 156:50]
      temp_6 <= 32'h0; // @[IST0.scala 156:50]
    end else begin
      temp_6 <= FADD_1_io_out; // @[IST0.scala 171:26]
    end
    if (reset) begin // @[IST0.scala 157:50]
      temp_7 <= 32'h0; // @[IST0.scala 157:50]
    end else begin
      temp_7 <= FADD_2_io_out; // @[IST0.scala 180:26]
    end
    if (reset) begin // @[IST0.scala 158:47]
      temp_0_2 <= 32'h0; // @[IST0.scala 158:47]
    end else begin
      temp_0_2 <= temp_0; // @[IST0.scala 161:41]
    end
    if (reset) begin // @[IST0.scala 159:46]
      temp_5_2 <= 32'h0; // @[IST0.scala 159:46]
    end else begin
      temp_5_2 <= temp_5; // @[IST0.scala 162:41]
    end
    if (reset) begin // @[IST0.scala 182:42]
      add_nodeid_ist0_temp_2 <= 32'sh0; // @[IST0.scala 182:42]
    end else begin
      add_nodeid_ist0_temp_2 <= nodeid_ist0_temp_2; // @[IST0.scala 194:33]
    end
    if (reset) begin // @[IST0.scala 183:45]
      add_rayid_ist0_temp_2 <= 32'h0; // @[IST0.scala 183:45]
    end else begin
      add_rayid_ist0_temp_2 <= rayid_ist0_temp_2; // @[IST0.scala 195:36]
    end
    if (reset) begin // @[IST0.scala 184:51]
      add_hitT_temp_2 <= 32'h0; // @[IST0.scala 184:51]
    end else begin
      add_hitT_temp_2 <= hitT_temp_2; // @[IST0.scala 196:42]
    end
    if (reset) begin // @[IST0.scala 185:60]
      add_v11_2 <= 128'h0; // @[IST0.scala 185:60]
    end else begin
      add_v11_2 <= v11_2; // @[IST0.scala 197:50]
    end
    if (reset) begin // @[IST0.scala 186:60]
      add_v22_2 <= 128'h0; // @[IST0.scala 186:60]
    end else begin
      add_v22_2 <= v22_2; // @[IST0.scala 198:50]
    end
    if (reset) begin // @[IST0.scala 187:54]
      add_ray_o_in_2 <= 96'h0; // @[IST0.scala 187:54]
    end else begin
      add_ray_o_in_2 <= ray_o_in_2; // @[IST0.scala 199:44]
    end
    if (reset) begin // @[IST0.scala 188:54]
      add_ray_d_in_2 <= 96'h0; // @[IST0.scala 188:54]
    end else begin
      add_ray_d_in_2 <= ray_d_in_2; // @[IST0.scala 200:44]
    end
    if (reset) begin // @[IST0.scala 189:55]
      add_enable_2 <= 1'h0; // @[IST0.scala 189:55]
    end else begin
      add_enable_2 <= enable_2; // @[IST0.scala 201:46]
    end
    if (reset) begin // @[IST0.scala 190:55]
      add_break_2 <= 1'h0; // @[IST0.scala 190:55]
    end else begin
      add_break_2 <= break_2; // @[IST0.scala 202:48]
    end
    if (reset) begin // @[IST0.scala 191:47]
      add_ray_aabb_1_2 <= 1'h0; // @[IST0.scala 191:47]
    end else begin
      add_ray_aabb_1_2 <= ray_aabb_1_2; // @[IST0.scala 203:41]
    end
    if (reset) begin // @[IST0.scala 192:48]
      add_ray_aabb_2_2 <= 1'h0; // @[IST0.scala 192:48]
    end else begin
      add_ray_aabb_2_2 <= ray_aabb_2_2; // @[IST0.scala 204:41]
    end
    if (reset) begin // @[IST0.scala 206:51]
      add_temp_0_2 <= 32'h0; // @[IST0.scala 206:51]
    end else begin
      add_temp_0_2 <= temp_0_2; // @[IST0.scala 209:45]
    end
    if (reset) begin // @[IST0.scala 207:50]
      add_temp_5_2 <= 32'h0; // @[IST0.scala 207:50]
    end else begin
      add_temp_5_2 <= temp_5_2; // @[IST0.scala 210:45]
    end
    if (reset) begin // @[IST0.scala 214:43]
      add2_nodeid_ist0_temp_2 <= 32'sh0; // @[IST0.scala 214:43]
    end else begin
      add2_nodeid_ist0_temp_2 <= add_nodeid_ist0_temp_2; // @[IST0.scala 226:34]
    end
    if (reset) begin // @[IST0.scala 215:46]
      add2_rayid_ist0_temp_2 <= 32'h0; // @[IST0.scala 215:46]
    end else begin
      add2_rayid_ist0_temp_2 <= add_rayid_ist0_temp_2; // @[IST0.scala 227:37]
    end
    if (reset) begin // @[IST0.scala 216:52]
      add2_hitT_temp_2 <= 32'h0; // @[IST0.scala 216:52]
    end else begin
      add2_hitT_temp_2 <= add_hitT_temp_2; // @[IST0.scala 228:43]
    end
    if (reset) begin // @[IST0.scala 217:61]
      add2_v11_2 <= 128'h0; // @[IST0.scala 217:61]
    end else begin
      add2_v11_2 <= add_v11_2; // @[IST0.scala 229:51]
    end
    if (reset) begin // @[IST0.scala 218:61]
      add2_v22_2 <= 128'h0; // @[IST0.scala 218:61]
    end else begin
      add2_v22_2 <= add_v22_2; // @[IST0.scala 230:51]
    end
    if (reset) begin // @[IST0.scala 219:55]
      add2_ray_o_in_2 <= 96'h0; // @[IST0.scala 219:55]
    end else begin
      add2_ray_o_in_2 <= add_ray_o_in_2; // @[IST0.scala 231:45]
    end
    if (reset) begin // @[IST0.scala 220:55]
      add2_ray_d_in_2 <= 96'h0; // @[IST0.scala 220:55]
    end else begin
      add2_ray_d_in_2 <= add_ray_d_in_2; // @[IST0.scala 232:45]
    end
    if (reset) begin // @[IST0.scala 221:56]
      add2_enable_2 <= 1'h0; // @[IST0.scala 221:56]
    end else begin
      add2_enable_2 <= add_enable_2; // @[IST0.scala 233:47]
    end
    if (reset) begin // @[IST0.scala 222:56]
      add2_break_2 <= 1'h0; // @[IST0.scala 222:56]
    end else begin
      add2_break_2 <= add_break_2; // @[IST0.scala 234:49]
    end
    if (reset) begin // @[IST0.scala 223:48]
      add2_ray_aabb_1_2 <= 1'h0; // @[IST0.scala 223:48]
    end else begin
      add2_ray_aabb_1_2 <= add_ray_aabb_1_2; // @[IST0.scala 235:42]
    end
    if (reset) begin // @[IST0.scala 224:49]
      add2_ray_aabb_2_2 <= 1'h0; // @[IST0.scala 224:49]
    end else begin
      add2_ray_aabb_2_2 <= add_ray_aabb_2_2; // @[IST0.scala 236:42]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  temp_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  temp_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  temp_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  temp_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  temp_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  temp_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  enable_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  nodeid_ist0_temp_1 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  rayid_ist0_temp_1 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  hitT_temp_1 = _RAND_9[31:0];
  _RAND_10 = {4{`RANDOM}};
  v11_1 = _RAND_10[127:0];
  _RAND_11 = {4{`RANDOM}};
  v22_1 = _RAND_11[127:0];
  _RAND_12 = {3{`RANDOM}};
  ray_o_in_1 = _RAND_12[95:0];
  _RAND_13 = {3{`RANDOM}};
  ray_d_in_1 = _RAND_13[95:0];
  _RAND_14 = {1{`RANDOM}};
  break_1 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  ray_aabb_1 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  ray_aabb_2 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  nodeid_ist0_temp_temp = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  rayid_ist0_temp_temp = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  hitT_temp_temp = _RAND_19[31:0];
  _RAND_20 = {4{`RANDOM}};
  v11_temp = _RAND_20[127:0];
  _RAND_21 = {4{`RANDOM}};
  v22_temp = _RAND_21[127:0];
  _RAND_22 = {3{`RANDOM}};
  ray_o_in_temp = _RAND_22[95:0];
  _RAND_23 = {3{`RANDOM}};
  ray_d_in_temp = _RAND_23[95:0];
  _RAND_24 = {1{`RANDOM}};
  enable_temp = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  break_temp = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  ray_aabb_1_temp = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  ray_aabb_2_temp = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  nodeid_ist0_temp_2 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  rayid_ist0_temp_2 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  hitT_temp_2 = _RAND_30[31:0];
  _RAND_31 = {4{`RANDOM}};
  v11_2 = _RAND_31[127:0];
  _RAND_32 = {4{`RANDOM}};
  v22_2 = _RAND_32[127:0];
  _RAND_33 = {3{`RANDOM}};
  ray_o_in_2 = _RAND_33[95:0];
  _RAND_34 = {3{`RANDOM}};
  ray_d_in_2 = _RAND_34[95:0];
  _RAND_35 = {1{`RANDOM}};
  enable_2 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  break_2 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  ray_aabb_1_2 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  ray_aabb_2_2 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  temp_6 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  temp_7 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  temp_0_2 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  temp_5_2 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  add_nodeid_ist0_temp_2 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  add_rayid_ist0_temp_2 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  add_hitT_temp_2 = _RAND_45[31:0];
  _RAND_46 = {4{`RANDOM}};
  add_v11_2 = _RAND_46[127:0];
  _RAND_47 = {4{`RANDOM}};
  add_v22_2 = _RAND_47[127:0];
  _RAND_48 = {3{`RANDOM}};
  add_ray_o_in_2 = _RAND_48[95:0];
  _RAND_49 = {3{`RANDOM}};
  add_ray_d_in_2 = _RAND_49[95:0];
  _RAND_50 = {1{`RANDOM}};
  add_enable_2 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  add_break_2 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  add_ray_aabb_1_2 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  add_ray_aabb_2_2 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  add_temp_0_2 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  add_temp_5_2 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  add2_nodeid_ist0_temp_2 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  add2_rayid_ist0_temp_2 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  add2_hitT_temp_2 = _RAND_58[31:0];
  _RAND_59 = {4{`RANDOM}};
  add2_v11_2 = _RAND_59[127:0];
  _RAND_60 = {4{`RANDOM}};
  add2_v22_2 = _RAND_60[127:0];
  _RAND_61 = {3{`RANDOM}};
  add2_ray_o_in_2 = _RAND_61[95:0];
  _RAND_62 = {3{`RANDOM}};
  add2_ray_d_in_2 = _RAND_62[95:0];
  _RAND_63 = {1{`RANDOM}};
  add2_enable_2 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  add2_break_2 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  add2_ray_aabb_1_2 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  add2_ray_aabb_2_2 = _RAND_66[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module lookupC(
  input  [5:0]  io_addr,
  output [23:0] io_out
);
  wire [9:0] _GEN_0 = io_addr == 6'h3f ? 10'h206 : 10'h0; // @[lookups.scala 386:43 lookups.scala 386:51 lookups.scala 387:27]
  wire [9:0] _GEN_1 = io_addr == 6'h3e ? 10'h212 : _GEN_0; // @[lookups.scala 385:43 lookups.scala 385:51]
  wire [9:0] _GEN_2 = io_addr == 6'h3d ? 10'h21f : _GEN_1; // @[lookups.scala 384:43 lookups.scala 384:51]
  wire [9:0] _GEN_3 = io_addr == 6'h3c ? 10'h22c : _GEN_2; // @[lookups.scala 383:43 lookups.scala 383:51]
  wire [9:0] _GEN_4 = io_addr == 6'h3b ? 10'h23a : _GEN_3; // @[lookups.scala 382:43 lookups.scala 382:51]
  wire [9:0] _GEN_5 = io_addr == 6'h3a ? 10'h248 : _GEN_4; // @[lookups.scala 381:43 lookups.scala 381:51]
  wire [9:0] _GEN_6 = io_addr == 6'h39 ? 10'h256 : _GEN_5; // @[lookups.scala 380:43 lookups.scala 380:51]
  wire [9:0] _GEN_7 = io_addr == 6'h38 ? 10'h265 : _GEN_6; // @[lookups.scala 379:43 lookups.scala 379:51]
  wire [9:0] _GEN_8 = io_addr == 6'h37 ? 10'h275 : _GEN_7; // @[lookups.scala 377:43 lookups.scala 377:51]
  wire [9:0] _GEN_9 = io_addr == 6'h36 ? 10'h285 : _GEN_8; // @[lookups.scala 376:43 lookups.scala 376:51]
  wire [9:0] _GEN_10 = io_addr == 6'h35 ? 10'h295 : _GEN_9; // @[lookups.scala 375:43 lookups.scala 375:51]
  wire [9:0] _GEN_11 = io_addr == 6'h34 ? 10'h2a7 : _GEN_10; // @[lookups.scala 374:43 lookups.scala 374:51]
  wire [9:0] _GEN_12 = io_addr == 6'h33 ? 10'h2b8 : _GEN_11; // @[lookups.scala 373:43 lookups.scala 373:51]
  wire [9:0] _GEN_13 = io_addr == 6'h32 ? 10'h2cb : _GEN_12; // @[lookups.scala 372:43 lookups.scala 372:51]
  wire [9:0] _GEN_14 = io_addr == 6'h31 ? 10'h2de : _GEN_13; // @[lookups.scala 371:43 lookups.scala 371:51]
  wire [9:0] _GEN_15 = io_addr == 6'h30 ? 10'h2f2 : _GEN_14; // @[lookups.scala 370:43 lookups.scala 370:51]
  wire [9:0] _GEN_16 = io_addr == 6'h2f ? 10'h306 : _GEN_15; // @[lookups.scala 368:43 lookups.scala 368:51]
  wire [9:0] _GEN_17 = io_addr == 6'h2e ? 10'h31b : _GEN_16; // @[lookups.scala 367:43 lookups.scala 367:51]
  wire [9:0] _GEN_18 = io_addr == 6'h2d ? 10'h331 : _GEN_17; // @[lookups.scala 366:43 lookups.scala 366:51]
  wire [9:0] _GEN_19 = io_addr == 6'h2c ? 10'h348 : _GEN_18; // @[lookups.scala 365:43 lookups.scala 365:51]
  wire [9:0] _GEN_20 = io_addr == 6'h2b ? 10'h360 : _GEN_19; // @[lookups.scala 364:43 lookups.scala 364:51]
  wire [9:0] _GEN_21 = io_addr == 6'h2a ? 10'h378 : _GEN_20; // @[lookups.scala 363:43 lookups.scala 363:51]
  wire [9:0] _GEN_22 = io_addr == 6'h29 ? 10'h392 : _GEN_21; // @[lookups.scala 362:43 lookups.scala 362:51]
  wire [9:0] _GEN_23 = io_addr == 6'h28 ? 10'h3ac : _GEN_22; // @[lookups.scala 361:43 lookups.scala 361:51]
  wire [9:0] _GEN_24 = io_addr == 6'h27 ? 10'h3c8 : _GEN_23; // @[lookups.scala 359:43 lookups.scala 359:51]
  wire [9:0] _GEN_25 = io_addr == 6'h26 ? 10'h3e5 : _GEN_24; // @[lookups.scala 358:43 lookups.scala 358:51]
  wire [10:0] _GEN_26 = io_addr == 6'h25 ? 11'h402 : {{1'd0}, _GEN_25}; // @[lookups.scala 357:43 lookups.scala 357:51]
  wire [10:0] _GEN_27 = io_addr == 6'h24 ? 11'h421 : _GEN_26; // @[lookups.scala 356:43 lookups.scala 356:51]
  wire [10:0] _GEN_28 = io_addr == 6'h23 ? 11'h442 : _GEN_27; // @[lookups.scala 355:43 lookups.scala 355:51]
  wire [10:0] _GEN_29 = io_addr == 6'h22 ? 11'h463 : _GEN_28; // @[lookups.scala 354:43 lookups.scala 354:51]
  wire [10:0] _GEN_30 = io_addr == 6'h21 ? 11'h486 : _GEN_29; // @[lookups.scala 353:43 lookups.scala 353:51]
  wire [10:0] _GEN_31 = io_addr == 6'h20 ? 11'h4aa : _GEN_30; // @[lookups.scala 352:43 lookups.scala 352:51]
  wire [10:0] _GEN_32 = io_addr == 6'h1f ? 11'h4d0 : _GEN_31; // @[lookups.scala 350:43 lookups.scala 350:51]
  wire [10:0] _GEN_33 = io_addr == 6'h1e ? 11'h4f8 : _GEN_32; // @[lookups.scala 349:43 lookups.scala 349:51]
  wire [10:0] _GEN_34 = io_addr == 6'h1d ? 11'h521 : _GEN_33; // @[lookups.scala 348:43 lookups.scala 348:51]
  wire [10:0] _GEN_35 = io_addr == 6'h1c ? 11'h54c : _GEN_34; // @[lookups.scala 347:43 lookups.scala 347:51]
  wire [10:0] _GEN_36 = io_addr == 6'h1b ? 11'h579 : _GEN_35; // @[lookups.scala 346:43 lookups.scala 346:51]
  wire [10:0] _GEN_37 = io_addr == 6'h1a ? 11'h5a8 : _GEN_36; // @[lookups.scala 345:43 lookups.scala 345:51]
  wire [10:0] _GEN_38 = io_addr == 6'h19 ? 11'h5d9 : _GEN_37; // @[lookups.scala 344:43 lookups.scala 344:51]
  wire [10:0] _GEN_39 = io_addr == 6'h18 ? 11'h60d : _GEN_38; // @[lookups.scala 343:43 lookups.scala 343:51]
  wire [10:0] _GEN_40 = io_addr == 6'h17 ? 11'h642 : _GEN_39; // @[lookups.scala 341:43 lookups.scala 341:51]
  wire [10:0] _GEN_41 = io_addr == 6'h16 ? 11'h67b : _GEN_40; // @[lookups.scala 340:43 lookups.scala 340:51]
  wire [10:0] _GEN_42 = io_addr == 6'h15 ? 11'h6b5 : _GEN_41; // @[lookups.scala 339:43 lookups.scala 339:51]
  wire [10:0] _GEN_43 = io_addr == 6'h14 ? 11'h6f3 : _GEN_42; // @[lookups.scala 338:43 lookups.scala 338:51]
  wire [10:0] _GEN_44 = io_addr == 6'h13 ? 11'h734 : _GEN_43; // @[lookups.scala 337:43 lookups.scala 337:51]
  wire [10:0] _GEN_45 = io_addr == 6'h12 ? 11'h778 : _GEN_44; // @[lookups.scala 336:43 lookups.scala 336:51]
  wire [10:0] _GEN_46 = io_addr == 6'h11 ? 11'h7bf : _GEN_45; // @[lookups.scala 335:43 lookups.scala 335:51]
  wire [11:0] _GEN_47 = io_addr == 6'h10 ? 12'h80a : {{1'd0}, _GEN_46}; // @[lookups.scala 334:43 lookups.scala 334:51]
  wire [11:0] _GEN_48 = io_addr == 6'hf ? 12'h859 : _GEN_47; // @[lookups.scala 332:43 lookups.scala 332:51]
  wire [11:0] _GEN_49 = io_addr == 6'he ? 12'h8ab : _GEN_48; // @[lookups.scala 331:43 lookups.scala 331:51]
  wire [11:0] _GEN_50 = io_addr == 6'hd ? 12'h902 : _GEN_49; // @[lookups.scala 330:43 lookups.scala 330:51]
  wire [11:0] _GEN_51 = io_addr == 6'hc ? 12'h95e : _GEN_50; // @[lookups.scala 329:43 lookups.scala 329:51]
  wire [11:0] _GEN_52 = io_addr == 6'hb ? 12'h9bf : _GEN_51; // @[lookups.scala 328:43 lookups.scala 328:51]
  wire [11:0] _GEN_53 = io_addr == 6'ha ? 12'ha24 : _GEN_52; // @[lookups.scala 327:43 lookups.scala 327:51]
  wire [11:0] _GEN_54 = io_addr == 6'h9 ? 12'ha90 : _GEN_53; // @[lookups.scala 326:43 lookups.scala 326:51]
  wire [11:0] _GEN_55 = io_addr == 6'h8 ? 12'hb01 : _GEN_54; // @[lookups.scala 325:43 lookups.scala 325:51]
  wire [11:0] _GEN_56 = io_addr == 6'h7 ? 12'hb79 : _GEN_55; // @[lookups.scala 323:43 lookups.scala 323:51]
  wire [11:0] _GEN_57 = io_addr == 6'h6 ? 12'hbf8 : _GEN_56; // @[lookups.scala 322:43 lookups.scala 322:51]
  wire [11:0] _GEN_58 = io_addr == 6'h5 ? 12'hc7e : _GEN_57; // @[lookups.scala 321:43 lookups.scala 321:51]
  wire [11:0] _GEN_59 = io_addr == 6'h4 ? 12'hd0c : _GEN_58; // @[lookups.scala 320:43 lookups.scala 320:51]
  wire [11:0] _GEN_60 = io_addr == 6'h3 ? 12'hda3 : _GEN_59; // @[lookups.scala 319:43 lookups.scala 319:51]
  wire [11:0] _GEN_61 = io_addr == 6'h2 ? 12'he43 : _GEN_60; // @[lookups.scala 318:43 lookups.scala 318:51]
  wire [11:0] _GEN_62 = io_addr == 6'h1 ? 12'heed : _GEN_61; // @[lookups.scala 317:43 lookups.scala 317:51]
  wire [11:0] _GEN_63 = io_addr == 6'h0 ? 12'hfa1 : _GEN_62; // @[lookups.scala 316:38 lookups.scala 316:46]
  assign io_out = {{12'd0}, _GEN_63}; // @[lookups.scala 316:38 lookups.scala 316:46]
endmodule
module lookupL(
  input  [5:0]  io_addr,
  output [26:0] io_out
);
  wire [26:0] _GEN_0 = io_addr == 6'h3f ? 27'h4081020 : 27'h0; // @[lookups.scala 134:43 lookups.scala 134:51 lookups.scala 135:27]
  wire [26:0] _GEN_1 = io_addr == 6'h3e ? 27'h4104104 : _GEN_0; // @[lookups.scala 133:43 lookups.scala 133:51]
  wire [26:0] _GEN_2 = io_addr == 6'h3d ? 27'h4189374 : _GEN_1; // @[lookups.scala 132:43 lookups.scala 132:51]
  wire [26:0] _GEN_3 = io_addr == 6'h3c ? 27'h4210842 : _GEN_2; // @[lookups.scala 131:43 lookups.scala 131:51]
  wire [26:0] _GEN_4 = io_addr == 6'h3b ? 27'h429a042 : _GEN_3; // @[lookups.scala 130:43 lookups.scala 130:51]
  wire [26:0] _GEN_5 = io_addr == 6'h3a ? 27'h4325c53 : _GEN_4; // @[lookups.scala 129:43 lookups.scala 129:51]
  wire [26:0] _GEN_6 = io_addr == 6'h39 ? 27'h43b3d5a : _GEN_5; // @[lookups.scala 128:43 lookups.scala 128:51]
  wire [26:0] _GEN_7 = io_addr == 6'h38 ? 27'h4444444 : _GEN_6; // @[lookups.scala 127:43 lookups.scala 127:51]
  wire [26:0] _GEN_8 = io_addr == 6'h37 ? 27'h44d7204 : _GEN_7; // @[lookups.scala 125:43 lookups.scala 125:51]
  wire [26:0] _GEN_9 = io_addr == 6'h36 ? 27'h456c797 : _GEN_8; // @[lookups.scala 124:43 lookups.scala 124:51]
  wire [26:0] _GEN_10 = io_addr == 6'h35 ? 27'h4604604 : _GEN_9; // @[lookups.scala 123:43 lookups.scala 123:51]
  wire [26:0] _GEN_11 = io_addr == 6'h34 ? 27'h469ee58 : _GEN_10; // @[lookups.scala 122:43 lookups.scala 122:51]
  wire [26:0] _GEN_12 = io_addr == 6'h33 ? 27'h473c1ab : _GEN_11; // @[lookups.scala 121:43 lookups.scala 121:51]
  wire [26:0] _GEN_13 = io_addr == 6'h32 ? 27'h47dc11f : _GEN_12; // @[lookups.scala 120:43 lookups.scala 120:51]
  wire [26:0] _GEN_14 = io_addr == 6'h31 ? 27'h487ede0 : _GEN_13; // @[lookups.scala 119:43 lookups.scala 119:51]
  wire [26:0] _GEN_15 = io_addr == 6'h30 ? 27'h4924924 : _GEN_14; // @[lookups.scala 118:43 lookups.scala 118:51]
  wire [26:0] _GEN_16 = io_addr == 6'h2f ? 27'h49cd42e : _GEN_15; // @[lookups.scala 116:43 lookups.scala 116:51]
  wire [26:0] _GEN_17 = io_addr == 6'h2e ? 27'h4a7904a : _GEN_16; // @[lookups.scala 115:43 lookups.scala 115:51]
  wire [26:0] _GEN_18 = io_addr == 6'h2d ? 27'h4b27ed3 : _GEN_17; // @[lookups.scala 114:43 lookups.scala 114:51]
  wire [26:0] _GEN_19 = io_addr == 6'h2c ? 27'h4bda12f : _GEN_18; // @[lookups.scala 113:43 lookups.scala 113:51]
  wire [26:0] _GEN_20 = io_addr == 6'h2b ? 27'h4c8f8d2 : _GEN_19; // @[lookups.scala 112:43 lookups.scala 112:51]
  wire [26:0] _GEN_21 = io_addr == 6'h2a ? 27'h4d4873e : _GEN_20; // @[lookups.scala 111:43 lookups.scala 111:51]
  wire [26:0] _GEN_22 = io_addr == 6'h29 ? 27'h4e04e04 : _GEN_21; // @[lookups.scala 110:43 lookups.scala 110:51]
  wire [26:0] _GEN_23 = io_addr == 6'h28 ? 27'h4ec4ec4 : _GEN_22; // @[lookups.scala 109:43 lookups.scala 109:51]
  wire [26:0] _GEN_24 = io_addr == 6'h27 ? 27'h4f88b2f : _GEN_23; // @[lookups.scala 107:43 lookups.scala 107:51]
  wire [26:0] _GEN_25 = io_addr == 6'h26 ? 27'h5050505 : _GEN_24; // @[lookups.scala 106:43 lookups.scala 106:51]
  wire [26:0] _GEN_26 = io_addr == 6'h25 ? 27'h511be19 : _GEN_25; // @[lookups.scala 105:43 lookups.scala 105:51]
  wire [26:0] _GEN_27 = io_addr == 6'h24 ? 27'h51eb851 : _GEN_26; // @[lookups.scala 104:43 lookups.scala 104:51]
  wire [26:0] _GEN_28 = io_addr == 6'h23 ? 27'h52bf5a8 : _GEN_27; // @[lookups.scala 103:43 lookups.scala 103:51]
  wire [26:0] _GEN_29 = io_addr == 6'h22 ? 27'h5397829 : _GEN_28; // @[lookups.scala 102:43 lookups.scala 102:51]
  wire [26:0] _GEN_30 = io_addr == 6'h21 ? 27'h54741fa : _GEN_29; // @[lookups.scala 101:43 lookups.scala 101:51]
  wire [26:0] _GEN_31 = io_addr == 6'h20 ? 27'h5555555 : _GEN_30; // @[lookups.scala 100:43 lookups.scala 100:51]
  wire [26:0] _GEN_32 = io_addr == 6'h1f ? 27'h563b48c : _GEN_31; // @[lookups.scala 98:43 lookups.scala 98:51]
  wire [26:0] _GEN_33 = io_addr == 6'h1e ? 27'h572620a : _GEN_32; // @[lookups.scala 97:43 lookups.scala 97:51]
  wire [26:0] _GEN_34 = io_addr == 6'h1d ? 27'h5816058 : _GEN_33; // @[lookups.scala 96:43 lookups.scala 96:51]
  wire [26:0] _GEN_35 = io_addr == 6'h1c ? 27'h590b216 : _GEN_34; // @[lookups.scala 95:43 lookups.scala 95:51]
  wire [26:0] _GEN_36 = io_addr == 6'h1b ? 27'h5a05a05 : _GEN_35; // @[lookups.scala 94:43 lookups.scala 94:51]
  wire [26:0] _GEN_37 = io_addr == 6'h1a ? 27'h5b05b05 : _GEN_36; // @[lookups.scala 93:43 lookups.scala 93:51]
  wire [26:0] _GEN_38 = io_addr == 6'h19 ? 27'h5c0b817 : _GEN_37; // @[lookups.scala 92:43 lookups.scala 92:51]
  wire [26:0] _GEN_39 = io_addr == 6'h18 ? 27'h5d1745d : _GEN_38; // @[lookups.scala 91:43 lookups.scala 91:51]
  wire [26:0] _GEN_40 = io_addr == 6'h17 ? 27'h5e29320 : _GEN_39; // @[lookups.scala 89:43 lookups.scala 89:51]
  wire [26:0] _GEN_41 = io_addr == 6'h16 ? 27'h5f417d0 : _GEN_40; // @[lookups.scala 88:43 lookups.scala 88:51]
  wire [26:0] _GEN_42 = io_addr == 6'h15 ? 27'h6060606 : _GEN_41; // @[lookups.scala 87:43 lookups.scala 87:51]
  wire [26:0] _GEN_43 = io_addr == 6'h14 ? 27'h6186186 : _GEN_42; // @[lookups.scala 86:43 lookups.scala 86:51]
  wire [26:0] _GEN_44 = io_addr == 6'h13 ? 27'h62b2e43 : _GEN_43; // @[lookups.scala 85:43 lookups.scala 85:51]
  wire [26:0] _GEN_45 = io_addr == 6'h12 ? 27'h63e7063 : _GEN_44; // @[lookups.scala 84:43 lookups.scala 84:51]
  wire [26:0] _GEN_46 = io_addr == 6'h11 ? 27'h6522c3f : _GEN_45; // @[lookups.scala 83:43 lookups.scala 83:51]
  wire [26:0] _GEN_47 = io_addr == 6'h10 ? 27'h6666666 : _GEN_46; // @[lookups.scala 82:43 lookups.scala 82:51]
  wire [26:0] _GEN_48 = io_addr == 6'hf ? 27'h67b23a5 : _GEN_47; // @[lookups.scala 80:43 lookups.scala 80:51]
  wire [26:0] _GEN_49 = io_addr == 6'he ? 27'h6906906 : _GEN_48; // @[lookups.scala 79:43 lookups.scala 79:51]
  wire [26:0] _GEN_50 = io_addr == 6'hd ? 27'h6a63bd8 : _GEN_49; // @[lookups.scala 78:43 lookups.scala 78:51]
  wire [26:0] _GEN_51 = io_addr == 6'hc ? 27'h6bca1af : _GEN_50; // @[lookups.scala 77:43 lookups.scala 77:51]
  wire [26:0] _GEN_52 = io_addr == 6'hb ? 27'h6d3a06d : _GEN_51; // @[lookups.scala 76:43 lookups.scala 76:51]
  wire [26:0] _GEN_53 = io_addr == 6'ha ? 27'h6eb3e45 : _GEN_52; // @[lookups.scala 75:43 lookups.scala 75:51]
  wire [26:0] _GEN_54 = io_addr == 6'h9 ? 27'h70381c0 : _GEN_53; // @[lookups.scala 74:43 lookups.scala 74:51]
  wire [26:0] _GEN_55 = io_addr == 6'h8 ? 27'h71c71c7 : _GEN_54; // @[lookups.scala 73:43 lookups.scala 73:51]
  wire [26:0] _GEN_56 = io_addr == 6'h7 ? 27'h73615a2 : _GEN_55; // @[lookups.scala 71:43 lookups.scala 71:51]
  wire [26:0] _GEN_57 = io_addr == 6'h6 ? 27'h7507507 : _GEN_56; // @[lookups.scala 70:43 lookups.scala 70:51]
  wire [26:0] _GEN_58 = io_addr == 6'h5 ? 27'h76b981d : _GEN_57; // @[lookups.scala 69:43 lookups.scala 69:51]
  wire [26:0] _GEN_59 = io_addr == 6'h4 ? 27'h7878787 : _GEN_58; // @[lookups.scala 68:43 lookups.scala 68:51]
  wire [26:0] _GEN_60 = io_addr == 6'h3 ? 27'h7a44c6a : _GEN_59; // @[lookups.scala 67:43 lookups.scala 67:51]
  wire [26:0] _GEN_61 = io_addr == 6'h2 ? 27'h7c1f07c : _GEN_60; // @[lookups.scala 66:43 lookups.scala 66:51]
  wire [26:0] _GEN_62 = io_addr == 6'h1 ? 27'h7e07e07 : _GEN_61; // @[lookups.scala 65:43 lookups.scala 65:51]
  assign io_out = io_addr == 6'h0 ? 27'h0 : _GEN_62; // @[lookups.scala 64:38 lookups.scala 64:46]
endmodule
module lookupJ(
  input  [5:0]  io_addr,
  output [22:0] io_out
);
  wire [15:0] _GEN_0 = io_addr == 6'h3f ? 16'h8205 : 16'h0; // @[lookups.scala 261:43 lookups.scala 261:51 lookups.scala 262:27]
  wire [15:0] _GEN_1 = io_addr == 6'h3e ? 16'h8417 : _GEN_0; // @[lookups.scala 260:43 lookups.scala 260:51]
  wire [15:0] _GEN_2 = io_addr == 6'h3d ? 16'h8636 : _GEN_1; // @[lookups.scala 259:43 lookups.scala 259:51]
  wire [15:0] _GEN_3 = io_addr == 6'h3c ? 16'h8863 : _GEN_2; // @[lookups.scala 258:43 lookups.scala 258:51]
  wire [15:0] _GEN_4 = io_addr == 6'h3b ? 16'h8a9d : _GEN_3; // @[lookups.scala 257:43 lookups.scala 257:51]
  wire [15:0] _GEN_5 = io_addr == 6'h3a ? 16'h8ce5 : _GEN_4; // @[lookups.scala 256:43 lookups.scala 256:51]
  wire [15:0] _GEN_6 = io_addr == 6'h39 ? 16'h8f3b : _GEN_5; // @[lookups.scala 255:43 lookups.scala 255:51]
  wire [15:0] _GEN_7 = io_addr == 6'h38 ? 16'h91a1 : _GEN_6; // @[lookups.scala 254:43 lookups.scala 254:51]
  wire [15:0] _GEN_8 = io_addr == 6'h37 ? 16'h9416 : _GEN_7; // @[lookups.scala 252:43 lookups.scala 252:51]
  wire [15:0] _GEN_9 = io_addr == 6'h36 ? 16'h969b : _GEN_8; // @[lookups.scala 251:43 lookups.scala 251:51]
  wire [15:0] _GEN_10 = io_addr == 6'h35 ? 16'h9931 : _GEN_9; // @[lookups.scala 250:43 lookups.scala 250:51]
  wire [15:0] _GEN_11 = io_addr == 6'h34 ? 16'h9bd8 : _GEN_10; // @[lookups.scala 249:43 lookups.scala 249:51]
  wire [15:0] _GEN_12 = io_addr == 6'h33 ? 16'h9e91 : _GEN_11; // @[lookups.scala 248:43 lookups.scala 248:51]
  wire [15:0] _GEN_13 = io_addr == 6'h32 ? 16'ha15c : _GEN_12; // @[lookups.scala 247:43 lookups.scala 247:51]
  wire [15:0] _GEN_14 = io_addr == 6'h31 ? 16'ha43b : _GEN_13; // @[lookups.scala 246:43 lookups.scala 246:51]
  wire [15:0] _GEN_15 = io_addr == 6'h30 ? 16'ha72d : _GEN_14; // @[lookups.scala 245:43 lookups.scala 245:51]
  wire [15:0] _GEN_16 = io_addr == 6'h2f ? 16'haa33 : _GEN_15; // @[lookups.scala 243:43 lookups.scala 243:51]
  wire [15:0] _GEN_17 = io_addr == 6'h2e ? 16'had4f : _GEN_16; // @[lookups.scala 242:43 lookups.scala 242:51]
  wire [15:0] _GEN_18 = io_addr == 6'h2d ? 16'hb081 : _GEN_17; // @[lookups.scala 241:43 lookups.scala 241:51]
  wire [15:0] _GEN_19 = io_addr == 6'h2c ? 16'hb3ca : _GEN_18; // @[lookups.scala 240:43 lookups.scala 240:51]
  wire [15:0] _GEN_20 = io_addr == 6'h2b ? 16'hb72a : _GEN_19; // @[lookups.scala 239:43 lookups.scala 239:51]
  wire [15:0] _GEN_21 = io_addr == 6'h2a ? 16'hbaa3 : _GEN_20; // @[lookups.scala 238:43 lookups.scala 238:51]
  wire [15:0] _GEN_22 = io_addr == 6'h29 ? 16'hbe35 : _GEN_21; // @[lookups.scala 237:43 lookups.scala 237:51]
  wire [15:0] _GEN_23 = io_addr == 6'h28 ? 16'hc1e2 : _GEN_22; // @[lookups.scala 236:43 lookups.scala 236:51]
  wire [15:0] _GEN_24 = io_addr == 6'h27 ? 16'hc5aa : _GEN_23; // @[lookups.scala 234:43 lookups.scala 234:51]
  wire [15:0] _GEN_25 = io_addr == 6'h26 ? 16'hc98f : _GEN_24; // @[lookups.scala 233:43 lookups.scala 233:51]
  wire [15:0] _GEN_26 = io_addr == 6'h25 ? 16'hcd92 : _GEN_25; // @[lookups.scala 232:43 lookups.scala 232:51]
  wire [15:0] _GEN_27 = io_addr == 6'h24 ? 16'hd1b4 : _GEN_26; // @[lookups.scala 231:43 lookups.scala 231:51]
  wire [15:0] _GEN_28 = io_addr == 6'h23 ? 16'hd5f6 : _GEN_27; // @[lookups.scala 230:43 lookups.scala 230:51]
  wire [15:0] _GEN_29 = io_addr == 6'h22 ? 16'hda59 : _GEN_28; // @[lookups.scala 229:43 lookups.scala 229:51]
  wire [15:0] _GEN_30 = io_addr == 6'h21 ? 16'hdee0 : _GEN_29; // @[lookups.scala 228:43 lookups.scala 228:51]
  wire [15:0] _GEN_31 = io_addr == 6'h20 ? 16'he38b : _GEN_30; // @[lookups.scala 227:43 lookups.scala 227:51]
  wire [15:0] _GEN_32 = io_addr == 6'h1f ? 16'he85b : _GEN_31; // @[lookups.scala 225:43 lookups.scala 225:51]
  wire [15:0] _GEN_33 = io_addr == 6'h1e ? 16'hed54 : _GEN_32; // @[lookups.scala 224:43 lookups.scala 224:51]
  wire [15:0] _GEN_34 = io_addr == 6'h1d ? 16'hf275 : _GEN_33; // @[lookups.scala 223:43 lookups.scala 223:51]
  wire [15:0] _GEN_35 = io_addr == 6'h1c ? 16'hf7c2 : _GEN_34; // @[lookups.scala 222:43 lookups.scala 222:51]
  wire [15:0] _GEN_36 = io_addr == 6'h1b ? 16'hfd3b : _GEN_35; // @[lookups.scala 221:43 lookups.scala 221:51]
  wire [16:0] _GEN_37 = io_addr == 6'h1a ? 17'h102e4 : {{1'd0}, _GEN_36}; // @[lookups.scala 220:43 lookups.scala 220:51]
  wire [16:0] _GEN_38 = io_addr == 6'h19 ? 17'h108bd : _GEN_37; // @[lookups.scala 219:43 lookups.scala 219:51]
  wire [16:0] _GEN_39 = io_addr == 6'h18 ? 17'h10eca : _GEN_38; // @[lookups.scala 218:43 lookups.scala 218:51]
  wire [16:0] _GEN_40 = io_addr == 6'h17 ? 17'h1150d : _GEN_39; // @[lookups.scala 216:43 lookups.scala 216:51]
  wire [16:0] _GEN_41 = io_addr == 6'h16 ? 17'h11b88 : _GEN_40; // @[lookups.scala 215:43 lookups.scala 215:51]
  wire [16:0] _GEN_42 = io_addr == 6'h15 ? 17'h1223e : _GEN_41; // @[lookups.scala 214:43 lookups.scala 214:51]
  wire [16:0] _GEN_43 = io_addr == 6'h14 ? 17'h12931 : _GEN_42; // @[lookups.scala 213:43 lookups.scala 213:51]
  wire [16:0] _GEN_44 = io_addr == 6'h13 ? 17'h13066 : _GEN_43; // @[lookups.scala 212:43 lookups.scala 212:51]
  wire [16:0] _GEN_45 = io_addr == 6'h12 ? 17'h137de : _GEN_44; // @[lookups.scala 211:43 lookups.scala 211:51]
  wire [16:0] _GEN_46 = io_addr == 6'h11 ? 17'h13f9d : _GEN_45; // @[lookups.scala 210:43 lookups.scala 210:51]
  wire [16:0] _GEN_47 = io_addr == 6'h10 ? 17'h147a7 : _GEN_46; // @[lookups.scala 209:43 lookups.scala 209:51]
  wire [16:0] _GEN_48 = io_addr == 6'hf ? 17'h15000 : _GEN_47; // @[lookups.scala 207:43 lookups.scala 207:51]
  wire [16:0] _GEN_49 = io_addr == 6'he ? 17'h158ab : _GEN_48; // @[lookups.scala 206:43 lookups.scala 206:51]
  wire [16:0] _GEN_50 = io_addr == 6'hd ? 17'h161ae : _GEN_49; // @[lookups.scala 205:43 lookups.scala 205:51]
  wire [16:0] _GEN_51 = io_addr == 6'hc ? 17'h16b0c : _GEN_50; // @[lookups.scala 204:43 lookups.scala 204:51]
  wire [16:0] _GEN_52 = io_addr == 6'hb ? 17'h174cb : _GEN_51; // @[lookups.scala 203:43 lookups.scala 203:51]
  wire [16:0] _GEN_53 = io_addr == 6'ha ? 17'h17eef : _GEN_52; // @[lookups.scala 202:43 lookups.scala 202:51]
  wire [16:0] _GEN_54 = io_addr == 6'h9 ? 17'h1897f : _GEN_53; // @[lookups.scala 201:43 lookups.scala 201:51]
  wire [16:0] _GEN_55 = io_addr == 6'h8 ? 17'h19481 : _GEN_54; // @[lookups.scala 200:43 lookups.scala 200:51]
  wire [16:0] _GEN_56 = io_addr == 6'h7 ? 17'h19ffa : _GEN_55; // @[lookups.scala 198:43 lookups.scala 198:51]
  wire [16:0] _GEN_57 = io_addr == 6'h6 ? 17'h1abf2 : _GEN_56; // @[lookups.scala 197:43 lookups.scala 197:51]
  wire [16:0] _GEN_58 = io_addr == 6'h5 ? 17'h1b870 : _GEN_57; // @[lookups.scala 196:43 lookups.scala 196:51]
  wire [16:0] _GEN_59 = io_addr == 6'h4 ? 17'h1c57d : _GEN_58; // @[lookups.scala 195:43 lookups.scala 195:51]
  wire [16:0] _GEN_60 = io_addr == 6'h3 ? 17'h1d31f : _GEN_59; // @[lookups.scala 194:43 lookups.scala 194:51]
  wire [16:0] _GEN_61 = io_addr == 6'h2 ? 17'h1e162 : _GEN_60; // @[lookups.scala 193:43 lookups.scala 193:51]
  wire [16:0] _GEN_62 = io_addr == 6'h1 ? 17'h1f04f : _GEN_61; // @[lookups.scala 192:43 lookups.scala 192:51]
  wire [16:0] _GEN_63 = io_addr == 6'h0 ? 17'h1fff0 : _GEN_62; // @[lookups.scala 191:38 lookups.scala 191:46]
  assign io_out = {{6'd0}, _GEN_63}; // @[lookups.scala 191:38 lookups.scala 191:46]
endmodule
module VarSizeMul(
  input  [22:0] io_in1,
  input  [16:0] io_in2,
  output [23:0] io_out
);
  wire [22:0] _GEN_0 = {{6'd0}, io_in2}; // @[VarSizeMul.scala 20:26]
  wire [39:0] result = io_in1 * _GEN_0; // @[VarSizeMul.scala 20:26]
  assign io_out = result[39:16]; // @[VarSizeMul.scala 22:25]
endmodule
module mul2(
  input  [23:0] io_in1,
  input  [16:0] io_in2,
  output [28:0] io_out
);
  wire [23:0] _GEN_0 = {{7'd0}, io_in2}; // @[VarSizeMul.scala 37:26]
  wire [40:0] result = io_in1 * _GEN_0; // @[VarSizeMul.scala 37:26]
  assign io_out = result[40:12]; // @[VarSizeMul.scala 38:25]
endmodule
module VarSizeSub(
  input  [26:0] io_in1,
  input  [26:0] io_in2,
  output [26:0] io_out
);
  assign io_out = io_in1 + io_in2; // @[VarSizeAdder.scala 36:27]
endmodule
module VarSizeAdder(
  input  [28:0] io_in1,
  input  [28:0] io_in2,
  output [24:0] io_out
);
  wire [28:0] _T_1 = io_in1 + io_in2; // @[VarSizeAdder.scala 21:27]
  assign io_out = _T_1[28:4]; // @[VarSizeAdder.scala 21:36]
endmodule
module mul3(
  input  [22:0] io_in1,
  input  [24:0] io_in2,
  output [23:0] io_out
);
  wire [24:0] _GEN_0 = {{2'd0}, io_in1}; // @[VarSizeMul.scala 54:26]
  wire [47:0] result = _GEN_0 * io_in2; // @[VarSizeMul.scala 54:26]
  assign io_out = result[47:24]; // @[VarSizeMul.scala 55:25]
endmodule
module fpInverter(
  input         clock,
  input         reset,
  input  [22:0] io_in1,
  output [23:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire [5:0] tableC_io_addr; // @[fpInverter.scala 19:28]
  wire [23:0] tableC_io_out; // @[fpInverter.scala 19:28]
  wire [5:0] tableL_io_addr; // @[fpInverter.scala 20:28]
  wire [26:0] tableL_io_out; // @[fpInverter.scala 20:28]
  wire [5:0] tableJ_io_addr; // @[fpInverter.scala 21:28]
  wire [22:0] tableJ_io_out; // @[fpInverter.scala 21:28]
  wire [22:0] mul1_io_in1; // @[fpInverter.scala 32:26]
  wire [16:0] mul1_io_in2; // @[fpInverter.scala 32:26]
  wire [23:0] mul1_io_out; // @[fpInverter.scala 32:26]
  wire [23:0] mul2_io_in1; // @[fpInverter.scala 37:26]
  wire [16:0] mul2_io_in2; // @[fpInverter.scala 37:26]
  wire [28:0] mul2_io_out; // @[fpInverter.scala 37:26]
  wire [26:0] sub2_io_in1; // @[fpInverter.scala 65:30]
  wire [26:0] sub2_io_in2; // @[fpInverter.scala 65:30]
  wire [26:0] sub2_io_out; // @[fpInverter.scala 65:30]
  wire [28:0] adder_io_in1; // @[fpInverter.scala 74:31]
  wire [28:0] adder_io_in2; // @[fpInverter.scala 74:31]
  wire [24:0] adder_io_out; // @[fpInverter.scala 74:31]
  wire [22:0] mul3_io_in1; // @[fpInverter.scala 89:30]
  wire [24:0] mul3_io_in2; // @[fpInverter.scala 89:30]
  wire [23:0] mul3_io_out; // @[fpInverter.scala 89:30]
  wire [22:0] _T = io_in1 ^ 23'h7fffff; // @[fpInverter.scala 30:28]
  wire [33:0] _T_5 = io_in1[16:0] * io_in1[16:0]; // @[fpInverter.scala 39:42]
  reg [22:0] w_sub1_reg; // @[fpInverter.scala 43:41]
  reg [23:0] w_mul1_reg; // @[fpInverter.scala 44:41]
  reg [28:0] w_mul2_reg; // @[fpInverter.scala 45:41]
  reg [26:0] tableL_out_reg; // @[fpInverter.scala 57:37]
  reg [22:0] sub1_out_reg1; // @[fpInverter.scala 59:37]
  reg [23:0] mul1_out_reg; // @[fpInverter.scala 60:37]
  reg [28:0] mul2_out_reg; // @[fpInverter.scala 61:37]
  wire [23:0] _T_7 = mul1_out_reg ^ 24'hffffff; // @[fpInverter.scala 66:38]
  wire [23:0] sub2_in2 = _T_7 + 24'h1; // @[fpInverter.scala 66:71]
  wire [25:0] temp4 = {sub2_in2,1'h0,1'h0}; // @[Cat.scala 30:58]
  wire [27:0] temp1 = {sub2_io_out,1'h0}; // @[Cat.scala 30:58]
  reg [22:0] sub1_out_reg2; // @[fpInverter.scala 82:36]
  reg [24:0] adder_out_reg; // @[fpInverter.scala 85:36]
  reg [24:0] adder_out_reg_2; // @[fpInverter.scala 87:38]
  lookupC tableC ( // @[fpInverter.scala 19:28]
    .io_addr(tableC_io_addr),
    .io_out(tableC_io_out)
  );
  lookupL tableL ( // @[fpInverter.scala 20:28]
    .io_addr(tableL_io_addr),
    .io_out(tableL_io_out)
  );
  lookupJ tableJ ( // @[fpInverter.scala 21:28]
    .io_addr(tableJ_io_addr),
    .io_out(tableJ_io_out)
  );
  VarSizeMul mul1 ( // @[fpInverter.scala 32:26]
    .io_in1(mul1_io_in1),
    .io_in2(mul1_io_in2),
    .io_out(mul1_io_out)
  );
  mul2 mul2 ( // @[fpInverter.scala 37:26]
    .io_in1(mul2_io_in1),
    .io_in2(mul2_io_in2),
    .io_out(mul2_io_out)
  );
  VarSizeSub sub2 ( // @[fpInverter.scala 65:30]
    .io_in1(sub2_io_in1),
    .io_in2(sub2_io_in2),
    .io_out(sub2_io_out)
  );
  VarSizeAdder adder ( // @[fpInverter.scala 74:31]
    .io_in1(adder_io_in1),
    .io_in2(adder_io_in2),
    .io_out(adder_io_out)
  );
  mul3 mul3 ( // @[fpInverter.scala 89:30]
    .io_in1(mul3_io_in1),
    .io_in2(mul3_io_in2),
    .io_out(mul3_io_out)
  );
  assign io_out = mul3_io_out; // @[fpInverter.scala 97:16]
  assign tableC_io_addr = io_in1[22:17]; // @[fpInverter.scala 25:33]
  assign tableL_io_addr = io_in1[22:17]; // @[fpInverter.scala 25:33]
  assign tableJ_io_addr = io_in1[22:17]; // @[fpInverter.scala 25:33]
  assign mul1_io_in1 = tableJ_io_out; // @[fpInverter.scala 33:21]
  assign mul1_io_in2 = io_in1[16:0]; // @[fpInverter.scala 34:30]
  assign mul2_io_in1 = tableC_io_out; // @[fpInverter.scala 38:21]
  assign mul2_io_in2 = _T_5[33:17]; // @[fpInverter.scala 39:61]
  assign sub2_io_in1 = tableL_out_reg; // @[fpInverter.scala 70:21]
  assign sub2_io_in2 = {temp4,1'h0}; // @[Cat.scala 30:58]
  assign adder_io_in1 = {temp1,1'h0}; // @[Cat.scala 30:58]
  assign adder_io_in2 = mul2_out_reg; // @[fpInverter.scala 78:22]
  assign mul3_io_in1 = sub1_out_reg2; // @[fpInverter.scala 91:21]
  assign mul3_io_in2 = adder_out_reg_2; // @[fpInverter.scala 92:21]
  always @(posedge clock) begin
    w_sub1_reg <= _T + 23'h1; // @[fpInverter.scala 30:60]
    w_mul1_reg <= mul1_io_out; // @[fpInverter.scala 44:41]
    w_mul2_reg <= mul2_io_out; // @[fpInverter.scala 45:41]
    tableL_out_reg <= tableL_io_out; // @[fpInverter.scala 57:37]
    sub1_out_reg1 <= w_sub1_reg; // @[fpInverter.scala 59:37]
    mul1_out_reg <= w_mul1_reg; // @[fpInverter.scala 60:37]
    mul2_out_reg <= w_mul2_reg; // @[fpInverter.scala 61:37]
    sub1_out_reg2 <= sub1_out_reg1; // @[fpInverter.scala 82:36]
    if (reset) begin // @[fpInverter.scala 85:36]
      adder_out_reg <= 25'h0; // @[fpInverter.scala 85:36]
    end else begin
      adder_out_reg <= adder_io_out; // @[fpInverter.scala 86:25]
    end
    if (reset) begin // @[fpInverter.scala 87:38]
      adder_out_reg_2 <= 25'h0; // @[fpInverter.scala 87:38]
    end else begin
      adder_out_reg_2 <= adder_out_reg; // @[fpInverter.scala 88:25]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  w_sub1_reg = _RAND_0[22:0];
  _RAND_1 = {1{`RANDOM}};
  w_mul1_reg = _RAND_1[23:0];
  _RAND_2 = {1{`RANDOM}};
  w_mul2_reg = _RAND_2[28:0];
  _RAND_3 = {1{`RANDOM}};
  tableL_out_reg = _RAND_3[26:0];
  _RAND_4 = {1{`RANDOM}};
  sub1_out_reg1 = _RAND_4[22:0];
  _RAND_5 = {1{`RANDOM}};
  mul1_out_reg = _RAND_5[23:0];
  _RAND_6 = {1{`RANDOM}};
  mul2_out_reg = _RAND_6[28:0];
  _RAND_7 = {1{`RANDOM}};
  sub1_out_reg2 = _RAND_7[22:0];
  _RAND_8 = {1{`RANDOM}};
  adder_out_reg = _RAND_8[24:0];
  _RAND_9 = {1{`RANDOM}};
  adder_out_reg_2 = _RAND_9[24:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module fp_inverter(
  input         clock,
  input         reset,
  input  [31:0] io_in1,
  output [31:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire  inverter_clock; // @[FP_inverter.scala 14:29]
  wire  inverter_reset; // @[FP_inverter.scala 14:29]
  wire [22:0] inverter_io_in1; // @[FP_inverter.scala 14:29]
  wire [23:0] inverter_io_out; // @[FP_inverter.scala 14:29]
  reg [7:0] in2ExpReg0; // @[FP_inverter.scala 18:42]
  reg  in2SignReg0; // @[FP_inverter.scala 20:42]
  reg [7:0] in2ExpReg1; // @[FP_inverter.scala 22:35]
  reg  in2SignReg1; // @[FP_inverter.scala 24:42]
  reg [7:0] in2ExpReg2; // @[FP_inverter.scala 27:35]
  reg  in2SignReg2; // @[FP_inverter.scala 29:42]
  reg [7:0] in2ExpReg3; // @[FP_inverter.scala 32:35]
  reg  in2SignReg3; // @[FP_inverter.scala 34:42]
  reg [23:0] invMant; // @[FP_inverter.scala 37:42]
  wire [23:0] _T_3 = inverter_io_out; // @[FP_inverter.scala 38:67]
  wire [7:0] negExpTmp = 8'hfe - in2ExpReg3; // @[FP_inverter.scala 41:35]
  wire [7:0] _T_7 = negExpTmp - 8'h1; // @[FP_inverter.scala 42:71]
  wire [7:0] negExp = invMant == 24'h0 ? negExpTmp : _T_7; // @[FP_inverter.scala 42:32]
  wire [22:0] lo = invMant[23:1]; // @[FP_inverter.scala 43:77]
  wire [8:0] hi = {in2SignReg3,negExp}; // @[Cat.scala 30:58]
  fpInverter inverter ( // @[FP_inverter.scala 14:29]
    .clock(inverter_clock),
    .reset(inverter_reset),
    .io_in1(inverter_io_in1),
    .io_out(inverter_io_out)
  );
  assign io_out = {hi,lo}; // @[Cat.scala 30:58]
  assign inverter_clock = clock;
  assign inverter_reset = reset;
  assign inverter_io_in1 = io_in1[22:0]; // @[FP_inverter.scala 16:30]
  always @(posedge clock) begin
    if (reset) begin // @[FP_inverter.scala 18:42]
      in2ExpReg0 <= 8'h0; // @[FP_inverter.scala 18:42]
    end else begin
      in2ExpReg0 <= io_in1[30:23]; // @[FP_inverter.scala 19:44]
    end
    if (reset) begin // @[FP_inverter.scala 20:42]
      in2SignReg0 <= 1'h0; // @[FP_inverter.scala 20:42]
    end else begin
      in2SignReg0 <= io_in1[31]; // @[FP_inverter.scala 21:43]
    end
    if (reset) begin // @[FP_inverter.scala 22:35]
      in2ExpReg1 <= 8'h0; // @[FP_inverter.scala 22:35]
    end else begin
      in2ExpReg1 <= in2ExpReg0; // @[FP_inverter.scala 23:43]
    end
    if (reset) begin // @[FP_inverter.scala 24:42]
      in2SignReg1 <= 1'h0; // @[FP_inverter.scala 24:42]
    end else begin
      in2SignReg1 <= in2SignReg0; // @[FP_inverter.scala 25:43]
    end
    if (reset) begin // @[FP_inverter.scala 27:35]
      in2ExpReg2 <= 8'h0; // @[FP_inverter.scala 27:35]
    end else begin
      in2ExpReg2 <= in2ExpReg1; // @[FP_inverter.scala 28:43]
    end
    if (reset) begin // @[FP_inverter.scala 29:42]
      in2SignReg2 <= 1'h0; // @[FP_inverter.scala 29:42]
    end else begin
      in2SignReg2 <= in2SignReg1; // @[FP_inverter.scala 30:43]
    end
    if (reset) begin // @[FP_inverter.scala 32:35]
      in2ExpReg3 <= 8'h0; // @[FP_inverter.scala 32:35]
    end else begin
      in2ExpReg3 <= in2ExpReg2; // @[FP_inverter.scala 33:43]
    end
    if (reset) begin // @[FP_inverter.scala 34:42]
      in2SignReg3 <= 1'h0; // @[FP_inverter.scala 34:42]
    end else begin
      in2SignReg3 <= in2SignReg2; // @[FP_inverter.scala 35:43]
    end
    if (reset) begin // @[FP_inverter.scala 37:42]
      invMant <= 24'h0; // @[FP_inverter.scala 37:42]
    end else begin
      invMant <= _T_3; // @[FP_inverter.scala 38:49]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  in2ExpReg0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  in2SignReg0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  in2ExpReg1 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  in2SignReg1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  in2ExpReg2 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  in2SignReg2 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  in2ExpReg3 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  in2SignReg3 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  invMant = _RAND_8[23:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Schedule_unit(
  input         clock,
  input         reset,
  input  [31:0] io_invDz_div,
  input         io_valid_in,
  input  [31:0] io_v11_x,
  input  [31:0] io_v11_y,
  input  [31:0] io_v11_z,
  input  [31:0] io_v11_w,
  input  [31:0] io_v22_x,
  input  [31:0] io_v22_y,
  input  [31:0] io_v22_z,
  input  [31:0] io_v22_w,
  input  [31:0] io_ray_in,
  input  [31:0] io_Oz,
  input  [31:0] io_ray_o_in_x,
  input  [31:0] io_ray_o_in_y,
  input  [31:0] io_ray_o_in_z,
  input  [31:0] io_ray_d_in_x,
  input  [31:0] io_ray_d_in_y,
  input  [31:0] io_ray_d_in_z,
  input  [31:0] io_node_id_in,
  input  [31:0] io_hitT_in,
  input         io_break_in,
  input         io_RAY_AABB_1,
  input         io_RAY_AABB_2,
  output [31:0] io_fdiv_out,
  output        io_valid_out,
  output [31:0] io_v11_out_x,
  output [31:0] io_v11_out_y,
  output [31:0] io_v11_out_z,
  output [31:0] io_v11_out_w,
  output [31:0] io_v22_out_x,
  output [31:0] io_v22_out_y,
  output [31:0] io_v22_out_z,
  output [31:0] io_v22_out_w,
  output [31:0] io_ray_out,
  output [31:0] io_Oz_out,
  output [31:0] io_ray_o_out_x,
  output [31:0] io_ray_o_out_y,
  output [31:0] io_ray_o_out_z,
  output [31:0] io_ray_d_out_x,
  output [31:0] io_ray_d_out_y,
  output [31:0] io_ray_d_out_z,
  output [31:0] io_node_id_out,
  output [31:0] io_hitT_out,
  output [31:0] io_counter_fdiv,
  output        io_break_out,
  output        io_RAY_AABB_1_out,
  output        io_RAY_AABB_2_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [95:0] _RAND_4;
  reg [95:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [127:0] _RAND_12;
  reg [127:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [95:0] _RAND_16;
  reg [95:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [127:0] _RAND_24;
  reg [127:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [95:0] _RAND_28;
  reg [95:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [127:0] _RAND_36;
  reg [127:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [95:0] _RAND_40;
  reg [95:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [63:0] _RAND_48;
`endif // RANDOMIZE_REG_INIT
  wire  FP_inverter_clock; // @[Schedule_unit_1.scala 39:39]
  wire  FP_inverter_reset; // @[Schedule_unit_1.scala 39:39]
  wire [31:0] FP_inverter_io_in1; // @[Schedule_unit_1.scala 39:39]
  wire [31:0] FP_inverter_io_out; // @[Schedule_unit_1.scala 39:39]
  reg [127:0] v11_temp_1; // @[Schedule_unit_1.scala 44:38]
  reg [127:0] v22_temp_1; // @[Schedule_unit_1.scala 45:42]
  reg [31:0] ray_temp_1; // @[Schedule_unit_1.scala 46:43]
  reg [31:0] Oz_temp_1; // @[Schedule_unit_1.scala 47:43]
  reg [95:0] ray_o_temp_1; // @[Schedule_unit_1.scala 48:40]
  reg [95:0] ray_d_temp_1; // @[Schedule_unit_1.scala 49:40]
  reg [31:0] node_id_temp_1; // @[Schedule_unit_1.scala 50:37]
  reg [31:0] hitT_temp_1; // @[Schedule_unit_1.scala 51:43]
  reg  inValid_1; // @[Schedule_unit_1.scala 52:61]
  reg  break_1; // @[Schedule_unit_1.scala 53:45]
  reg  ray_aabb_1; // @[Schedule_unit_1.scala 54:46]
  reg  ray_aabb_2; // @[Schedule_unit_1.scala 55:46]
  wire [127:0] _T = {io_v11_w,io_v11_z,io_v11_y,io_v11_x}; // @[Cat.scala 30:58]
  wire [127:0] _T_1 = {io_v22_w,io_v22_z,io_v22_y,io_v22_x}; // @[Cat.scala 30:58]
  wire [95:0] _T_2 = {io_ray_o_in_z,io_ray_o_in_y,io_ray_o_in_x}; // @[Cat.scala 30:58]
  wire [95:0] _T_3 = {io_ray_d_in_z,io_ray_d_in_y,io_ray_d_in_x}; // @[Cat.scala 30:58]
  reg [127:0] v11_temp_2; // @[Schedule_unit_1.scala 70:42]
  reg [127:0] v22_temp_2; // @[Schedule_unit_1.scala 71:42]
  reg [31:0] ray_temp_2; // @[Schedule_unit_1.scala 72:43]
  reg [31:0] Oz_temp_2; // @[Schedule_unit_1.scala 73:43]
  reg [95:0] ray_o_temp_2; // @[Schedule_unit_1.scala 74:40]
  reg [95:0] ray_d_temp_2; // @[Schedule_unit_1.scala 75:40]
  reg [31:0] node_id_temp_2; // @[Schedule_unit_1.scala 76:37]
  reg [31:0] hitT_temp_2; // @[Schedule_unit_1.scala 77:43]
  reg  inValid_2; // @[Schedule_unit_1.scala 78:61]
  reg  break_2; // @[Schedule_unit_1.scala 79:45]
  reg  ray_aabb_1_2; // @[Schedule_unit_1.scala 80:43]
  reg  ray_aabb_2_2; // @[Schedule_unit_1.scala 81:43]
  reg [127:0] v11_temp_3; // @[Schedule_unit_1.scala 96:42]
  reg [127:0] v22_temp_3; // @[Schedule_unit_1.scala 97:42]
  reg [31:0] ray_temp_3; // @[Schedule_unit_1.scala 98:43]
  reg [31:0] Oz_temp_3; // @[Schedule_unit_1.scala 99:43]
  reg [95:0] ray_o_temp_3; // @[Schedule_unit_1.scala 100:40]
  reg [95:0] ray_d_temp_3; // @[Schedule_unit_1.scala 101:40]
  reg [31:0] node_id_temp_3; // @[Schedule_unit_1.scala 102:37]
  reg [31:0] hitT_temp_3; // @[Schedule_unit_1.scala 103:43]
  reg  inValid_3; // @[Schedule_unit_1.scala 104:61]
  reg  break_3; // @[Schedule_unit_1.scala 105:45]
  reg  ray_aabb_1_3; // @[Schedule_unit_1.scala 106:43]
  reg  ray_aabb_2_3; // @[Schedule_unit_1.scala 107:43]
  reg [127:0] v11_temp_4; // @[Schedule_unit_1.scala 121:38]
  reg [127:0] v22_temp_4; // @[Schedule_unit_1.scala 122:42]
  reg [31:0] ray_temp_4; // @[Schedule_unit_1.scala 123:43]
  reg [31:0] Oz_temp_4; // @[Schedule_unit_1.scala 124:43]
  reg [95:0] ray_o_temp_4; // @[Schedule_unit_1.scala 125:40]
  reg [95:0] ray_d_temp_4; // @[Schedule_unit_1.scala 126:40]
  reg [31:0] node_id_temp_4; // @[Schedule_unit_1.scala 127:37]
  reg [31:0] hitT_temp_4; // @[Schedule_unit_1.scala 128:43]
  reg  inValid_4; // @[Schedule_unit_1.scala 129:61]
  reg  break_4; // @[Schedule_unit_1.scala 130:45]
  reg  ray_aabb_1_4; // @[Schedule_unit_1.scala 131:43]
  reg  ray_aabb_2_4; // @[Schedule_unit_1.scala 132:43]
  reg [63:0] count; // @[Schedule_unit_1.scala 171:46]
  wire [63:0] _T_19 = count + 64'h1; // @[Schedule_unit_1.scala 191:26]
  fp_inverter FP_inverter ( // @[Schedule_unit_1.scala 39:39]
    .clock(FP_inverter_clock),
    .reset(FP_inverter_reset),
    .io_in1(FP_inverter_io_in1),
    .io_out(FP_inverter_io_out)
  );
  assign io_fdiv_out = FP_inverter_io_out; // @[Schedule_unit_1.scala 42:45]
  assign io_valid_out = inValid_4; // @[Schedule_unit_1.scala 147:65]
  assign io_v11_out_x = v11_temp_4[31:0]; // @[Schedule_unit_1.scala 148:61]
  assign io_v11_out_y = v11_temp_4[63:32]; // @[Schedule_unit_1.scala 149:61]
  assign io_v11_out_z = v11_temp_4[95:64]; // @[Schedule_unit_1.scala 150:61]
  assign io_v11_out_w = v11_temp_4[127:96]; // @[Schedule_unit_1.scala 151:60]
  assign io_v22_out_x = v22_temp_4[31:0]; // @[Schedule_unit_1.scala 152:61]
  assign io_v22_out_y = v22_temp_4[63:32]; // @[Schedule_unit_1.scala 153:61]
  assign io_v22_out_z = v22_temp_4[95:64]; // @[Schedule_unit_1.scala 154:61]
  assign io_v22_out_w = v22_temp_4[127:96]; // @[Schedule_unit_1.scala 155:59]
  assign io_ray_out = ray_temp_4; // @[Schedule_unit_1.scala 157:50]
  assign io_Oz_out = Oz_temp_4; // @[Schedule_unit_1.scala 158:50]
  assign io_ray_o_out_x = ray_o_temp_4[31:0]; // @[Schedule_unit_1.scala 159:60]
  assign io_ray_o_out_y = ray_o_temp_4[63:32]; // @[Schedule_unit_1.scala 160:60]
  assign io_ray_o_out_z = ray_o_temp_4[95:64]; // @[Schedule_unit_1.scala 161:60]
  assign io_ray_d_out_x = ray_d_temp_4[31:0]; // @[Schedule_unit_1.scala 162:60]
  assign io_ray_d_out_y = ray_d_temp_4[63:32]; // @[Schedule_unit_1.scala 163:60]
  assign io_ray_d_out_z = ray_d_temp_4[95:64]; // @[Schedule_unit_1.scala 164:60]
  assign io_node_id_out = node_id_temp_4; // @[Schedule_unit_1.scala 165:59]
  assign io_hitT_out = hitT_temp_4; // @[Schedule_unit_1.scala 166:73]
  assign io_counter_fdiv = count[31:0]; // @[Schedule_unit_1.scala 196:21]
  assign io_break_out = break_4; // @[Schedule_unit_1.scala 167:42]
  assign io_RAY_AABB_1_out = ray_aabb_1_4; // @[Schedule_unit_1.scala 168:33]
  assign io_RAY_AABB_2_out = ray_aabb_2_4; // @[Schedule_unit_1.scala 169:33]
  assign FP_inverter_clock = clock;
  assign FP_inverter_reset = reset;
  assign FP_inverter_io_in1 = io_invDz_div; // @[Schedule_unit_1.scala 41:37]
  always @(posedge clock) begin
    if (reset) begin // @[Schedule_unit_1.scala 44:38]
      v11_temp_1 <= 128'h0; // @[Schedule_unit_1.scala 44:38]
    end else begin
      v11_temp_1 <= _T; // @[Schedule_unit_1.scala 57:48]
    end
    if (reset) begin // @[Schedule_unit_1.scala 45:42]
      v22_temp_1 <= 128'h0; // @[Schedule_unit_1.scala 45:42]
    end else begin
      v22_temp_1 <= _T_1; // @[Schedule_unit_1.scala 58:48]
    end
    if (reset) begin // @[Schedule_unit_1.scala 46:43]
      ray_temp_1 <= 32'h0; // @[Schedule_unit_1.scala 46:43]
    end else begin
      ray_temp_1 <= io_ray_in; // @[Schedule_unit_1.scala 59:49]
    end
    if (reset) begin // @[Schedule_unit_1.scala 47:43]
      Oz_temp_1 <= 32'h0; // @[Schedule_unit_1.scala 47:43]
    end else begin
      Oz_temp_1 <= io_Oz; // @[Schedule_unit_1.scala 60:49]
    end
    if (reset) begin // @[Schedule_unit_1.scala 48:40]
      ray_o_temp_1 <= 96'h0; // @[Schedule_unit_1.scala 48:40]
    end else begin
      ray_o_temp_1 <= _T_2; // @[Schedule_unit_1.scala 61:46]
    end
    if (reset) begin // @[Schedule_unit_1.scala 49:40]
      ray_d_temp_1 <= 96'h0; // @[Schedule_unit_1.scala 49:40]
    end else begin
      ray_d_temp_1 <= _T_3; // @[Schedule_unit_1.scala 62:46]
    end
    if (reset) begin // @[Schedule_unit_1.scala 50:37]
      node_id_temp_1 <= 32'sh0; // @[Schedule_unit_1.scala 50:37]
    end else begin
      node_id_temp_1 <= io_node_id_in; // @[Schedule_unit_1.scala 63:43]
    end
    if (reset) begin // @[Schedule_unit_1.scala 51:43]
      hitT_temp_1 <= 32'h0; // @[Schedule_unit_1.scala 51:43]
    end else begin
      hitT_temp_1 <= io_hitT_in; // @[Schedule_unit_1.scala 64:49]
    end
    if (reset) begin // @[Schedule_unit_1.scala 52:61]
      inValid_1 <= 1'h0; // @[Schedule_unit_1.scala 52:61]
    end else begin
      inValid_1 <= io_valid_in; // @[Schedule_unit_1.scala 65:50]
    end
    if (reset) begin // @[Schedule_unit_1.scala 53:45]
      break_1 <= 1'h0; // @[Schedule_unit_1.scala 53:45]
    end else begin
      break_1 <= io_break_in; // @[Schedule_unit_1.scala 66:51]
    end
    if (reset) begin // @[Schedule_unit_1.scala 54:46]
      ray_aabb_1 <= 1'h0; // @[Schedule_unit_1.scala 54:46]
    end else begin
      ray_aabb_1 <= io_RAY_AABB_1; // @[Schedule_unit_1.scala 67:40]
    end
    if (reset) begin // @[Schedule_unit_1.scala 55:46]
      ray_aabb_2 <= 1'h0; // @[Schedule_unit_1.scala 55:46]
    end else begin
      ray_aabb_2 <= io_RAY_AABB_2; // @[Schedule_unit_1.scala 68:40]
    end
    if (reset) begin // @[Schedule_unit_1.scala 70:42]
      v11_temp_2 <= 128'h0; // @[Schedule_unit_1.scala 70:42]
    end else begin
      v11_temp_2 <= v11_temp_1; // @[Schedule_unit_1.scala 83:57]
    end
    if (reset) begin // @[Schedule_unit_1.scala 71:42]
      v22_temp_2 <= 128'h0; // @[Schedule_unit_1.scala 71:42]
    end else begin
      v22_temp_2 <= v22_temp_1; // @[Schedule_unit_1.scala 84:57]
    end
    if (reset) begin // @[Schedule_unit_1.scala 72:43]
      ray_temp_2 <= 32'h0; // @[Schedule_unit_1.scala 72:43]
    end else begin
      ray_temp_2 <= ray_temp_1; // @[Schedule_unit_1.scala 85:58]
    end
    if (reset) begin // @[Schedule_unit_1.scala 73:43]
      Oz_temp_2 <= 32'h0; // @[Schedule_unit_1.scala 73:43]
    end else begin
      Oz_temp_2 <= Oz_temp_1; // @[Schedule_unit_1.scala 86:54]
    end
    if (reset) begin // @[Schedule_unit_1.scala 74:40]
      ray_o_temp_2 <= 96'h0; // @[Schedule_unit_1.scala 74:40]
    end else begin
      ray_o_temp_2 <= ray_o_temp_1; // @[Schedule_unit_1.scala 87:39]
    end
    if (reset) begin // @[Schedule_unit_1.scala 75:40]
      ray_d_temp_2 <= 96'h0; // @[Schedule_unit_1.scala 75:40]
    end else begin
      ray_d_temp_2 <= ray_d_temp_1; // @[Schedule_unit_1.scala 88:39]
    end
    if (reset) begin // @[Schedule_unit_1.scala 76:37]
      node_id_temp_2 <= 32'sh0; // @[Schedule_unit_1.scala 76:37]
    end else begin
      node_id_temp_2 <= node_id_temp_1; // @[Schedule_unit_1.scala 89:35]
    end
    if (reset) begin // @[Schedule_unit_1.scala 77:43]
      hitT_temp_2 <= 32'h0; // @[Schedule_unit_1.scala 77:43]
    end else begin
      hitT_temp_2 <= hitT_temp_1; // @[Schedule_unit_1.scala 90:57]
    end
    if (reset) begin // @[Schedule_unit_1.scala 78:61]
      inValid_2 <= 1'h0; // @[Schedule_unit_1.scala 78:61]
    end else begin
      inValid_2 <= inValid_1; // @[Schedule_unit_1.scala 91:66]
    end
    if (reset) begin // @[Schedule_unit_1.scala 79:45]
      break_2 <= 1'h0; // @[Schedule_unit_1.scala 79:45]
    end else begin
      break_2 <= break_1; // @[Schedule_unit_1.scala 92:39]
    end
    if (reset) begin // @[Schedule_unit_1.scala 80:43]
      ray_aabb_1_2 <= 1'h0; // @[Schedule_unit_1.scala 80:43]
    end else begin
      ray_aabb_1_2 <= ray_aabb_1; // @[Schedule_unit_1.scala 93:37]
    end
    if (reset) begin // @[Schedule_unit_1.scala 81:43]
      ray_aabb_2_2 <= 1'h0; // @[Schedule_unit_1.scala 81:43]
    end else begin
      ray_aabb_2_2 <= ray_aabb_2; // @[Schedule_unit_1.scala 94:37]
    end
    if (reset) begin // @[Schedule_unit_1.scala 96:42]
      v11_temp_3 <= 128'h0; // @[Schedule_unit_1.scala 96:42]
    end else begin
      v11_temp_3 <= v11_temp_2; // @[Schedule_unit_1.scala 109:57]
    end
    if (reset) begin // @[Schedule_unit_1.scala 97:42]
      v22_temp_3 <= 128'h0; // @[Schedule_unit_1.scala 97:42]
    end else begin
      v22_temp_3 <= v22_temp_2; // @[Schedule_unit_1.scala 110:57]
    end
    if (reset) begin // @[Schedule_unit_1.scala 98:43]
      ray_temp_3 <= 32'h0; // @[Schedule_unit_1.scala 98:43]
    end else begin
      ray_temp_3 <= ray_temp_2; // @[Schedule_unit_1.scala 111:58]
    end
    if (reset) begin // @[Schedule_unit_1.scala 99:43]
      Oz_temp_3 <= 32'h0; // @[Schedule_unit_1.scala 99:43]
    end else begin
      Oz_temp_3 <= Oz_temp_2; // @[Schedule_unit_1.scala 112:54]
    end
    if (reset) begin // @[Schedule_unit_1.scala 100:40]
      ray_o_temp_3 <= 96'h0; // @[Schedule_unit_1.scala 100:40]
    end else begin
      ray_o_temp_3 <= ray_o_temp_2; // @[Schedule_unit_1.scala 113:39]
    end
    if (reset) begin // @[Schedule_unit_1.scala 101:40]
      ray_d_temp_3 <= 96'h0; // @[Schedule_unit_1.scala 101:40]
    end else begin
      ray_d_temp_3 <= ray_d_temp_2; // @[Schedule_unit_1.scala 114:39]
    end
    if (reset) begin // @[Schedule_unit_1.scala 102:37]
      node_id_temp_3 <= 32'sh0; // @[Schedule_unit_1.scala 102:37]
    end else begin
      node_id_temp_3 <= node_id_temp_2; // @[Schedule_unit_1.scala 115:35]
    end
    if (reset) begin // @[Schedule_unit_1.scala 103:43]
      hitT_temp_3 <= 32'h0; // @[Schedule_unit_1.scala 103:43]
    end else begin
      hitT_temp_3 <= hitT_temp_2; // @[Schedule_unit_1.scala 116:49]
    end
    if (reset) begin // @[Schedule_unit_1.scala 104:61]
      inValid_3 <= 1'h0; // @[Schedule_unit_1.scala 104:61]
    end else begin
      inValid_3 <= inValid_2; // @[Schedule_unit_1.scala 117:66]
    end
    if (reset) begin // @[Schedule_unit_1.scala 105:45]
      break_3 <= 1'h0; // @[Schedule_unit_1.scala 105:45]
    end else begin
      break_3 <= break_2; // @[Schedule_unit_1.scala 118:39]
    end
    if (reset) begin // @[Schedule_unit_1.scala 106:43]
      ray_aabb_1_3 <= 1'h0; // @[Schedule_unit_1.scala 106:43]
    end else begin
      ray_aabb_1_3 <= ray_aabb_1_2; // @[Schedule_unit_1.scala 119:37]
    end
    if (reset) begin // @[Schedule_unit_1.scala 107:43]
      ray_aabb_2_3 <= 1'h0; // @[Schedule_unit_1.scala 107:43]
    end else begin
      ray_aabb_2_3 <= ray_aabb_2_2; // @[Schedule_unit_1.scala 120:37]
    end
    if (reset) begin // @[Schedule_unit_1.scala 121:38]
      v11_temp_4 <= 128'h0; // @[Schedule_unit_1.scala 121:38]
    end else begin
      v11_temp_4 <= v11_temp_3; // @[Schedule_unit_1.scala 134:57]
    end
    if (reset) begin // @[Schedule_unit_1.scala 122:42]
      v22_temp_4 <= 128'h0; // @[Schedule_unit_1.scala 122:42]
    end else begin
      v22_temp_4 <= v22_temp_3; // @[Schedule_unit_1.scala 135:57]
    end
    if (reset) begin // @[Schedule_unit_1.scala 123:43]
      ray_temp_4 <= 32'h0; // @[Schedule_unit_1.scala 123:43]
    end else begin
      ray_temp_4 <= ray_temp_3; // @[Schedule_unit_1.scala 136:58]
    end
    if (reset) begin // @[Schedule_unit_1.scala 124:43]
      Oz_temp_4 <= 32'h0; // @[Schedule_unit_1.scala 124:43]
    end else begin
      Oz_temp_4 <= Oz_temp_3; // @[Schedule_unit_1.scala 137:54]
    end
    if (reset) begin // @[Schedule_unit_1.scala 125:40]
      ray_o_temp_4 <= 96'h0; // @[Schedule_unit_1.scala 125:40]
    end else begin
      ray_o_temp_4 <= ray_o_temp_3; // @[Schedule_unit_1.scala 138:39]
    end
    if (reset) begin // @[Schedule_unit_1.scala 126:40]
      ray_d_temp_4 <= 96'h0; // @[Schedule_unit_1.scala 126:40]
    end else begin
      ray_d_temp_4 <= ray_d_temp_3; // @[Schedule_unit_1.scala 139:39]
    end
    if (reset) begin // @[Schedule_unit_1.scala 127:37]
      node_id_temp_4 <= 32'sh0; // @[Schedule_unit_1.scala 127:37]
    end else begin
      node_id_temp_4 <= node_id_temp_3; // @[Schedule_unit_1.scala 140:35]
    end
    if (reset) begin // @[Schedule_unit_1.scala 128:43]
      hitT_temp_4 <= 32'h0; // @[Schedule_unit_1.scala 128:43]
    end else begin
      hitT_temp_4 <= hitT_temp_3; // @[Schedule_unit_1.scala 141:49]
    end
    if (reset) begin // @[Schedule_unit_1.scala 129:61]
      inValid_4 <= 1'h0; // @[Schedule_unit_1.scala 129:61]
    end else begin
      inValid_4 <= inValid_3; // @[Schedule_unit_1.scala 142:66]
    end
    if (reset) begin // @[Schedule_unit_1.scala 130:45]
      break_4 <= 1'h0; // @[Schedule_unit_1.scala 130:45]
    end else begin
      break_4 <= break_3; // @[Schedule_unit_1.scala 143:39]
    end
    if (reset) begin // @[Schedule_unit_1.scala 131:43]
      ray_aabb_1_4 <= 1'h0; // @[Schedule_unit_1.scala 131:43]
    end else begin
      ray_aabb_1_4 <= ray_aabb_1_3; // @[Schedule_unit_1.scala 144:37]
    end
    if (reset) begin // @[Schedule_unit_1.scala 132:43]
      ray_aabb_2_4 <= 1'h0; // @[Schedule_unit_1.scala 132:43]
    end else begin
      ray_aabb_2_4 <= ray_aabb_2_3; // @[Schedule_unit_1.scala 145:37]
    end
    if (reset) begin // @[Schedule_unit_1.scala 171:46]
      count <= 64'h0; // @[Schedule_unit_1.scala 171:46]
    end else if (io_valid_in) begin // @[Schedule_unit_1.scala 190:22]
      count <= _T_19; // @[Schedule_unit_1.scala 191:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  v11_temp_1 = _RAND_0[127:0];
  _RAND_1 = {4{`RANDOM}};
  v22_temp_1 = _RAND_1[127:0];
  _RAND_2 = {1{`RANDOM}};
  ray_temp_1 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  Oz_temp_1 = _RAND_3[31:0];
  _RAND_4 = {3{`RANDOM}};
  ray_o_temp_1 = _RAND_4[95:0];
  _RAND_5 = {3{`RANDOM}};
  ray_d_temp_1 = _RAND_5[95:0];
  _RAND_6 = {1{`RANDOM}};
  node_id_temp_1 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  hitT_temp_1 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  inValid_1 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  break_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  ray_aabb_1 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ray_aabb_2 = _RAND_11[0:0];
  _RAND_12 = {4{`RANDOM}};
  v11_temp_2 = _RAND_12[127:0];
  _RAND_13 = {4{`RANDOM}};
  v22_temp_2 = _RAND_13[127:0];
  _RAND_14 = {1{`RANDOM}};
  ray_temp_2 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  Oz_temp_2 = _RAND_15[31:0];
  _RAND_16 = {3{`RANDOM}};
  ray_o_temp_2 = _RAND_16[95:0];
  _RAND_17 = {3{`RANDOM}};
  ray_d_temp_2 = _RAND_17[95:0];
  _RAND_18 = {1{`RANDOM}};
  node_id_temp_2 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  hitT_temp_2 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  inValid_2 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  break_2 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  ray_aabb_1_2 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  ray_aabb_2_2 = _RAND_23[0:0];
  _RAND_24 = {4{`RANDOM}};
  v11_temp_3 = _RAND_24[127:0];
  _RAND_25 = {4{`RANDOM}};
  v22_temp_3 = _RAND_25[127:0];
  _RAND_26 = {1{`RANDOM}};
  ray_temp_3 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  Oz_temp_3 = _RAND_27[31:0];
  _RAND_28 = {3{`RANDOM}};
  ray_o_temp_3 = _RAND_28[95:0];
  _RAND_29 = {3{`RANDOM}};
  ray_d_temp_3 = _RAND_29[95:0];
  _RAND_30 = {1{`RANDOM}};
  node_id_temp_3 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  hitT_temp_3 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  inValid_3 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  break_3 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  ray_aabb_1_3 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  ray_aabb_2_3 = _RAND_35[0:0];
  _RAND_36 = {4{`RANDOM}};
  v11_temp_4 = _RAND_36[127:0];
  _RAND_37 = {4{`RANDOM}};
  v22_temp_4 = _RAND_37[127:0];
  _RAND_38 = {1{`RANDOM}};
  ray_temp_4 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  Oz_temp_4 = _RAND_39[31:0];
  _RAND_40 = {3{`RANDOM}};
  ray_o_temp_4 = _RAND_40[95:0];
  _RAND_41 = {3{`RANDOM}};
  ray_d_temp_4 = _RAND_41[95:0];
  _RAND_42 = {1{`RANDOM}};
  node_id_temp_4 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  hitT_temp_4 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  inValid_4 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  break_4 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  ray_aabb_1_4 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  ray_aabb_2_4 = _RAND_47[0:0];
  _RAND_48 = {2{`RANDOM}};
  count = _RAND_48[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IST1(
  input         clock,
  input         reset,
  input         io_enable_IST1,
  input  [31:0] io_nodeid_leaf_1,
  input  [31:0] io_rayid_leaf_1,
  input  [31:0] io_hiT_in,
  input  [31:0] io_Oz,
  input  [31:0] io_invDz,
  input  [31:0] io_v11_in_x,
  input  [31:0] io_v11_in_y,
  input  [31:0] io_v11_in_z,
  input  [31:0] io_v11_in_w,
  input  [31:0] io_v22_in_x,
  input  [31:0] io_v22_in_y,
  input  [31:0] io_v22_in_z,
  input  [31:0] io_v22_in_w,
  input  [31:0] io_ray_o_in_x,
  input  [31:0] io_ray_o_in_y,
  input  [31:0] io_ray_o_in_z,
  input  [31:0] io_ray_d_in_x,
  input  [31:0] io_ray_d_in_y,
  input  [31:0] io_ray_d_in_z,
  input         io_break_in,
  input         io_RAY_AABB_1,
  input         io_RAY_AABB_2,
  output [31:0] io_nodeid_ist1_out,
  output [31:0] io_rayid_ist1_out,
  output [31:0] io_hiT_out,
  output [31:0] io_t,
  output        io_pop_1,
  output [31:0] io_v11_out_x,
  output [31:0] io_v11_out_y,
  output [31:0] io_v11_out_z,
  output [31:0] io_v11_out_w,
  output [31:0] io_v22_out_x,
  output [31:0] io_v22_out_y,
  output [31:0] io_v22_out_z,
  output [31:0] io_v22_out_w,
  output [31:0] io_ray_o_out_x,
  output [31:0] io_ray_o_out_y,
  output [31:0] io_ray_o_out_z,
  output [31:0] io_ray_d_out_x,
  output [31:0] io_ray_d_out_y,
  output [31:0] io_ray_d_out_z,
  output        io_enable_IST2,
  output        io_break_out,
  output        io_break_ist1,
  output        io_RAY_AABB_1_out,
  output        io_RAY_AABB_2_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [127:0] _RAND_5;
  reg [127:0] _RAND_6;
  reg [95:0] _RAND_7;
  reg [95:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [127:0] _RAND_16;
  reg [127:0] _RAND_17;
  reg [95:0] _RAND_18;
  reg [95:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [127:0] _RAND_29;
  reg [127:0] _RAND_30;
  reg [95:0] _RAND_31;
  reg [95:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
`endif // RANDOMIZE_REG_INIT
  wire  FMUL_6_clock; // @[IST1.scala 69:24]
  wire  FMUL_6_reset; // @[IST1.scala 69:24]
  wire [31:0] FMUL_6_io_a; // @[IST1.scala 69:24]
  wire [31:0] FMUL_6_io_b; // @[IST1.scala 69:24]
  wire [31:0] FMUL_6_io_out; // @[IST1.scala 69:24]
  wire [31:0] FCMP_21_io_a; // @[IST1.scala 131:25]
  wire [31:0] FCMP_21_io_b; // @[IST1.scala 131:25]
  wire  FCMP_21_io_actual_out; // @[IST1.scala 131:25]
  wire [31:0] FCMP_22_io_a; // @[IST1.scala 141:25]
  wire [31:0] FCMP_22_io_b; // @[IST1.scala 141:25]
  wire  FCMP_22_io_actual_out; // @[IST1.scala 141:25]
  reg  enable_1; // @[IST1.scala 45:52]
  reg [31:0] nodeid_ist1_temp_1; // @[IST1.scala 46:38]
  reg [31:0] rayid_ist1_temp_1; // @[IST1.scala 47:41]
  reg [31:0] hitT_temp_1; // @[IST1.scala 48:47]
  reg [31:0] t_1; // @[IST1.scala 49:59]
  reg [127:0] v11_1; // @[IST1.scala 50:56]
  reg [127:0] v22_1; // @[IST1.scala 51:56]
  reg [95:0] ray_o_in_1; // @[IST1.scala 52:50]
  reg [95:0] ray_d_in_1; // @[IST1.scala 53:50]
  reg  break_1; // @[IST1.scala 54:54]
  reg  ray_aabb_1; // @[IST1.scala 55:46]
  reg  ray_aabb_2; // @[IST1.scala 56:46]
  wire [127:0] _T = {io_v11_in_w,io_v11_in_z,io_v11_in_y,io_v11_in_x}; // @[Cat.scala 30:58]
  wire [127:0] _T_1 = {io_v22_in_w,io_v22_in_z,io_v22_in_y,io_v22_in_x}; // @[Cat.scala 30:58]
  wire [95:0] _T_2 = {io_ray_o_in_z,io_ray_o_in_y,io_ray_o_in_x}; // @[Cat.scala 30:58]
  wire [95:0] _T_3 = {io_ray_d_in_z,io_ray_d_in_y,io_ray_d_in_x}; // @[Cat.scala 30:58]
  reg  mul_enable_1; // @[IST1.scala 78:56]
  reg [31:0] mul_nodeid_ist1_temp_1; // @[IST1.scala 79:42]
  reg [31:0] mul_rayid_ist1_temp_1; // @[IST1.scala 80:45]
  reg [31:0] mul_hitT_temp_1; // @[IST1.scala 81:51]
  reg [127:0] mul_v11_1; // @[IST1.scala 83:60]
  reg [127:0] mul_v22_1; // @[IST1.scala 84:60]
  reg [95:0] mul_ray_o_in_1; // @[IST1.scala 85:54]
  reg [95:0] mul_ray_d_in_1; // @[IST1.scala 86:54]
  reg  mul_break_1; // @[IST1.scala 87:58]
  reg  mul_ray_aabb_1; // @[IST1.scala 88:50]
  reg  mul_ray_aabb_2; // @[IST1.scala 89:50]
  reg [31:0] nodeid_ist1_temp_2; // @[IST1.scala 104:38]
  reg [31:0] rayid_ist1_temp_2; // @[IST1.scala 105:41]
  reg [31:0] hitT_temp_2; // @[IST1.scala 106:47]
  reg [31:0] t_2; // @[IST1.scala 107:59]
  reg  t_min; // @[IST1.scala 108:54]
  reg  t_hitT; // @[IST1.scala 109:55]
  reg [127:0] v11_2; // @[IST1.scala 110:56]
  reg [127:0] v22_2; // @[IST1.scala 111:56]
  reg [95:0] ray_o_in_2; // @[IST1.scala 112:50]
  reg [95:0] ray_d_in_2; // @[IST1.scala 113:50]
  reg  enable_2; // @[IST1.scala 114:50]
  reg  break_2; // @[IST1.scala 115:52]
  reg  ray_aabb_1_2; // @[IST1.scala 116:43]
  reg  ray_aabb_2_2; // @[IST1.scala 117:43]
  wire  _T_4 = FCMP_21_io_actual_out > 1'h0; // @[IST1.scala 136:36]
  wire  _T_5 = FCMP_22_io_actual_out > 1'h0; // @[IST1.scala 146:36]
  wire  _T_20 = t_min & t_hitT; // @[IST1.scala 173:19]
  wire  _T_23 = t_min & t_hitT & enable_2; // @[IST1.scala 173:36]
  wire  _T_24 = ~break_2; // @[IST1.scala 173:64]
  wire  _T_29 = ~_T_20 & enable_2; // @[IST1.scala 178:41]
  wire  _T_31 = ~_T_20 & enable_2 & _T_24; // @[IST1.scala 178:59]
  wire  _T_37 = _T_23 & break_2; // @[IST1.scala 183:59]
  wire  _T_43 = _T_29 & break_2; // @[IST1.scala 188:59]
  wire  _GEN_6 = _T_23 & break_2 ? 1'h0 : _T_43; // @[IST1.scala 183:77 IST1.scala 187:31]
  wire  _GEN_7 = ~_T_20 & enable_2 & _T_24 ? 1'h0 : _T_37; // @[IST1.scala 178:77 IST1.scala 179:28]
  wire  _GEN_9 = ~_T_20 & enable_2 & _T_24 ? 1'h0 : _GEN_6; // @[IST1.scala 178:77 IST1.scala 182:31]
  MY_MUL FMUL_6 ( // @[IST1.scala 69:24]
    .clock(FMUL_6_clock),
    .reset(FMUL_6_reset),
    .io_a(FMUL_6_io_a),
    .io_b(FMUL_6_io_b),
    .io_out(FMUL_6_io_out)
  );
  ValExec_CompareRecF32_lt FCMP_21 ( // @[IST1.scala 131:25]
    .io_a(FCMP_21_io_a),
    .io_b(FCMP_21_io_b),
    .io_actual_out(FCMP_21_io_actual_out)
  );
  ValExec_CompareRecF32_lt FCMP_22 ( // @[IST1.scala 141:25]
    .io_a(FCMP_22_io_a),
    .io_b(FCMP_22_io_b),
    .io_actual_out(FCMP_22_io_actual_out)
  );
  assign io_nodeid_ist1_out = nodeid_ist1_temp_2; // @[IST1.scala 160:39]
  assign io_rayid_ist1_out = rayid_ist1_temp_2; // @[IST1.scala 161:42]
  assign io_hiT_out = hitT_temp_2; // @[IST1.scala 163:49]
  assign io_t = t_2; // @[IST1.scala 162:58]
  assign io_pop_1 = t_min & t_hitT & enable_2 & ~break_2 ? 1'h0 : _T_31; // @[IST1.scala 173:72 IST1.scala 175:35]
  assign io_v11_out_x = v11_2[31:0]; // @[IST1.scala 152:52]
  assign io_v11_out_y = v11_2[63:32]; // @[IST1.scala 153:52]
  assign io_v11_out_z = v11_2[95:64]; // @[IST1.scala 154:52]
  assign io_v11_out_w = v11_2[127:96]; // @[IST1.scala 155:51]
  assign io_v22_out_x = v22_2[31:0]; // @[IST1.scala 156:56]
  assign io_v22_out_y = v22_2[63:32]; // @[IST1.scala 157:56]
  assign io_v22_out_z = v22_2[95:64]; // @[IST1.scala 158:56]
  assign io_v22_out_w = v22_2[127:96]; // @[IST1.scala 159:54]
  assign io_ray_o_out_x = ray_o_in_2[31:0]; // @[IST1.scala 164:58]
  assign io_ray_o_out_y = ray_o_in_2[63:32]; // @[IST1.scala 165:58]
  assign io_ray_o_out_z = ray_o_in_2[95:64]; // @[IST1.scala 166:58]
  assign io_ray_d_out_x = ray_d_in_2[31:0]; // @[IST1.scala 167:58]
  assign io_ray_d_out_y = ray_d_in_2[63:32]; // @[IST1.scala 168:58]
  assign io_ray_d_out_z = ray_d_in_2[95:64]; // @[IST1.scala 169:58]
  assign io_enable_IST2 = t_min & t_hitT & enable_2 & ~break_2 | _GEN_7; // @[IST1.scala 173:72 IST1.scala 174:28]
  assign io_break_out = t_min & t_hitT & enable_2 & ~break_2 ? 1'h0 : _GEN_9; // @[IST1.scala 173:72 IST1.scala 177:31]
  assign io_break_ist1 = break_2; // @[IST1.scala 170:47]
  assign io_RAY_AABB_1_out = ray_aabb_1_2; // @[IST1.scala 171:36]
  assign io_RAY_AABB_2_out = ray_aabb_2_2; // @[IST1.scala 172:36]
  assign FMUL_6_clock = clock;
  assign FMUL_6_reset = reset;
  assign FMUL_6_io_a = io_Oz; // @[IST1.scala 70:21]
  assign FMUL_6_io_b = io_invDz; // @[IST1.scala 71:21]
  assign FCMP_21_io_a = 32'h0; // @[IST1.scala 132:22]
  assign FCMP_21_io_b = t_1; // @[IST1.scala 133:22]
  assign FCMP_22_io_a = t_1; // @[IST1.scala 142:22]
  assign FCMP_22_io_b = mul_hitT_temp_1; // @[IST1.scala 143:22]
  always @(posedge clock) begin
    if (reset) begin // @[IST1.scala 45:52]
      enable_1 <= 1'h0; // @[IST1.scala 45:52]
    end else begin
      enable_1 <= io_enable_IST1; // @[IST1.scala 65:43]
    end
    if (reset) begin // @[IST1.scala 46:38]
      nodeid_ist1_temp_1 <= 32'sh0; // @[IST1.scala 46:38]
    end else begin
      nodeid_ist1_temp_1 <= io_nodeid_leaf_1; // @[IST1.scala 58:29]
    end
    if (reset) begin // @[IST1.scala 47:41]
      rayid_ist1_temp_1 <= 32'h0; // @[IST1.scala 47:41]
    end else begin
      rayid_ist1_temp_1 <= io_rayid_leaf_1; // @[IST1.scala 59:32]
    end
    if (reset) begin // @[IST1.scala 48:47]
      hitT_temp_1 <= 32'h0; // @[IST1.scala 48:47]
    end else begin
      hitT_temp_1 <= io_hiT_in; // @[IST1.scala 60:38]
    end
    if (reset) begin // @[IST1.scala 49:59]
      t_1 <= 32'h0; // @[IST1.scala 49:59]
    end else begin
      t_1 <= FMUL_6_io_out; // @[IST1.scala 76:46]
    end
    if (reset) begin // @[IST1.scala 50:56]
      v11_1 <= 128'h0; // @[IST1.scala 50:56]
    end else begin
      v11_1 <= _T; // @[IST1.scala 61:46]
    end
    if (reset) begin // @[IST1.scala 51:56]
      v22_1 <= 128'h0; // @[IST1.scala 51:56]
    end else begin
      v22_1 <= _T_1; // @[IST1.scala 62:46]
    end
    if (reset) begin // @[IST1.scala 52:50]
      ray_o_in_1 <= 96'h0; // @[IST1.scala 52:50]
    end else begin
      ray_o_in_1 <= _T_2; // @[IST1.scala 63:40]
    end
    if (reset) begin // @[IST1.scala 53:50]
      ray_d_in_1 <= 96'h0; // @[IST1.scala 53:50]
    end else begin
      ray_d_in_1 <= _T_3; // @[IST1.scala 64:40]
    end
    if (reset) begin // @[IST1.scala 54:54]
      break_1 <= 1'h0; // @[IST1.scala 54:54]
    end else begin
      break_1 <= io_break_in; // @[IST1.scala 66:45]
    end
    if (reset) begin // @[IST1.scala 55:46]
      ray_aabb_1 <= 1'h0; // @[IST1.scala 55:46]
    end else begin
      ray_aabb_1 <= io_RAY_AABB_1; // @[IST1.scala 67:40]
    end
    if (reset) begin // @[IST1.scala 56:46]
      ray_aabb_2 <= 1'h0; // @[IST1.scala 56:46]
    end else begin
      ray_aabb_2 <= io_RAY_AABB_2; // @[IST1.scala 68:40]
    end
    if (reset) begin // @[IST1.scala 78:56]
      mul_enable_1 <= 1'h0; // @[IST1.scala 78:56]
    end else begin
      mul_enable_1 <= enable_1; // @[IST1.scala 98:47]
    end
    if (reset) begin // @[IST1.scala 79:42]
      mul_nodeid_ist1_temp_1 <= 32'sh0; // @[IST1.scala 79:42]
    end else begin
      mul_nodeid_ist1_temp_1 <= nodeid_ist1_temp_1; // @[IST1.scala 91:33]
    end
    if (reset) begin // @[IST1.scala 80:45]
      mul_rayid_ist1_temp_1 <= 32'h0; // @[IST1.scala 80:45]
    end else begin
      mul_rayid_ist1_temp_1 <= rayid_ist1_temp_1; // @[IST1.scala 92:36]
    end
    if (reset) begin // @[IST1.scala 81:51]
      mul_hitT_temp_1 <= 32'h0; // @[IST1.scala 81:51]
    end else begin
      mul_hitT_temp_1 <= hitT_temp_1; // @[IST1.scala 93:42]
    end
    if (reset) begin // @[IST1.scala 83:60]
      mul_v11_1 <= 128'h0; // @[IST1.scala 83:60]
    end else begin
      mul_v11_1 <= v11_1; // @[IST1.scala 94:50]
    end
    if (reset) begin // @[IST1.scala 84:60]
      mul_v22_1 <= 128'h0; // @[IST1.scala 84:60]
    end else begin
      mul_v22_1 <= v22_1; // @[IST1.scala 95:50]
    end
    if (reset) begin // @[IST1.scala 85:54]
      mul_ray_o_in_1 <= 96'h0; // @[IST1.scala 85:54]
    end else begin
      mul_ray_o_in_1 <= ray_o_in_1; // @[IST1.scala 96:44]
    end
    if (reset) begin // @[IST1.scala 86:54]
      mul_ray_d_in_1 <= 96'h0; // @[IST1.scala 86:54]
    end else begin
      mul_ray_d_in_1 <= ray_d_in_1; // @[IST1.scala 97:44]
    end
    if (reset) begin // @[IST1.scala 87:58]
      mul_break_1 <= 1'h0; // @[IST1.scala 87:58]
    end else begin
      mul_break_1 <= break_1; // @[IST1.scala 99:49]
    end
    if (reset) begin // @[IST1.scala 88:50]
      mul_ray_aabb_1 <= 1'h0; // @[IST1.scala 88:50]
    end else begin
      mul_ray_aabb_1 <= ray_aabb_1; // @[IST1.scala 100:45]
    end
    if (reset) begin // @[IST1.scala 89:50]
      mul_ray_aabb_2 <= 1'h0; // @[IST1.scala 89:50]
    end else begin
      mul_ray_aabb_2 <= ray_aabb_2; // @[IST1.scala 101:46]
    end
    if (reset) begin // @[IST1.scala 104:38]
      nodeid_ist1_temp_2 <= 32'sh0; // @[IST1.scala 104:38]
    end else begin
      nodeid_ist1_temp_2 <= mul_nodeid_ist1_temp_1; // @[IST1.scala 119:29]
    end
    if (reset) begin // @[IST1.scala 105:41]
      rayid_ist1_temp_2 <= 32'h0; // @[IST1.scala 105:41]
    end else begin
      rayid_ist1_temp_2 <= mul_rayid_ist1_temp_1; // @[IST1.scala 120:32]
    end
    if (reset) begin // @[IST1.scala 106:47]
      hitT_temp_2 <= 32'h0; // @[IST1.scala 106:47]
    end else begin
      hitT_temp_2 <= mul_hitT_temp_1; // @[IST1.scala 121:38]
    end
    if (reset) begin // @[IST1.scala 107:59]
      t_2 <= 32'h0; // @[IST1.scala 107:59]
    end else begin
      t_2 <= t_1; // @[IST1.scala 122:50]
    end
    if (reset) begin // @[IST1.scala 108:54]
      t_min <= 1'h0; // @[IST1.scala 108:54]
    end else begin
      t_min <= _T_4;
    end
    if (reset) begin // @[IST1.scala 109:55]
      t_hitT <= 1'h0; // @[IST1.scala 109:55]
    end else begin
      t_hitT <= _T_5;
    end
    if (reset) begin // @[IST1.scala 110:56]
      v11_2 <= 128'h0; // @[IST1.scala 110:56]
    end else begin
      v11_2 <= mul_v11_1; // @[IST1.scala 123:46]
    end
    if (reset) begin // @[IST1.scala 111:56]
      v22_2 <= 128'h0; // @[IST1.scala 111:56]
    end else begin
      v22_2 <= mul_v22_1; // @[IST1.scala 124:46]
    end
    if (reset) begin // @[IST1.scala 112:50]
      ray_o_in_2 <= 96'h0; // @[IST1.scala 112:50]
    end else begin
      ray_o_in_2 <= mul_ray_o_in_1; // @[IST1.scala 125:40]
    end
    if (reset) begin // @[IST1.scala 113:50]
      ray_d_in_2 <= 96'h0; // @[IST1.scala 113:50]
    end else begin
      ray_d_in_2 <= mul_ray_d_in_1; // @[IST1.scala 126:40]
    end
    if (reset) begin // @[IST1.scala 114:50]
      enable_2 <= 1'h0; // @[IST1.scala 114:50]
    end else begin
      enable_2 <= mul_enable_1; // @[IST1.scala 127:42]
    end
    if (reset) begin // @[IST1.scala 115:52]
      break_2 <= 1'h0; // @[IST1.scala 115:52]
    end else begin
      break_2 <= mul_break_1; // @[IST1.scala 128:44]
    end
    if (reset) begin // @[IST1.scala 116:43]
      ray_aabb_1_2 <= 1'h0; // @[IST1.scala 116:43]
    end else begin
      ray_aabb_1_2 <= mul_ray_aabb_1; // @[IST1.scala 129:37]
    end
    if (reset) begin // @[IST1.scala 117:43]
      ray_aabb_2_2 <= 1'h0; // @[IST1.scala 117:43]
    end else begin
      ray_aabb_2_2 <= mul_ray_aabb_2; // @[IST1.scala 130:37]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_1 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  nodeid_ist1_temp_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  rayid_ist1_temp_1 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  hitT_temp_1 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  t_1 = _RAND_4[31:0];
  _RAND_5 = {4{`RANDOM}};
  v11_1 = _RAND_5[127:0];
  _RAND_6 = {4{`RANDOM}};
  v22_1 = _RAND_6[127:0];
  _RAND_7 = {3{`RANDOM}};
  ray_o_in_1 = _RAND_7[95:0];
  _RAND_8 = {3{`RANDOM}};
  ray_d_in_1 = _RAND_8[95:0];
  _RAND_9 = {1{`RANDOM}};
  break_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  ray_aabb_1 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ray_aabb_2 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  mul_enable_1 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  mul_nodeid_ist1_temp_1 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  mul_rayid_ist1_temp_1 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  mul_hitT_temp_1 = _RAND_15[31:0];
  _RAND_16 = {4{`RANDOM}};
  mul_v11_1 = _RAND_16[127:0];
  _RAND_17 = {4{`RANDOM}};
  mul_v22_1 = _RAND_17[127:0];
  _RAND_18 = {3{`RANDOM}};
  mul_ray_o_in_1 = _RAND_18[95:0];
  _RAND_19 = {3{`RANDOM}};
  mul_ray_d_in_1 = _RAND_19[95:0];
  _RAND_20 = {1{`RANDOM}};
  mul_break_1 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  mul_ray_aabb_1 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  mul_ray_aabb_2 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  nodeid_ist1_temp_2 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  rayid_ist1_temp_2 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  hitT_temp_2 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  t_2 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  t_min = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  t_hitT = _RAND_28[0:0];
  _RAND_29 = {4{`RANDOM}};
  v11_2 = _RAND_29[127:0];
  _RAND_30 = {4{`RANDOM}};
  v22_2 = _RAND_30[127:0];
  _RAND_31 = {3{`RANDOM}};
  ray_o_in_2 = _RAND_31[95:0];
  _RAND_32 = {3{`RANDOM}};
  ray_d_in_2 = _RAND_32[95:0];
  _RAND_33 = {1{`RANDOM}};
  enable_2 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  break_2 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  ray_aabb_1_2 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  ray_aabb_2_2 = _RAND_36[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IST2(
  input         clock,
  input         reset,
  input         io_enable_IST2,
  input  [31:0] io_nodeid_leaf_2,
  input  [31:0] io_rayid_leaf_2,
  input  [31:0] io_hiT_in,
  input  [31:0] io_v11_in_x,
  input  [31:0] io_v11_in_y,
  input  [31:0] io_v11_in_z,
  input  [31:0] io_v11_in_w,
  input  [31:0] io_v22_in_x,
  input  [31:0] io_v22_in_y,
  input  [31:0] io_v22_in_z,
  input  [31:0] io_v22_in_w,
  input  [31:0] io_ray_o_in_x,
  input  [31:0] io_ray_o_in_y,
  input  [31:0] io_ray_o_in_z,
  input  [31:0] io_ray_d_in_x,
  input  [31:0] io_ray_d_in_y,
  input  [31:0] io_ray_d_in_z,
  input  [31:0] io_t,
  input         io_break_in,
  input         io_RAY_AABB_1,
  input         io_RAY_AABB_2,
  output [31:0] io_nodeid_ist2_out,
  output [31:0] io_rayid_ist2_out,
  output [31:0] io_hiT_out,
  output [31:0] io_u,
  output        io_pop_2,
  output [31:0] io_t_out,
  output [31:0] io_v22_out_x,
  output [31:0] io_v22_out_y,
  output [31:0] io_v22_out_z,
  output [31:0] io_v22_out_w,
  output [31:0] io_ray_o_out_x,
  output [31:0] io_ray_o_out_y,
  output [31:0] io_ray_o_out_z,
  output [31:0] io_ray_d_out_x,
  output [31:0] io_ray_d_out_y,
  output [31:0] io_ray_d_out_z,
  output        io_enable_IST3,
  output        io_break_ist2,
  output        io_break_out,
  output        io_RAY_AABB_1_out,
  output        io_RAY_AABB_2_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [127:0] _RAND_10;
  reg [95:0] _RAND_11;
  reg [95:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [127:0] _RAND_21;
  reg [95:0] _RAND_22;
  reg [95:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [127:0] _RAND_32;
  reg [95:0] _RAND_33;
  reg [95:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [127:0] _RAND_49;
  reg [95:0] _RAND_50;
  reg [95:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [127:0] _RAND_60;
  reg [95:0] _RAND_61;
  reg [95:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [127:0] _RAND_73;
  reg [95:0] _RAND_74;
  reg [95:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [127:0] _RAND_85;
  reg [95:0] _RAND_86;
  reg [95:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [127:0] _RAND_96;
  reg [95:0] _RAND_97;
  reg [95:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
`endif // RANDOMIZE_REG_INIT
  wire  FADD_MUL_14_clock; // @[IST2.scala 74:33]
  wire  FADD_MUL_14_reset; // @[IST2.scala 74:33]
  wire [31:0] FADD_MUL_14_io_a; // @[IST2.scala 74:33]
  wire [31:0] FADD_MUL_14_io_b; // @[IST2.scala 74:33]
  wire [31:0] FADD_MUL_14_io_c; // @[IST2.scala 74:33]
  wire [31:0] FADD_MUL_14_io_out; // @[IST2.scala 74:33]
  wire  FMUL_7_clock; // @[IST2.scala 84:24]
  wire  FMUL_7_reset; // @[IST2.scala 84:24]
  wire [31:0] FMUL_7_io_a; // @[IST2.scala 84:24]
  wire [31:0] FMUL_7_io_b; // @[IST2.scala 84:24]
  wire [31:0] FMUL_7_io_out; // @[IST2.scala 84:24]
  wire  FMUL_8_clock; // @[IST2.scala 93:24]
  wire  FMUL_8_reset; // @[IST2.scala 93:24]
  wire [31:0] FMUL_8_io_a; // @[IST2.scala 93:24]
  wire [31:0] FMUL_8_io_b; // @[IST2.scala 93:24]
  wire [31:0] FMUL_8_io_out; // @[IST2.scala 93:24]
  wire  FMUL_9_clock; // @[IST2.scala 102:24]
  wire  FMUL_9_reset; // @[IST2.scala 102:24]
  wire [31:0] FMUL_9_io_a; // @[IST2.scala 102:24]
  wire [31:0] FMUL_9_io_b; // @[IST2.scala 102:24]
  wire [31:0] FMUL_9_io_out; // @[IST2.scala 102:24]
  wire  FMUL_10_clock; // @[IST2.scala 111:25]
  wire  FMUL_10_reset; // @[IST2.scala 111:25]
  wire [31:0] FMUL_10_io_a; // @[IST2.scala 111:25]
  wire [31:0] FMUL_10_io_b; // @[IST2.scala 111:25]
  wire [31:0] FMUL_10_io_out; // @[IST2.scala 111:25]
  wire  FMUL_11_clock; // @[IST2.scala 120:25]
  wire  FMUL_11_reset; // @[IST2.scala 120:25]
  wire [31:0] FMUL_11_io_a; // @[IST2.scala 120:25]
  wire [31:0] FMUL_11_io_b; // @[IST2.scala 120:25]
  wire [31:0] FMUL_11_io_out; // @[IST2.scala 120:25]
  wire  FADD_5_clock; // @[IST2.scala 192:24]
  wire  FADD_5_reset; // @[IST2.scala 192:24]
  wire [31:0] FADD_5_io_a; // @[IST2.scala 192:24]
  wire [31:0] FADD_5_io_b; // @[IST2.scala 192:24]
  wire [31:0] FADD_5_io_out; // @[IST2.scala 192:24]
  wire  FADD_6_clock; // @[IST2.scala 201:24]
  wire  FADD_6_reset; // @[IST2.scala 201:24]
  wire [31:0] FADD_6_io_a; // @[IST2.scala 201:24]
  wire [31:0] FADD_6_io_b; // @[IST2.scala 201:24]
  wire [31:0] FADD_6_io_out; // @[IST2.scala 201:24]
  wire  FADD_7_clock; // @[IST2.scala 264:24]
  wire  FADD_7_reset; // @[IST2.scala 264:24]
  wire [31:0] FADD_7_io_a; // @[IST2.scala 264:24]
  wire [31:0] FADD_7_io_b; // @[IST2.scala 264:24]
  wire [31:0] FADD_7_io_out; // @[IST2.scala 264:24]
  wire  FADD_8_clock; // @[IST2.scala 273:24]
  wire  FADD_8_reset; // @[IST2.scala 273:24]
  wire [31:0] FADD_8_io_a; // @[IST2.scala 273:24]
  wire [31:0] FADD_8_io_b; // @[IST2.scala 273:24]
  wire [31:0] FADD_8_io_out; // @[IST2.scala 273:24]
  wire  FADD_MUL_15_clock; // @[IST2.scala 332:33]
  wire  FADD_MUL_15_reset; // @[IST2.scala 332:33]
  wire [31:0] FADD_MUL_15_io_a; // @[IST2.scala 332:33]
  wire [31:0] FADD_MUL_15_io_b; // @[IST2.scala 332:33]
  wire [31:0] FADD_MUL_15_io_c; // @[IST2.scala 332:33]
  wire [31:0] FADD_MUL_15_io_out; // @[IST2.scala 332:33]
  wire [31:0] FCMP_23_io_a; // @[IST2.scala 384:25]
  wire [31:0] FCMP_23_io_b; // @[IST2.scala 384:25]
  wire  FCMP_23_io_actual_out; // @[IST2.scala 384:25]
  reg [31:0] temp_0; // @[IST2.scala 44:33]
  reg [31:0] temp_1; // @[IST2.scala 45:33]
  reg [31:0] temp_2; // @[IST2.scala 46:33]
  reg [31:0] temp_3; // @[IST2.scala 47:33]
  reg [31:0] temp_4; // @[IST2.scala 48:33]
  reg [31:0] temp_5; // @[IST2.scala 49:33]
  reg [31:0] nodeid_ist2_temp_1_temp; // @[IST2.scala 51:42]
  reg [31:0] rayid_ist2_temp_1_temp; // @[IST2.scala 52:46]
  reg [31:0] t_temp_1_temp; // @[IST2.scala 53:56]
  reg [31:0] hitT_temp_1_temp; // @[IST2.scala 54:52]
  reg [127:0] v22_1_temp; // @[IST2.scala 55:60]
  reg [95:0] ray_o_in_1_temp; // @[IST2.scala 56:55]
  reg [95:0] ray_d_in_1_temp; // @[IST2.scala 57:55]
  reg  enable_1_temp; // @[IST2.scala 58:57]
  reg  break_1_temp; // @[IST2.scala 59:58]
  reg  ray_aabb_1_temp; // @[IST2.scala 60:51]
  reg  ray_aabb_2_temp; // @[IST2.scala 61:51]
  wire [127:0] _T = {io_v22_in_w,io_v22_in_z,io_v22_in_y,io_v22_in_x}; // @[Cat.scala 30:58]
  wire [95:0] _T_1 = {io_ray_o_in_z,io_ray_o_in_y,io_ray_o_in_x}; // @[Cat.scala 30:58]
  wire [95:0] _T_2 = {io_ray_d_in_z,io_ray_d_in_y,io_ray_d_in_x}; // @[Cat.scala 30:58]
  reg [31:0] nodeid_ist2_temp_1; // @[IST2.scala 129:37]
  reg [31:0] rayid_ist2_temp_1; // @[IST2.scala 130:41]
  reg [31:0] t_temp_1; // @[IST2.scala 131:51]
  reg [31:0] hitT_temp_1; // @[IST2.scala 132:47]
  reg [127:0] v22_1; // @[IST2.scala 133:55]
  reg [95:0] ray_o_in_1; // @[IST2.scala 134:50]
  reg [95:0] ray_d_in_1; // @[IST2.scala 135:50]
  reg  enable_1; // @[IST2.scala 136:52]
  reg  break_1; // @[IST2.scala 137:53]
  reg  ray_aabb_1; // @[IST2.scala 138:46]
  reg  ray_aabb_2; // @[IST2.scala 139:46]
  reg [31:0] nodeid_ist2_temp_2_temp; // @[IST2.scala 155:43]
  reg [31:0] rayid_ist2_temp_2_temp; // @[IST2.scala 156:46]
  reg [31:0] t_temp_2_temp; // @[IST2.scala 157:56]
  reg [31:0] hitT_temp_2_temp; // @[IST2.scala 158:52]
  reg [127:0] v22_2_temp; // @[IST2.scala 159:60]
  reg [95:0] ray_o_in_2_temp; // @[IST2.scala 160:55]
  reg [95:0] ray_d_in_2_temp; // @[IST2.scala 161:55]
  reg  enable_2_temp; // @[IST2.scala 162:55]
  reg  break_2_temp; // @[IST2.scala 163:58]
  reg  ray_aabb_1_2_temp; // @[IST2.scala 164:48]
  reg  ray_aabb_2_2_temp; // @[IST2.scala 165:48]
  reg [31:0] temp_6; // @[IST2.scala 179:50]
  reg [31:0] temp_7; // @[IST2.scala 180:50]
  reg [31:0] temp_0_2; // @[IST2.scala 181:47]
  reg [31:0] temp_0_3; // @[IST2.scala 182:47]
  reg [31:0] temp_5_2; // @[IST2.scala 184:46]
  reg [31:0] temp_5_3; // @[IST2.scala 185:46]
  reg [31:0] nodeid_ist2_temp_2; // @[IST2.scala 210:38]
  reg [31:0] rayid_ist2_temp_2; // @[IST2.scala 211:41]
  reg [31:0] t_temp_2; // @[IST2.scala 212:51]
  reg [31:0] hitT_temp_2; // @[IST2.scala 213:47]
  reg [127:0] v22_2; // @[IST2.scala 214:55]
  reg [95:0] ray_o_in_2; // @[IST2.scala 215:50]
  reg [95:0] ray_d_in_2; // @[IST2.scala 216:50]
  reg  enable_2; // @[IST2.scala 217:50]
  reg  break_2; // @[IST2.scala 218:53]
  reg  ray_aabb_1_2; // @[IST2.scala 219:43]
  reg  ray_aabb_2_2; // @[IST2.scala 220:43]
  reg [31:0] nodeid_ist2_temp_3_temp; // @[IST2.scala 236:43]
  reg [31:0] rayid_ist2_temp_3_temp; // @[IST2.scala 237:46]
  reg [31:0] t_temp_3_temp; // @[IST2.scala 238:56]
  reg [31:0] hitT_temp_3_temp; // @[IST2.scala 239:52]
  reg [127:0] v22_3_temp; // @[IST2.scala 240:60]
  reg [95:0] ray_o_in_3_temp; // @[IST2.scala 241:55]
  reg [95:0] ray_d_in_3_temp; // @[IST2.scala 242:55]
  reg  enable_3_temp; // @[IST2.scala 243:55]
  reg  break_3_temp; // @[IST2.scala 244:58]
  reg  ray_aabb_1_3_temp; // @[IST2.scala 245:48]
  reg  ray_aabb_2_3_temp; // @[IST2.scala 246:48]
  reg [31:0] Ox; // @[IST2.scala 261:58]
  reg [31:0] Dx; // @[IST2.scala 262:58]
  reg [31:0] nodeid_ist2_temp_3; // @[IST2.scala 282:38]
  reg [31:0] rayid_ist2_temp_3; // @[IST2.scala 283:41]
  reg [31:0] t_temp_3; // @[IST2.scala 284:51]
  reg [31:0] hitT_temp_3; // @[IST2.scala 285:47]
  reg [127:0] v22_3; // @[IST2.scala 286:55]
  reg [95:0] ray_o_in_3; // @[IST2.scala 287:50]
  reg [95:0] ray_d_in_3; // @[IST2.scala 288:50]
  reg  enable_3; // @[IST2.scala 289:50]
  reg  break_3; // @[IST2.scala 290:53]
  reg  ray_aabb_1_3; // @[IST2.scala 291:43]
  reg  ray_aabb_2_3; // @[IST2.scala 292:43]
  reg [31:0] nodeid_ist2_temp_4_temp; // @[IST2.scala 307:43]
  reg [31:0] rayid_ist2_temp_4_temp; // @[IST2.scala 308:46]
  reg [31:0] temp_u; // @[IST2.scala 309:53]
  reg [31:0] t_temp_4_temp; // @[IST2.scala 311:56]
  reg [31:0] hitT_temp_4_temp; // @[IST2.scala 312:52]
  reg [127:0] v22_4_temp; // @[IST2.scala 313:60]
  reg [95:0] ray_o_in_4_temp; // @[IST2.scala 314:55]
  reg [95:0] ray_d_in_4_temp; // @[IST2.scala 315:55]
  reg  enable_4_temp; // @[IST2.scala 316:55]
  reg  break_4_temp; // @[IST2.scala 317:58]
  reg  ray_aabb_1_4_temp; // @[IST2.scala 318:48]
  reg  ray_aabb_2_4_temp; // @[IST2.scala 319:48]
  reg [31:0] nodeid_ist2_temp_4; // @[IST2.scala 342:38]
  reg [31:0] rayid_ist2_temp_4; // @[IST2.scala 343:41]
  reg [31:0] t_temp_4; // @[IST2.scala 345:51]
  reg [31:0] hitT_temp_4; // @[IST2.scala 346:47]
  reg [127:0] v22_4; // @[IST2.scala 347:55]
  reg [95:0] ray_o_in_4; // @[IST2.scala 348:50]
  reg [95:0] ray_d_in_4; // @[IST2.scala 349:50]
  reg  enable_4; // @[IST2.scala 350:50]
  reg  break_4; // @[IST2.scala 351:53]
  reg  ray_aabb_1_4; // @[IST2.scala 352:43]
  reg  ray_aabb_2_4; // @[IST2.scala 353:43]
  wire  _T_15 = FCMP_23_io_actual_out > 1'h0 & enable_4; // @[IST2.scala 389:41]
  wire  _T_16 = ~break_4; // @[IST2.scala 389:69]
  wire  _T_20 = FCMP_23_io_actual_out < 1'h1 & enable_4; // @[IST2.scala 395:47]
  wire  _T_22 = FCMP_23_io_actual_out < 1'h1 & enable_4 & _T_16; // @[IST2.scala 395:65]
  wire  _T_27 = _T_15 & break_4; // @[IST2.scala 401:65]
  wire  _T_32 = _T_20 & break_4; // @[IST2.scala 407:65]
  wire  _GEN_6 = _T_15 & break_4 ? 1'h0 : _T_32; // @[IST2.scala 401:83 IST2.scala 406:34]
  wire  _GEN_9 = FCMP_23_io_actual_out < 1'h1 & enable_4 & _T_16 ? 1'h0 : _T_27; // @[IST2.scala 395:84 IST2.scala 399:32]
  wire  _GEN_10 = FCMP_23_io_actual_out < 1'h1 & enable_4 & _T_16 ? 1'h0 : _GEN_6; // @[IST2.scala 395:84 IST2.scala 400:34]
  MY_MULADD FADD_MUL_14 ( // @[IST2.scala 74:33]
    .clock(FADD_MUL_14_clock),
    .reset(FADD_MUL_14_reset),
    .io_a(FADD_MUL_14_io_a),
    .io_b(FADD_MUL_14_io_b),
    .io_c(FADD_MUL_14_io_c),
    .io_out(FADD_MUL_14_io_out)
  );
  MY_MUL FMUL_7 ( // @[IST2.scala 84:24]
    .clock(FMUL_7_clock),
    .reset(FMUL_7_reset),
    .io_a(FMUL_7_io_a),
    .io_b(FMUL_7_io_b),
    .io_out(FMUL_7_io_out)
  );
  MY_MUL FMUL_8 ( // @[IST2.scala 93:24]
    .clock(FMUL_8_clock),
    .reset(FMUL_8_reset),
    .io_a(FMUL_8_io_a),
    .io_b(FMUL_8_io_b),
    .io_out(FMUL_8_io_out)
  );
  MY_MUL FMUL_9 ( // @[IST2.scala 102:24]
    .clock(FMUL_9_clock),
    .reset(FMUL_9_reset),
    .io_a(FMUL_9_io_a),
    .io_b(FMUL_9_io_b),
    .io_out(FMUL_9_io_out)
  );
  MY_MUL FMUL_10 ( // @[IST2.scala 111:25]
    .clock(FMUL_10_clock),
    .reset(FMUL_10_reset),
    .io_a(FMUL_10_io_a),
    .io_b(FMUL_10_io_b),
    .io_out(FMUL_10_io_out)
  );
  MY_MUL FMUL_11 ( // @[IST2.scala 120:25]
    .clock(FMUL_11_clock),
    .reset(FMUL_11_reset),
    .io_a(FMUL_11_io_a),
    .io_b(FMUL_11_io_b),
    .io_out(FMUL_11_io_out)
  );
  MY_ADD FADD_5 ( // @[IST2.scala 192:24]
    .clock(FADD_5_clock),
    .reset(FADD_5_reset),
    .io_a(FADD_5_io_a),
    .io_b(FADD_5_io_b),
    .io_out(FADD_5_io_out)
  );
  MY_ADD FADD_6 ( // @[IST2.scala 201:24]
    .clock(FADD_6_clock),
    .reset(FADD_6_reset),
    .io_a(FADD_6_io_a),
    .io_b(FADD_6_io_b),
    .io_out(FADD_6_io_out)
  );
  MY_ADD FADD_7 ( // @[IST2.scala 264:24]
    .clock(FADD_7_clock),
    .reset(FADD_7_reset),
    .io_a(FADD_7_io_a),
    .io_b(FADD_7_io_b),
    .io_out(FADD_7_io_out)
  );
  MY_ADD FADD_8 ( // @[IST2.scala 273:24]
    .clock(FADD_8_clock),
    .reset(FADD_8_reset),
    .io_a(FADD_8_io_a),
    .io_b(FADD_8_io_b),
    .io_out(FADD_8_io_out)
  );
  MY_MULADD FADD_MUL_15 ( // @[IST2.scala 332:33]
    .clock(FADD_MUL_15_clock),
    .reset(FADD_MUL_15_reset),
    .io_a(FADD_MUL_15_io_a),
    .io_b(FADD_MUL_15_io_b),
    .io_c(FADD_MUL_15_io_c),
    .io_out(FADD_MUL_15_io_out)
  );
  ValExec_CompareRecF32_lt FCMP_23 ( // @[IST2.scala 384:25]
    .io_a(FCMP_23_io_a),
    .io_b(FCMP_23_io_b),
    .io_actual_out(FCMP_23_io_actual_out)
  );
  assign io_nodeid_ist2_out = nodeid_ist2_temp_4; // @[IST2.scala 367:37]
  assign io_rayid_ist2_out = rayid_ist2_temp_4; // @[IST2.scala 368:40]
  assign io_hiT_out = hitT_temp_4; // @[IST2.scala 370:47]
  assign io_u = temp_u; // @[IST2.scala 389:77 IST2.scala 390:45]
  assign io_pop_2 = FCMP_23_io_actual_out > 1'h0 & enable_4 & ~break_4 ? 1'h0 : _T_22; // @[IST2.scala 389:77 IST2.scala 392:38]
  assign io_t_out = t_temp_4; // @[IST2.scala 369:50]
  assign io_v22_out_x = v22_4[31:0]; // @[IST2.scala 371:53]
  assign io_v22_out_y = v22_4[63:32]; // @[IST2.scala 372:53]
  assign io_v22_out_z = v22_4[95:64]; // @[IST2.scala 373:53]
  assign io_v22_out_w = v22_4[127:96]; // @[IST2.scala 374:52]
  assign io_ray_o_out_x = ray_o_in_4[31:0]; // @[IST2.scala 375:54]
  assign io_ray_o_out_y = ray_o_in_4[63:32]; // @[IST2.scala 376:54]
  assign io_ray_o_out_z = ray_o_in_4[95:64]; // @[IST2.scala 377:54]
  assign io_ray_d_out_x = ray_d_in_4[31:0]; // @[IST2.scala 378:54]
  assign io_ray_d_out_y = ray_d_in_4[63:32]; // @[IST2.scala 379:54]
  assign io_ray_d_out_z = ray_d_in_4[95:64]; // @[IST2.scala 380:54]
  assign io_enable_IST3 = FCMP_23_io_actual_out > 1'h0 & enable_4 & ~break_4 | _GEN_9; // @[IST2.scala 389:77 IST2.scala 393:32]
  assign io_break_ist2 = break_4; // @[IST2.scala 381:43]
  assign io_break_out = FCMP_23_io_actual_out > 1'h0 & enable_4 & ~break_4 ? 1'h0 : _GEN_10; // @[IST2.scala 389:77 IST2.scala 394:34]
  assign io_RAY_AABB_1_out = ray_aabb_1_4; // @[IST2.scala 382:33]
  assign io_RAY_AABB_2_out = ray_aabb_2_4; // @[IST2.scala 383:33]
  assign FADD_MUL_14_clock = clock;
  assign FADD_MUL_14_reset = reset;
  assign FADD_MUL_14_io_a = io_ray_o_in_x; // @[IST2.scala 75:26]
  assign FADD_MUL_14_io_b = io_v11_in_x; // @[IST2.scala 76:26]
  assign FADD_MUL_14_io_c = io_v11_in_w; // @[IST2.scala 77:26]
  assign FMUL_7_clock = clock;
  assign FMUL_7_reset = reset;
  assign FMUL_7_io_a = io_ray_o_in_y; // @[IST2.scala 85:21]
  assign FMUL_7_io_b = io_v11_in_y; // @[IST2.scala 86:21]
  assign FMUL_8_clock = clock;
  assign FMUL_8_reset = reset;
  assign FMUL_8_io_a = io_ray_o_in_z; // @[IST2.scala 94:21]
  assign FMUL_8_io_b = io_v11_in_z; // @[IST2.scala 95:21]
  assign FMUL_9_clock = clock;
  assign FMUL_9_reset = reset;
  assign FMUL_9_io_a = io_ray_d_in_x; // @[IST2.scala 103:21]
  assign FMUL_9_io_b = io_v11_in_x; // @[IST2.scala 104:21]
  assign FMUL_10_clock = clock;
  assign FMUL_10_reset = reset;
  assign FMUL_10_io_a = io_ray_d_in_y; // @[IST2.scala 112:22]
  assign FMUL_10_io_b = io_v11_in_y; // @[IST2.scala 113:22]
  assign FMUL_11_clock = clock;
  assign FMUL_11_reset = reset;
  assign FMUL_11_io_a = io_ray_d_in_z; // @[IST2.scala 121:22]
  assign FMUL_11_io_b = io_v11_in_z; // @[IST2.scala 122:22]
  assign FADD_5_clock = clock;
  assign FADD_5_reset = reset;
  assign FADD_5_io_a = temp_1; // @[IST2.scala 193:21]
  assign FADD_5_io_b = temp_2; // @[IST2.scala 194:21]
  assign FADD_6_clock = clock;
  assign FADD_6_reset = reset;
  assign FADD_6_io_a = temp_3; // @[IST2.scala 202:21]
  assign FADD_6_io_b = temp_4; // @[IST2.scala 203:21]
  assign FADD_7_clock = clock;
  assign FADD_7_reset = reset;
  assign FADD_7_io_a = temp_0_3; // @[IST2.scala 265:21]
  assign FADD_7_io_b = temp_6; // @[IST2.scala 266:21]
  assign FADD_8_clock = clock;
  assign FADD_8_reset = reset;
  assign FADD_8_io_a = temp_5_3; // @[IST2.scala 274:21]
  assign FADD_8_io_b = temp_7; // @[IST2.scala 275:21]
  assign FADD_MUL_15_clock = clock;
  assign FADD_MUL_15_reset = reset;
  assign FADD_MUL_15_io_a = t_temp_3; // @[IST2.scala 333:26]
  assign FADD_MUL_15_io_b = Dx; // @[IST2.scala 334:26]
  assign FADD_MUL_15_io_c = Ox; // @[IST2.scala 335:26]
  assign FCMP_23_io_a = 32'h0; // @[IST2.scala 385:22]
  assign FCMP_23_io_b = temp_u; // @[IST2.scala 386:22]
  always @(posedge clock) begin
    if (reset) begin // @[IST2.scala 44:33]
      temp_0 <= 32'h0; // @[IST2.scala 44:33]
    end else begin
      temp_0 <= FADD_MUL_14_io_out; // @[IST2.scala 82:42]
    end
    if (reset) begin // @[IST2.scala 45:33]
      temp_1 <= 32'h0; // @[IST2.scala 45:33]
    end else begin
      temp_1 <= FMUL_7_io_out; // @[IST2.scala 91:42]
    end
    if (reset) begin // @[IST2.scala 46:33]
      temp_2 <= 32'h0; // @[IST2.scala 46:33]
    end else begin
      temp_2 <= FMUL_8_io_out; // @[IST2.scala 100:42]
    end
    if (reset) begin // @[IST2.scala 47:33]
      temp_3 <= 32'h0; // @[IST2.scala 47:33]
    end else begin
      temp_3 <= FMUL_9_io_out; // @[IST2.scala 109:42]
    end
    if (reset) begin // @[IST2.scala 48:33]
      temp_4 <= 32'h0; // @[IST2.scala 48:33]
    end else begin
      temp_4 <= FMUL_10_io_out; // @[IST2.scala 118:42]
    end
    if (reset) begin // @[IST2.scala 49:33]
      temp_5 <= 32'h0; // @[IST2.scala 49:33]
    end else begin
      temp_5 <= FMUL_11_io_out; // @[IST2.scala 127:42]
    end
    if (reset) begin // @[IST2.scala 51:42]
      nodeid_ist2_temp_1_temp <= 32'sh0; // @[IST2.scala 51:42]
    end else begin
      nodeid_ist2_temp_1_temp <= io_nodeid_leaf_2; // @[IST2.scala 63:34]
    end
    if (reset) begin // @[IST2.scala 52:46]
      rayid_ist2_temp_1_temp <= 32'h0; // @[IST2.scala 52:46]
    end else begin
      rayid_ist2_temp_1_temp <= io_rayid_leaf_2; // @[IST2.scala 64:37]
    end
    if (reset) begin // @[IST2.scala 53:56]
      t_temp_1_temp <= 32'h0; // @[IST2.scala 53:56]
    end else begin
      t_temp_1_temp <= io_t; // @[IST2.scala 65:47]
    end
    if (reset) begin // @[IST2.scala 54:52]
      hitT_temp_1_temp <= 32'h0; // @[IST2.scala 54:52]
    end else begin
      hitT_temp_1_temp <= io_hiT_in; // @[IST2.scala 66:43]
    end
    if (reset) begin // @[IST2.scala 55:60]
      v22_1_temp <= 128'h0; // @[IST2.scala 55:60]
    end else begin
      v22_1_temp <= _T; // @[IST2.scala 67:51]
    end
    if (reset) begin // @[IST2.scala 56:55]
      ray_o_in_1_temp <= 96'h0; // @[IST2.scala 56:55]
    end else begin
      ray_o_in_1_temp <= _T_1; // @[IST2.scala 68:45]
    end
    if (reset) begin // @[IST2.scala 57:55]
      ray_d_in_1_temp <= 96'h0; // @[IST2.scala 57:55]
    end else begin
      ray_d_in_1_temp <= _T_2; // @[IST2.scala 69:45]
    end
    if (reset) begin // @[IST2.scala 58:57]
      enable_1_temp <= 1'h0; // @[IST2.scala 58:57]
    end else begin
      enable_1_temp <= io_enable_IST2; // @[IST2.scala 70:48]
    end
    if (reset) begin // @[IST2.scala 59:58]
      break_1_temp <= 1'h0; // @[IST2.scala 59:58]
    end else begin
      break_1_temp <= io_break_in; // @[IST2.scala 71:50]
    end
    if (reset) begin // @[IST2.scala 60:51]
      ray_aabb_1_temp <= 1'h0; // @[IST2.scala 60:51]
    end else begin
      ray_aabb_1_temp <= io_RAY_AABB_1; // @[IST2.scala 72:45]
    end
    if (reset) begin // @[IST2.scala 61:51]
      ray_aabb_2_temp <= 1'h0; // @[IST2.scala 61:51]
    end else begin
      ray_aabb_2_temp <= io_RAY_AABB_2; // @[IST2.scala 73:45]
    end
    if (reset) begin // @[IST2.scala 129:37]
      nodeid_ist2_temp_1 <= 32'sh0; // @[IST2.scala 129:37]
    end else begin
      nodeid_ist2_temp_1 <= nodeid_ist2_temp_1_temp; // @[IST2.scala 141:29]
    end
    if (reset) begin // @[IST2.scala 130:41]
      rayid_ist2_temp_1 <= 32'h0; // @[IST2.scala 130:41]
    end else begin
      rayid_ist2_temp_1 <= rayid_ist2_temp_1_temp; // @[IST2.scala 142:32]
    end
    if (reset) begin // @[IST2.scala 131:51]
      t_temp_1 <= 32'h0; // @[IST2.scala 131:51]
    end else begin
      t_temp_1 <= t_temp_1_temp; // @[IST2.scala 143:42]
    end
    if (reset) begin // @[IST2.scala 132:47]
      hitT_temp_1 <= 32'h0; // @[IST2.scala 132:47]
    end else begin
      hitT_temp_1 <= hitT_temp_1_temp; // @[IST2.scala 144:38]
    end
    if (reset) begin // @[IST2.scala 133:55]
      v22_1 <= 128'h0; // @[IST2.scala 133:55]
    end else begin
      v22_1 <= v22_1_temp; // @[IST2.scala 145:46]
    end
    if (reset) begin // @[IST2.scala 134:50]
      ray_o_in_1 <= 96'h0; // @[IST2.scala 134:50]
    end else begin
      ray_o_in_1 <= ray_o_in_1_temp; // @[IST2.scala 146:40]
    end
    if (reset) begin // @[IST2.scala 135:50]
      ray_d_in_1 <= 96'h0; // @[IST2.scala 135:50]
    end else begin
      ray_d_in_1 <= ray_d_in_1_temp; // @[IST2.scala 147:40]
    end
    if (reset) begin // @[IST2.scala 136:52]
      enable_1 <= 1'h0; // @[IST2.scala 136:52]
    end else begin
      enable_1 <= enable_1_temp; // @[IST2.scala 148:43]
    end
    if (reset) begin // @[IST2.scala 137:53]
      break_1 <= 1'h0; // @[IST2.scala 137:53]
    end else begin
      break_1 <= break_1_temp; // @[IST2.scala 149:45]
    end
    if (reset) begin // @[IST2.scala 138:46]
      ray_aabb_1 <= 1'h0; // @[IST2.scala 138:46]
    end else begin
      ray_aabb_1 <= ray_aabb_1_temp; // @[IST2.scala 150:40]
    end
    if (reset) begin // @[IST2.scala 139:46]
      ray_aabb_2 <= 1'h0; // @[IST2.scala 139:46]
    end else begin
      ray_aabb_2 <= ray_aabb_2_temp; // @[IST2.scala 151:40]
    end
    if (reset) begin // @[IST2.scala 155:43]
      nodeid_ist2_temp_2_temp <= 32'sh0; // @[IST2.scala 155:43]
    end else begin
      nodeid_ist2_temp_2_temp <= nodeid_ist2_temp_1; // @[IST2.scala 167:34]
    end
    if (reset) begin // @[IST2.scala 156:46]
      rayid_ist2_temp_2_temp <= 32'h0; // @[IST2.scala 156:46]
    end else begin
      rayid_ist2_temp_2_temp <= rayid_ist2_temp_1; // @[IST2.scala 168:37]
    end
    if (reset) begin // @[IST2.scala 157:56]
      t_temp_2_temp <= 32'h0; // @[IST2.scala 157:56]
    end else begin
      t_temp_2_temp <= t_temp_1; // @[IST2.scala 169:47]
    end
    if (reset) begin // @[IST2.scala 158:52]
      hitT_temp_2_temp <= 32'h0; // @[IST2.scala 158:52]
    end else begin
      hitT_temp_2_temp <= hitT_temp_1; // @[IST2.scala 170:43]
    end
    if (reset) begin // @[IST2.scala 159:60]
      v22_2_temp <= 128'h0; // @[IST2.scala 159:60]
    end else begin
      v22_2_temp <= v22_1; // @[IST2.scala 171:51]
    end
    if (reset) begin // @[IST2.scala 160:55]
      ray_o_in_2_temp <= 96'h0; // @[IST2.scala 160:55]
    end else begin
      ray_o_in_2_temp <= ray_o_in_1; // @[IST2.scala 172:45]
    end
    if (reset) begin // @[IST2.scala 161:55]
      ray_d_in_2_temp <= 96'h0; // @[IST2.scala 161:55]
    end else begin
      ray_d_in_2_temp <= ray_d_in_1; // @[IST2.scala 173:45]
    end
    if (reset) begin // @[IST2.scala 162:55]
      enable_2_temp <= 1'h0; // @[IST2.scala 162:55]
    end else begin
      enable_2_temp <= enable_1; // @[IST2.scala 174:47]
    end
    if (reset) begin // @[IST2.scala 163:58]
      break_2_temp <= 1'h0; // @[IST2.scala 163:58]
    end else begin
      break_2_temp <= break_1; // @[IST2.scala 175:50]
    end
    if (reset) begin // @[IST2.scala 164:48]
      ray_aabb_1_2_temp <= 1'h0; // @[IST2.scala 164:48]
    end else begin
      ray_aabb_1_2_temp <= ray_aabb_1; // @[IST2.scala 176:41]
    end
    if (reset) begin // @[IST2.scala 165:48]
      ray_aabb_2_2_temp <= 1'h0; // @[IST2.scala 165:48]
    end else begin
      ray_aabb_2_2_temp <= ray_aabb_2; // @[IST2.scala 177:41]
    end
    if (reset) begin // @[IST2.scala 179:50]
      temp_6 <= 32'h0; // @[IST2.scala 179:50]
    end else begin
      temp_6 <= FADD_5_io_out; // @[IST2.scala 199:26]
    end
    if (reset) begin // @[IST2.scala 180:50]
      temp_7 <= 32'h0; // @[IST2.scala 180:50]
    end else begin
      temp_7 <= FADD_6_io_out; // @[IST2.scala 208:26]
    end
    if (reset) begin // @[IST2.scala 181:47]
      temp_0_2 <= 32'h0; // @[IST2.scala 181:47]
    end else begin
      temp_0_2 <= temp_0; // @[IST2.scala 186:41]
    end
    if (reset) begin // @[IST2.scala 182:47]
      temp_0_3 <= 32'h0; // @[IST2.scala 182:47]
    end else begin
      temp_0_3 <= temp_0_2; // @[IST2.scala 187:41]
    end
    if (reset) begin // @[IST2.scala 184:46]
      temp_5_2 <= 32'h0; // @[IST2.scala 184:46]
    end else begin
      temp_5_2 <= temp_5; // @[IST2.scala 188:41]
    end
    if (reset) begin // @[IST2.scala 185:46]
      temp_5_3 <= 32'h0; // @[IST2.scala 185:46]
    end else begin
      temp_5_3 <= temp_5_2; // @[IST2.scala 189:41]
    end
    if (reset) begin // @[IST2.scala 210:38]
      nodeid_ist2_temp_2 <= 32'sh0; // @[IST2.scala 210:38]
    end else begin
      nodeid_ist2_temp_2 <= nodeid_ist2_temp_2_temp; // @[IST2.scala 222:29]
    end
    if (reset) begin // @[IST2.scala 211:41]
      rayid_ist2_temp_2 <= 32'h0; // @[IST2.scala 211:41]
    end else begin
      rayid_ist2_temp_2 <= rayid_ist2_temp_2_temp; // @[IST2.scala 223:32]
    end
    if (reset) begin // @[IST2.scala 212:51]
      t_temp_2 <= 32'h0; // @[IST2.scala 212:51]
    end else begin
      t_temp_2 <= t_temp_2_temp; // @[IST2.scala 224:42]
    end
    if (reset) begin // @[IST2.scala 213:47]
      hitT_temp_2 <= 32'h0; // @[IST2.scala 213:47]
    end else begin
      hitT_temp_2 <= hitT_temp_2_temp; // @[IST2.scala 225:38]
    end
    if (reset) begin // @[IST2.scala 214:55]
      v22_2 <= 128'h0; // @[IST2.scala 214:55]
    end else begin
      v22_2 <= v22_2_temp; // @[IST2.scala 226:46]
    end
    if (reset) begin // @[IST2.scala 215:50]
      ray_o_in_2 <= 96'h0; // @[IST2.scala 215:50]
    end else begin
      ray_o_in_2 <= ray_o_in_2_temp; // @[IST2.scala 227:40]
    end
    if (reset) begin // @[IST2.scala 216:50]
      ray_d_in_2 <= 96'h0; // @[IST2.scala 216:50]
    end else begin
      ray_d_in_2 <= ray_d_in_2_temp; // @[IST2.scala 228:40]
    end
    if (reset) begin // @[IST2.scala 217:50]
      enable_2 <= 1'h0; // @[IST2.scala 217:50]
    end else begin
      enable_2 <= enable_2_temp; // @[IST2.scala 229:42]
    end
    if (reset) begin // @[IST2.scala 218:53]
      break_2 <= 1'h0; // @[IST2.scala 218:53]
    end else begin
      break_2 <= break_2_temp; // @[IST2.scala 230:45]
    end
    if (reset) begin // @[IST2.scala 219:43]
      ray_aabb_1_2 <= 1'h0; // @[IST2.scala 219:43]
    end else begin
      ray_aabb_1_2 <= ray_aabb_1_2_temp; // @[IST2.scala 231:37]
    end
    if (reset) begin // @[IST2.scala 220:43]
      ray_aabb_2_2 <= 1'h0; // @[IST2.scala 220:43]
    end else begin
      ray_aabb_2_2 <= ray_aabb_2_2_temp; // @[IST2.scala 232:37]
    end
    if (reset) begin // @[IST2.scala 236:43]
      nodeid_ist2_temp_3_temp <= 32'sh0; // @[IST2.scala 236:43]
    end else begin
      nodeid_ist2_temp_3_temp <= nodeid_ist2_temp_2; // @[IST2.scala 248:37]
    end
    if (reset) begin // @[IST2.scala 237:46]
      rayid_ist2_temp_3_temp <= 32'h0; // @[IST2.scala 237:46]
    end else begin
      rayid_ist2_temp_3_temp <= rayid_ist2_temp_2; // @[IST2.scala 249:40]
    end
    if (reset) begin // @[IST2.scala 238:56]
      t_temp_3_temp <= 32'h0; // @[IST2.scala 238:56]
    end else begin
      t_temp_3_temp <= t_temp_2; // @[IST2.scala 250:50]
    end
    if (reset) begin // @[IST2.scala 239:52]
      hitT_temp_3_temp <= 32'h0; // @[IST2.scala 239:52]
    end else begin
      hitT_temp_3_temp <= hitT_temp_2; // @[IST2.scala 251:46]
    end
    if (reset) begin // @[IST2.scala 240:60]
      v22_3_temp <= 128'h0; // @[IST2.scala 240:60]
    end else begin
      v22_3_temp <= v22_2; // @[IST2.scala 252:54]
    end
    if (reset) begin // @[IST2.scala 241:55]
      ray_o_in_3_temp <= 96'h0; // @[IST2.scala 241:55]
    end else begin
      ray_o_in_3_temp <= ray_o_in_2; // @[IST2.scala 253:45]
    end
    if (reset) begin // @[IST2.scala 242:55]
      ray_d_in_3_temp <= 96'h0; // @[IST2.scala 242:55]
    end else begin
      ray_d_in_3_temp <= ray_d_in_2; // @[IST2.scala 254:45]
    end
    if (reset) begin // @[IST2.scala 243:55]
      enable_3_temp <= 1'h0; // @[IST2.scala 243:55]
    end else begin
      enable_3_temp <= enable_2; // @[IST2.scala 255:47]
    end
    if (reset) begin // @[IST2.scala 244:58]
      break_3_temp <= 1'h0; // @[IST2.scala 244:58]
    end else begin
      break_3_temp <= break_2; // @[IST2.scala 256:49]
    end
    if (reset) begin // @[IST2.scala 245:48]
      ray_aabb_1_3_temp <= 1'h0; // @[IST2.scala 245:48]
    end else begin
      ray_aabb_1_3_temp <= ray_aabb_1_2; // @[IST2.scala 257:41]
    end
    if (reset) begin // @[IST2.scala 246:48]
      ray_aabb_2_3_temp <= 1'h0; // @[IST2.scala 246:48]
    end else begin
      ray_aabb_2_3_temp <= ray_aabb_2_2; // @[IST2.scala 258:41]
    end
    if (reset) begin // @[IST2.scala 261:58]
      Ox <= 32'h0; // @[IST2.scala 261:58]
    end else begin
      Ox <= FADD_7_io_out; // @[IST2.scala 271:26]
    end
    if (reset) begin // @[IST2.scala 262:58]
      Dx <= 32'h0; // @[IST2.scala 262:58]
    end else begin
      Dx <= FADD_8_io_out; // @[IST2.scala 280:26]
    end
    if (reset) begin // @[IST2.scala 282:38]
      nodeid_ist2_temp_3 <= 32'sh0; // @[IST2.scala 282:38]
    end else begin
      nodeid_ist2_temp_3 <= nodeid_ist2_temp_3_temp; // @[IST2.scala 294:32]
    end
    if (reset) begin // @[IST2.scala 283:41]
      rayid_ist2_temp_3 <= 32'h0; // @[IST2.scala 283:41]
    end else begin
      rayid_ist2_temp_3 <= rayid_ist2_temp_3_temp; // @[IST2.scala 295:35]
    end
    if (reset) begin // @[IST2.scala 284:51]
      t_temp_3 <= 32'h0; // @[IST2.scala 284:51]
    end else begin
      t_temp_3 <= t_temp_3_temp; // @[IST2.scala 296:45]
    end
    if (reset) begin // @[IST2.scala 285:47]
      hitT_temp_3 <= 32'h0; // @[IST2.scala 285:47]
    end else begin
      hitT_temp_3 <= hitT_temp_3_temp; // @[IST2.scala 297:41]
    end
    if (reset) begin // @[IST2.scala 286:55]
      v22_3 <= 128'h0; // @[IST2.scala 286:55]
    end else begin
      v22_3 <= v22_3_temp; // @[IST2.scala 298:49]
    end
    if (reset) begin // @[IST2.scala 287:50]
      ray_o_in_3 <= 96'h0; // @[IST2.scala 287:50]
    end else begin
      ray_o_in_3 <= ray_o_in_3_temp; // @[IST2.scala 299:40]
    end
    if (reset) begin // @[IST2.scala 288:50]
      ray_d_in_3 <= 96'h0; // @[IST2.scala 288:50]
    end else begin
      ray_d_in_3 <= ray_d_in_3_temp; // @[IST2.scala 300:40]
    end
    if (reset) begin // @[IST2.scala 289:50]
      enable_3 <= 1'h0; // @[IST2.scala 289:50]
    end else begin
      enable_3 <= enable_3_temp; // @[IST2.scala 301:42]
    end
    if (reset) begin // @[IST2.scala 290:53]
      break_3 <= 1'h0; // @[IST2.scala 290:53]
    end else begin
      break_3 <= break_3_temp; // @[IST2.scala 302:44]
    end
    if (reset) begin // @[IST2.scala 291:43]
      ray_aabb_1_3 <= 1'h0; // @[IST2.scala 291:43]
    end else begin
      ray_aabb_1_3 <= ray_aabb_1_3_temp; // @[IST2.scala 303:37]
    end
    if (reset) begin // @[IST2.scala 292:43]
      ray_aabb_2_3 <= 1'h0; // @[IST2.scala 292:43]
    end else begin
      ray_aabb_2_3 <= ray_aabb_2_3_temp; // @[IST2.scala 304:37]
    end
    if (reset) begin // @[IST2.scala 307:43]
      nodeid_ist2_temp_4_temp <= 32'sh0; // @[IST2.scala 307:43]
    end else begin
      nodeid_ist2_temp_4_temp <= nodeid_ist2_temp_3; // @[IST2.scala 321:37]
    end
    if (reset) begin // @[IST2.scala 308:46]
      rayid_ist2_temp_4_temp <= 32'h0; // @[IST2.scala 308:46]
    end else begin
      rayid_ist2_temp_4_temp <= rayid_ist2_temp_3; // @[IST2.scala 322:40]
    end
    if (reset) begin // @[IST2.scala 309:53]
      temp_u <= 32'h0; // @[IST2.scala 309:53]
    end else begin
      temp_u <= FADD_MUL_15_io_out; // @[IST2.scala 340:42]
    end
    if (reset) begin // @[IST2.scala 311:56]
      t_temp_4_temp <= 32'h0; // @[IST2.scala 311:56]
    end else begin
      t_temp_4_temp <= t_temp_3; // @[IST2.scala 323:50]
    end
    if (reset) begin // @[IST2.scala 312:52]
      hitT_temp_4_temp <= 32'h0; // @[IST2.scala 312:52]
    end else begin
      hitT_temp_4_temp <= hitT_temp_3; // @[IST2.scala 324:46]
    end
    if (reset) begin // @[IST2.scala 313:60]
      v22_4_temp <= 128'h0; // @[IST2.scala 313:60]
    end else begin
      v22_4_temp <= v22_3; // @[IST2.scala 325:54]
    end
    if (reset) begin // @[IST2.scala 314:55]
      ray_o_in_4_temp <= 96'h0; // @[IST2.scala 314:55]
    end else begin
      ray_o_in_4_temp <= ray_o_in_3; // @[IST2.scala 327:45]
    end
    if (reset) begin // @[IST2.scala 315:55]
      ray_d_in_4_temp <= 96'h0; // @[IST2.scala 315:55]
    end else begin
      ray_d_in_4_temp <= ray_d_in_3; // @[IST2.scala 326:45]
    end
    if (reset) begin // @[IST2.scala 316:55]
      enable_4_temp <= 1'h0; // @[IST2.scala 316:55]
    end else begin
      enable_4_temp <= enable_3; // @[IST2.scala 328:47]
    end
    if (reset) begin // @[IST2.scala 317:58]
      break_4_temp <= 1'h0; // @[IST2.scala 317:58]
    end else begin
      break_4_temp <= break_3; // @[IST2.scala 329:48]
    end
    if (reset) begin // @[IST2.scala 318:48]
      ray_aabb_1_4_temp <= 1'h0; // @[IST2.scala 318:48]
    end else begin
      ray_aabb_1_4_temp <= ray_aabb_1_3; // @[IST2.scala 330:42]
    end
    if (reset) begin // @[IST2.scala 319:48]
      ray_aabb_2_4_temp <= 1'h0; // @[IST2.scala 319:48]
    end else begin
      ray_aabb_2_4_temp <= ray_aabb_2_3; // @[IST2.scala 331:42]
    end
    if (reset) begin // @[IST2.scala 342:38]
      nodeid_ist2_temp_4 <= 32'sh0; // @[IST2.scala 342:38]
    end else begin
      nodeid_ist2_temp_4 <= nodeid_ist2_temp_4_temp; // @[IST2.scala 355:32]
    end
    if (reset) begin // @[IST2.scala 343:41]
      rayid_ist2_temp_4 <= 32'h0; // @[IST2.scala 343:41]
    end else begin
      rayid_ist2_temp_4 <= rayid_ist2_temp_4_temp; // @[IST2.scala 356:35]
    end
    if (reset) begin // @[IST2.scala 345:51]
      t_temp_4 <= 32'h0; // @[IST2.scala 345:51]
    end else begin
      t_temp_4 <= t_temp_4_temp; // @[IST2.scala 357:45]
    end
    if (reset) begin // @[IST2.scala 346:47]
      hitT_temp_4 <= 32'h0; // @[IST2.scala 346:47]
    end else begin
      hitT_temp_4 <= hitT_temp_4_temp; // @[IST2.scala 358:41]
    end
    if (reset) begin // @[IST2.scala 347:55]
      v22_4 <= 128'h0; // @[IST2.scala 347:55]
    end else begin
      v22_4 <= v22_4_temp; // @[IST2.scala 359:49]
    end
    if (reset) begin // @[IST2.scala 348:50]
      ray_o_in_4 <= 96'h0; // @[IST2.scala 348:50]
    end else begin
      ray_o_in_4 <= ray_o_in_4_temp; // @[IST2.scala 361:40]
    end
    if (reset) begin // @[IST2.scala 349:50]
      ray_d_in_4 <= 96'h0; // @[IST2.scala 349:50]
    end else begin
      ray_d_in_4 <= ray_d_in_4_temp; // @[IST2.scala 360:40]
    end
    if (reset) begin // @[IST2.scala 350:50]
      enable_4 <= 1'h0; // @[IST2.scala 350:50]
    end else begin
      enable_4 <= enable_4_temp; // @[IST2.scala 362:42]
    end
    if (reset) begin // @[IST2.scala 351:53]
      break_4 <= 1'h0; // @[IST2.scala 351:53]
    end else begin
      break_4 <= break_4_temp; // @[IST2.scala 363:43]
    end
    if (reset) begin // @[IST2.scala 352:43]
      ray_aabb_1_4 <= 1'h0; // @[IST2.scala 352:43]
    end else begin
      ray_aabb_1_4 <= ray_aabb_1_4_temp; // @[IST2.scala 364:37]
    end
    if (reset) begin // @[IST2.scala 353:43]
      ray_aabb_2_4 <= 1'h0; // @[IST2.scala 353:43]
    end else begin
      ray_aabb_2_4 <= ray_aabb_2_4_temp; // @[IST2.scala 365:37]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  temp_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  temp_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  temp_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  temp_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  temp_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  temp_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  nodeid_ist2_temp_1_temp = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  rayid_ist2_temp_1_temp = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  t_temp_1_temp = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  hitT_temp_1_temp = _RAND_9[31:0];
  _RAND_10 = {4{`RANDOM}};
  v22_1_temp = _RAND_10[127:0];
  _RAND_11 = {3{`RANDOM}};
  ray_o_in_1_temp = _RAND_11[95:0];
  _RAND_12 = {3{`RANDOM}};
  ray_d_in_1_temp = _RAND_12[95:0];
  _RAND_13 = {1{`RANDOM}};
  enable_1_temp = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  break_1_temp = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  ray_aabb_1_temp = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  ray_aabb_2_temp = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  nodeid_ist2_temp_1 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  rayid_ist2_temp_1 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  t_temp_1 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  hitT_temp_1 = _RAND_20[31:0];
  _RAND_21 = {4{`RANDOM}};
  v22_1 = _RAND_21[127:0];
  _RAND_22 = {3{`RANDOM}};
  ray_o_in_1 = _RAND_22[95:0];
  _RAND_23 = {3{`RANDOM}};
  ray_d_in_1 = _RAND_23[95:0];
  _RAND_24 = {1{`RANDOM}};
  enable_1 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  break_1 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  ray_aabb_1 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  ray_aabb_2 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  nodeid_ist2_temp_2_temp = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  rayid_ist2_temp_2_temp = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  t_temp_2_temp = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  hitT_temp_2_temp = _RAND_31[31:0];
  _RAND_32 = {4{`RANDOM}};
  v22_2_temp = _RAND_32[127:0];
  _RAND_33 = {3{`RANDOM}};
  ray_o_in_2_temp = _RAND_33[95:0];
  _RAND_34 = {3{`RANDOM}};
  ray_d_in_2_temp = _RAND_34[95:0];
  _RAND_35 = {1{`RANDOM}};
  enable_2_temp = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  break_2_temp = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  ray_aabb_1_2_temp = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  ray_aabb_2_2_temp = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  temp_6 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  temp_7 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  temp_0_2 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  temp_0_3 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  temp_5_2 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  temp_5_3 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  nodeid_ist2_temp_2 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  rayid_ist2_temp_2 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  t_temp_2 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  hitT_temp_2 = _RAND_48[31:0];
  _RAND_49 = {4{`RANDOM}};
  v22_2 = _RAND_49[127:0];
  _RAND_50 = {3{`RANDOM}};
  ray_o_in_2 = _RAND_50[95:0];
  _RAND_51 = {3{`RANDOM}};
  ray_d_in_2 = _RAND_51[95:0];
  _RAND_52 = {1{`RANDOM}};
  enable_2 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  break_2 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  ray_aabb_1_2 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  ray_aabb_2_2 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  nodeid_ist2_temp_3_temp = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  rayid_ist2_temp_3_temp = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  t_temp_3_temp = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  hitT_temp_3_temp = _RAND_59[31:0];
  _RAND_60 = {4{`RANDOM}};
  v22_3_temp = _RAND_60[127:0];
  _RAND_61 = {3{`RANDOM}};
  ray_o_in_3_temp = _RAND_61[95:0];
  _RAND_62 = {3{`RANDOM}};
  ray_d_in_3_temp = _RAND_62[95:0];
  _RAND_63 = {1{`RANDOM}};
  enable_3_temp = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  break_3_temp = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  ray_aabb_1_3_temp = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  ray_aabb_2_3_temp = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  Ox = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  Dx = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  nodeid_ist2_temp_3 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  rayid_ist2_temp_3 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  t_temp_3 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  hitT_temp_3 = _RAND_72[31:0];
  _RAND_73 = {4{`RANDOM}};
  v22_3 = _RAND_73[127:0];
  _RAND_74 = {3{`RANDOM}};
  ray_o_in_3 = _RAND_74[95:0];
  _RAND_75 = {3{`RANDOM}};
  ray_d_in_3 = _RAND_75[95:0];
  _RAND_76 = {1{`RANDOM}};
  enable_3 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  break_3 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  ray_aabb_1_3 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  ray_aabb_2_3 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  nodeid_ist2_temp_4_temp = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  rayid_ist2_temp_4_temp = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  temp_u = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  t_temp_4_temp = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  hitT_temp_4_temp = _RAND_84[31:0];
  _RAND_85 = {4{`RANDOM}};
  v22_4_temp = _RAND_85[127:0];
  _RAND_86 = {3{`RANDOM}};
  ray_o_in_4_temp = _RAND_86[95:0];
  _RAND_87 = {3{`RANDOM}};
  ray_d_in_4_temp = _RAND_87[95:0];
  _RAND_88 = {1{`RANDOM}};
  enable_4_temp = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  break_4_temp = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  ray_aabb_1_4_temp = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  ray_aabb_2_4_temp = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  nodeid_ist2_temp_4 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  rayid_ist2_temp_4 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  t_temp_4 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  hitT_temp_4 = _RAND_95[31:0];
  _RAND_96 = {4{`RANDOM}};
  v22_4 = _RAND_96[127:0];
  _RAND_97 = {3{`RANDOM}};
  ray_o_in_4 = _RAND_97[95:0];
  _RAND_98 = {3{`RANDOM}};
  ray_d_in_4 = _RAND_98[95:0];
  _RAND_99 = {1{`RANDOM}};
  enable_4 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  break_4 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  ray_aabb_1_4 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  ray_aabb_2_4 = _RAND_102[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IST3(
  input         clock,
  input         reset,
  input         io_enable_IST3,
  input  [31:0] io_nodeid_leaf_3,
  input  [31:0] io_rayid_leaf_3,
  input  [31:0] io_hiT_in,
  input  [31:0] io_t_in,
  input  [31:0] io_v22_in_x,
  input  [31:0] io_v22_in_y,
  input  [31:0] io_v22_in_z,
  input  [31:0] io_v22_in_w,
  input  [31:0] io_ray_o_in_x,
  input  [31:0] io_ray_o_in_y,
  input  [31:0] io_ray_o_in_z,
  input  [31:0] io_ray_d_in_x,
  input  [31:0] io_ray_d_in_y,
  input  [31:0] io_ray_d_in_z,
  input  [31:0] io_u_in,
  input         io_break_in,
  input         io_RAY_AABB_1,
  input         io_RAY_AABB_2,
  output [31:0] io_nodeid_ist3_out,
  output [31:0] io_rayid_ist3_out,
  output [31:0] io_hiT_out,
  output        io_hitT_en,
  output        io_pop_3,
  output [31:0] io_hitIndex,
  output        io_break_out,
  output        io_RAY_AABB_1_out,
  output        io_RAY_AABB_2_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
`endif // RANDOMIZE_REG_INIT
  wire  FADD_MUL_16_clock; // @[IST3.scala 70:33]
  wire  FADD_MUL_16_reset; // @[IST3.scala 70:33]
  wire [31:0] FADD_MUL_16_io_a; // @[IST3.scala 70:33]
  wire [31:0] FADD_MUL_16_io_b; // @[IST3.scala 70:33]
  wire [31:0] FADD_MUL_16_io_c; // @[IST3.scala 70:33]
  wire [31:0] FADD_MUL_16_io_out; // @[IST3.scala 70:33]
  wire  FMUL_12_clock; // @[IST3.scala 80:25]
  wire  FMUL_12_reset; // @[IST3.scala 80:25]
  wire [31:0] FMUL_12_io_a; // @[IST3.scala 80:25]
  wire [31:0] FMUL_12_io_b; // @[IST3.scala 80:25]
  wire [31:0] FMUL_12_io_out; // @[IST3.scala 80:25]
  wire  FMUL_13_clock; // @[IST3.scala 89:25]
  wire  FMUL_13_reset; // @[IST3.scala 89:25]
  wire [31:0] FMUL_13_io_a; // @[IST3.scala 89:25]
  wire [31:0] FMUL_13_io_b; // @[IST3.scala 89:25]
  wire [31:0] FMUL_13_io_out; // @[IST3.scala 89:25]
  wire  FMUL_14_clock; // @[IST3.scala 98:25]
  wire  FMUL_14_reset; // @[IST3.scala 98:25]
  wire [31:0] FMUL_14_io_a; // @[IST3.scala 98:25]
  wire [31:0] FMUL_14_io_b; // @[IST3.scala 98:25]
  wire [31:0] FMUL_14_io_out; // @[IST3.scala 98:25]
  wire  FMUL_15_clock; // @[IST3.scala 107:25]
  wire  FMUL_15_reset; // @[IST3.scala 107:25]
  wire [31:0] FMUL_15_io_a; // @[IST3.scala 107:25]
  wire [31:0] FMUL_15_io_b; // @[IST3.scala 107:25]
  wire [31:0] FMUL_15_io_out; // @[IST3.scala 107:25]
  wire  FMUL_16_clock; // @[IST3.scala 116:25]
  wire  FMUL_16_reset; // @[IST3.scala 116:25]
  wire [31:0] FMUL_16_io_a; // @[IST3.scala 116:25]
  wire [31:0] FMUL_16_io_b; // @[IST3.scala 116:25]
  wire [31:0] FMUL_16_io_out; // @[IST3.scala 116:25]
  wire  FADD_9_clock; // @[IST3.scala 178:24]
  wire  FADD_9_reset; // @[IST3.scala 178:24]
  wire [31:0] FADD_9_io_a; // @[IST3.scala 178:24]
  wire [31:0] FADD_9_io_b; // @[IST3.scala 178:24]
  wire [31:0] FADD_9_io_out; // @[IST3.scala 178:24]
  wire  FADD_10_clock; // @[IST3.scala 187:25]
  wire  FADD_10_reset; // @[IST3.scala 187:25]
  wire [31:0] FADD_10_io_a; // @[IST3.scala 187:25]
  wire [31:0] FADD_10_io_b; // @[IST3.scala 187:25]
  wire [31:0] FADD_10_io_out; // @[IST3.scala 187:25]
  wire  FADD_11_clock; // @[IST3.scala 238:25]
  wire  FADD_11_reset; // @[IST3.scala 238:25]
  wire [31:0] FADD_11_io_a; // @[IST3.scala 238:25]
  wire [31:0] FADD_11_io_b; // @[IST3.scala 238:25]
  wire [31:0] FADD_11_io_out; // @[IST3.scala 238:25]
  wire  FADD_12_clock; // @[IST3.scala 247:25]
  wire  FADD_12_reset; // @[IST3.scala 247:25]
  wire [31:0] FADD_12_io_a; // @[IST3.scala 247:25]
  wire [31:0] FADD_12_io_b; // @[IST3.scala 247:25]
  wire [31:0] FADD_12_io_out; // @[IST3.scala 247:25]
  wire  FADD_MUL_17_clock; // @[IST3.scala 299:33]
  wire  FADD_MUL_17_reset; // @[IST3.scala 299:33]
  wire [31:0] FADD_MUL_17_io_a; // @[IST3.scala 299:33]
  wire [31:0] FADD_MUL_17_io_b; // @[IST3.scala 299:33]
  wire [31:0] FADD_MUL_17_io_c; // @[IST3.scala 299:33]
  wire [31:0] FADD_MUL_17_io_out; // @[IST3.scala 299:33]
  wire [31:0] FCMP_24_io_a; // @[IST3.scala 350:25]
  wire [31:0] FCMP_24_io_b; // @[IST3.scala 350:25]
  wire  FCMP_24_io_actual_out; // @[IST3.scala 350:25]
  wire  FADD_13_clock; // @[IST3.scala 364:25]
  wire  FADD_13_reset; // @[IST3.scala 364:25]
  wire [31:0] FADD_13_io_a; // @[IST3.scala 364:25]
  wire [31:0] FADD_13_io_b; // @[IST3.scala 364:25]
  wire [31:0] FADD_13_io_out; // @[IST3.scala 364:25]
  wire [31:0] FCMP_25_io_a; // @[IST3.scala 398:25]
  wire [31:0] FCMP_25_io_b; // @[IST3.scala 398:25]
  wire  FCMP_25_io_actual_out; // @[IST3.scala 398:25]
  reg [31:0] temp_0; // @[IST3.scala 44:33]
  reg [31:0] temp_1; // @[IST3.scala 45:33]
  reg [31:0] temp_2; // @[IST3.scala 46:33]
  reg [31:0] temp_3; // @[IST3.scala 47:33]
  reg [31:0] temp_4; // @[IST3.scala 48:33]
  reg [31:0] temp_5; // @[IST3.scala 49:33]
  reg [31:0] nodeid_ist3_temp_1_temp; // @[IST3.scala 51:42]
  reg [31:0] rayid_ist3_temp_1_temp; // @[IST3.scala 52:46]
  reg [31:0] t_temp_1_temp; // @[IST3.scala 53:56]
  reg [31:0] u_temp_1_temp; // @[IST3.scala 54:54]
  reg [31:0] hitT_temp_1_temp; // @[IST3.scala 55:52]
  reg  enable_1_temp; // @[IST3.scala 56:55]
  reg  break_1_temp; // @[IST3.scala 57:56]
  reg  ray_aabb_1_temp; // @[IST3.scala 58:51]
  reg  ray_aabb_2_temp; // @[IST3.scala 59:51]
  reg [31:0] nodeid_ist3_temp_1; // @[IST3.scala 126:37]
  reg [31:0] rayid_ist3_temp_1; // @[IST3.scala 127:41]
  reg [31:0] t_temp_1; // @[IST3.scala 128:51]
  reg [31:0] u_temp_1; // @[IST3.scala 129:49]
  reg [31:0] hitT_temp_1; // @[IST3.scala 130:47]
  reg  enable_1; // @[IST3.scala 131:50]
  reg  break_1; // @[IST3.scala 132:51]
  reg  ray_aabb_1; // @[IST3.scala 133:46]
  reg  ray_aabb_2; // @[IST3.scala 134:46]
  reg [31:0] nodeid_ist3_temp_2_temp; // @[IST3.scala 145:43]
  reg [31:0] rayid_ist3_temp_2_temp; // @[IST3.scala 146:46]
  reg [31:0] t_temp_2_temp; // @[IST3.scala 147:56]
  reg [31:0] u_temp_2_temp; // @[IST3.scala 148:55]
  reg [31:0] hitT_temp_2_temp; // @[IST3.scala 149:52]
  reg  enable_2_temp; // @[IST3.scala 150:55]
  reg  break_2_temp; // @[IST3.scala 151:56]
  reg  ray_aabb_1_2_temp; // @[IST3.scala 152:48]
  reg  ray_aabb_2_2_temp; // @[IST3.scala 153:48]
  reg [31:0] temp_6; // @[IST3.scala 164:50]
  reg [31:0] temp_7; // @[IST3.scala 165:50]
  reg [31:0] temp_0_2; // @[IST3.scala 166:47]
  reg [31:0] temp_0_3; // @[IST3.scala 167:47]
  reg [31:0] temp_5_2; // @[IST3.scala 168:46]
  reg [31:0] temp_5_3; // @[IST3.scala 169:46]
  reg [31:0] nodeid_ist3_temp_2; // @[IST3.scala 196:38]
  reg [31:0] rayid_ist3_temp_2; // @[IST3.scala 197:41]
  reg [31:0] t_temp_2; // @[IST3.scala 198:51]
  reg [31:0] u_temp_2; // @[IST3.scala 199:50]
  reg [31:0] hitT_temp_2; // @[IST3.scala 200:47]
  reg  enable_2; // @[IST3.scala 201:50]
  reg  break_2; // @[IST3.scala 202:51]
  reg  ray_aabb_1_2; // @[IST3.scala 203:44]
  reg  ray_aabb_2_2; // @[IST3.scala 204:43]
  reg [31:0] nodeid_ist3_temp_3_temp; // @[IST3.scala 217:43]
  reg [31:0] rayid_ist3_temp_3_temp; // @[IST3.scala 218:46]
  reg [31:0] t_temp_3_temp; // @[IST3.scala 219:56]
  reg [31:0] u_temp_3_temp; // @[IST3.scala 220:55]
  reg [31:0] hitT_temp_3_temp; // @[IST3.scala 221:52]
  reg  enable_3_temp; // @[IST3.scala 222:55]
  reg  break_3_temp; // @[IST3.scala 223:56]
  reg  ray_aabb_1_3_temp; // @[IST3.scala 224:48]
  reg  ray_aabb_2_3_temp; // @[IST3.scala 225:48]
  reg [31:0] Oy; // @[IST3.scala 235:58]
  reg [31:0] Dy; // @[IST3.scala 236:58]
  reg [31:0] nodeid_ist3_temp_3; // @[IST3.scala 258:38]
  reg [31:0] rayid_ist3_temp_3; // @[IST3.scala 259:41]
  reg [31:0] t_temp_3; // @[IST3.scala 260:51]
  reg [31:0] u_temp_3; // @[IST3.scala 261:50]
  reg [31:0] hitT_temp_3; // @[IST3.scala 262:47]
  reg  enable_3; // @[IST3.scala 263:50]
  reg  break_3; // @[IST3.scala 264:51]
  reg  ray_aabb_1_3; // @[IST3.scala 265:43]
  reg  ray_aabb_2_3; // @[IST3.scala 266:43]
  reg [31:0] nodeid_ist3_temp_4_temp; // @[IST3.scala 279:47]
  reg [31:0] rayid_ist3_temp_4_temp; // @[IST3.scala 280:50]
  reg [31:0] t_temp_4_temp; // @[IST3.scala 281:60]
  reg [31:0] u_temp_4_temp; // @[IST3.scala 282:59]
  reg [31:0] hitT_temp_4_temp; // @[IST3.scala 283:56]
  reg  enable_4_temp; // @[IST3.scala 284:59]
  reg  break_4_temp; // @[IST3.scala 285:60]
  reg  ray_aabb_1_4_temp; // @[IST3.scala 286:52]
  reg  ray_aabb_2_4_temp; // @[IST3.scala 287:52]
  reg [31:0] temp_v; // @[IST3.scala 297:67]
  reg [31:0] nodeid_ist3_temp_4; // @[IST3.scala 309:42]
  reg [31:0] rayid_ist3_temp_4; // @[IST3.scala 310:45]
  reg [31:0] t_temp_4; // @[IST3.scala 311:55]
  reg [31:0] u_temp_4; // @[IST3.scala 312:54]
  reg [31:0] hitT_temp_4; // @[IST3.scala 313:51]
  reg  enable_4; // @[IST3.scala 314:54]
  reg  break_4; // @[IST3.scala 315:55]
  reg  ray_aabb_1_4; // @[IST3.scala 316:47]
  reg  ray_aabb_2_4; // @[IST3.scala 317:47]
  reg [31:0] u_add_v; // @[IST3.scala 331:52]
  reg [31:0] nodeid_ist3_temp_5_temp; // @[IST3.scala 332:43]
  reg [31:0] rayid_ist3_temp_5_temp; // @[IST3.scala 333:46]
  reg [31:0] t_temp_5_temp; // @[IST3.scala 334:56]
  reg  v_cmp_0_0; // @[IST3.scala 335:61]
  reg [31:0] hitT_temp_5_temp; // @[IST3.scala 336:52]
  reg  enable_5_temp; // @[IST3.scala 337:55]
  reg  break_5_temp; // @[IST3.scala 339:56]
  reg  ray_aabb_1_5_temp; // @[IST3.scala 340:48]
  reg  ray_aabb_2_5_temp; // @[IST3.scala 341:48]
  wire  _T = FCMP_24_io_actual_out > 1'h0; // @[IST3.scala 355:36]
  reg  v_cmp_0; // @[IST3.scala 361:52]
  reg [31:0] nodeid_ist3_temp_5; // @[IST3.scala 377:38]
  reg [31:0] rayid_ist3_temp_5; // @[IST3.scala 378:41]
  reg [31:0] t_temp_5; // @[IST3.scala 379:51]
  reg [31:0] hitT_temp_5; // @[IST3.scala 382:47]
  reg  enable_5; // @[IST3.scala 383:50]
  reg  break_5; // @[IST3.scala 385:51]
  reg  ray_aabb_1_5; // @[IST3.scala 386:43]
  reg  ray_aabb_2_5; // @[IST3.scala 387:43]
  wire  _T_3 = FCMP_25_io_actual_out & enable_5; // @[IST3.scala 403:43]
  wire  _T_5 = FCMP_25_io_actual_out & enable_5 & v_cmp_0; // @[IST3.scala 403:61]
  wire  _T_6 = ~break_5; // @[IST3.scala 403:90]
  wire  _T_10 = ~FCMP_25_io_actual_out & enable_5; // @[IST3.scala 411:49]
  wire  _T_12 = ~FCMP_25_io_actual_out & enable_5 & v_cmp_0; // @[IST3.scala 411:67]
  wire  _T_18 = ~v_cmp_0; // @[IST3.scala 419:78]
  wire  _T_19 = _T_10 & ~v_cmp_0; // @[IST3.scala 419:67]
  wire  _T_26 = _T_3 & _T_18; // @[IST3.scala 427:67]
  wire  _T_28 = _T_3 & _T_18 & _T_6; // @[IST3.scala 427:86]
  wire  _T_35 = _T_5 & break_5; // @[IST3.scala 435:86]
  wire  _T_56 = _T_26 & break_5; // @[IST3.scala 459:86]
  wire [31:0] _GEN_1 = _T_26 & break_5 ? hitT_temp_5 : 32'h0; // @[IST3.scala 459:104 IST3.scala 460:45 IST3.scala 468:45]
  wire [32:0] _GEN_2 = _T_26 & break_5 ? $signed(33'shbf800000) : $signed(33'sh0); // @[IST3.scala 459:104 IST3.scala 461:45 IST3.scala 469:45]
  wire [31:0] _GEN_4 = _T_26 & break_5 ? rayid_ist3_temp_5 : 32'h0; // @[IST3.scala 459:104 IST3.scala 463:38 IST3.scala 471:38]
  wire [31:0] _GEN_6 = _T_19 & break_5 ? hitT_temp_5 : _GEN_1; // @[IST3.scala 451:104 IST3.scala 452:45]
  wire [32:0] _GEN_7 = _T_19 & break_5 ? $signed(33'shbf800000) : $signed(_GEN_2); // @[IST3.scala 451:104 IST3.scala 453:45]
  wire [31:0] _GEN_9 = _T_19 & break_5 ? rayid_ist3_temp_5 : _GEN_4; // @[IST3.scala 451:104 IST3.scala 455:38]
  wire  _GEN_10 = _T_19 & break_5 | _T_56; // @[IST3.scala 451:104 IST3.scala 458:41]
  wire [31:0] _GEN_11 = _T_12 & break_5 ? hitT_temp_5 : _GEN_6; // @[IST3.scala 443:104 IST3.scala 444:45]
  wire [32:0] _GEN_12 = _T_12 & break_5 ? $signed(33'shbf800000) : $signed(_GEN_7); // @[IST3.scala 443:104 IST3.scala 445:45]
  wire [31:0] _GEN_14 = _T_12 & break_5 ? rayid_ist3_temp_5 : _GEN_9; // @[IST3.scala 443:104 IST3.scala 447:38]
  wire  _GEN_15 = _T_12 & break_5 | _GEN_10; // @[IST3.scala 443:104 IST3.scala 450:41]
  wire [31:0] _GEN_16 = _T_5 & break_5 ? t_temp_5 : _GEN_11; // @[IST3.scala 435:104 IST3.scala 436:45]
  wire [32:0] _GEN_17 = _T_5 & break_5 ? $signed({{1{nodeid_ist3_temp_5[31]}},nodeid_ist3_temp_5}) : $signed(_GEN_12); // @[IST3.scala 435:104 IST3.scala 437:45]
  wire [31:0] _GEN_19 = _T_5 & break_5 ? rayid_ist3_temp_5 : _GEN_14; // @[IST3.scala 435:104 IST3.scala 439:38]
  wire  _GEN_21 = _T_5 & break_5 | _GEN_15; // @[IST3.scala 435:104 IST3.scala 442:41]
  wire [31:0] _GEN_22 = _T_3 & _T_18 & _T_6 ? hitT_temp_5 : _GEN_16; // @[IST3.scala 427:104 IST3.scala 428:45]
  wire [32:0] _GEN_23 = _T_3 & _T_18 & _T_6 ? $signed(33'shbf800000) : $signed(_GEN_17); // @[IST3.scala 427:104 IST3.scala 429:45]
  wire [31:0] _GEN_25 = _T_3 & _T_18 & _T_6 ? rayid_ist3_temp_5 : _GEN_19; // @[IST3.scala 427:104 IST3.scala 431:38]
  wire  _GEN_26 = _T_3 & _T_18 & _T_6 ? 1'h0 : _T_35; // @[IST3.scala 427:104 IST3.scala 432:45]
  wire  _GEN_27 = _T_3 & _T_18 & _T_6 ? 1'h0 : _GEN_21; // @[IST3.scala 427:104 IST3.scala 434:41]
  wire [31:0] _GEN_28 = _T_10 & ~v_cmp_0 & _T_6 ? hitT_temp_5 : _GEN_22; // @[IST3.scala 419:104 IST3.scala 420:45]
  wire [32:0] _GEN_29 = _T_10 & ~v_cmp_0 & _T_6 ? $signed(33'shbf800000) : $signed(_GEN_23); // @[IST3.scala 419:104 IST3.scala 421:45]
  wire  _GEN_30 = _T_10 & ~v_cmp_0 & _T_6 | _T_28; // @[IST3.scala 419:104 IST3.scala 422:46]
  wire [31:0] _GEN_31 = _T_10 & ~v_cmp_0 & _T_6 ? rayid_ist3_temp_5 : _GEN_25; // @[IST3.scala 419:104 IST3.scala 423:38]
  wire  _GEN_32 = _T_10 & ~v_cmp_0 & _T_6 ? 1'h0 : _GEN_26; // @[IST3.scala 419:104 IST3.scala 424:45]
  wire  _GEN_33 = _T_10 & ~v_cmp_0 & _T_6 ? 1'h0 : _GEN_27; // @[IST3.scala 419:104 IST3.scala 426:41]
  wire [31:0] _GEN_34 = ~FCMP_25_io_actual_out & enable_5 & v_cmp_0 & _T_6 ? hitT_temp_5 : _GEN_28; // @[IST3.scala 411:104 IST3.scala 412:45]
  wire [32:0] _GEN_35 = ~FCMP_25_io_actual_out & enable_5 & v_cmp_0 & _T_6 ? $signed(33'shbf800000) : $signed(_GEN_29); // @[IST3.scala 411:104 IST3.scala 413:45]
  wire  _GEN_36 = ~FCMP_25_io_actual_out & enable_5 & v_cmp_0 & _T_6 | _GEN_30; // @[IST3.scala 411:104 IST3.scala 414:46]
  wire [31:0] _GEN_37 = ~FCMP_25_io_actual_out & enable_5 & v_cmp_0 & _T_6 ? rayid_ist3_temp_5 : _GEN_31; // @[IST3.scala 411:104 IST3.scala 415:38]
  wire  _GEN_38 = ~FCMP_25_io_actual_out & enable_5 & v_cmp_0 & _T_6 ? 1'h0 : _GEN_32; // @[IST3.scala 411:104 IST3.scala 416:45]
  wire  _GEN_39 = ~FCMP_25_io_actual_out & enable_5 & v_cmp_0 & _T_6 ? 1'h0 : _GEN_33; // @[IST3.scala 411:104 IST3.scala 418:41]
  wire [32:0] _GEN_41 = FCMP_25_io_actual_out & enable_5 & v_cmp_0 & ~break_5 ? $signed({{1{nodeid_ist3_temp_5[31]}},
    nodeid_ist3_temp_5}) : $signed(_GEN_35); // @[IST3.scala 403:98 IST3.scala 405:45]
  MY_MULADD FADD_MUL_16 ( // @[IST3.scala 70:33]
    .clock(FADD_MUL_16_clock),
    .reset(FADD_MUL_16_reset),
    .io_a(FADD_MUL_16_io_a),
    .io_b(FADD_MUL_16_io_b),
    .io_c(FADD_MUL_16_io_c),
    .io_out(FADD_MUL_16_io_out)
  );
  MY_MUL FMUL_12 ( // @[IST3.scala 80:25]
    .clock(FMUL_12_clock),
    .reset(FMUL_12_reset),
    .io_a(FMUL_12_io_a),
    .io_b(FMUL_12_io_b),
    .io_out(FMUL_12_io_out)
  );
  MY_MUL FMUL_13 ( // @[IST3.scala 89:25]
    .clock(FMUL_13_clock),
    .reset(FMUL_13_reset),
    .io_a(FMUL_13_io_a),
    .io_b(FMUL_13_io_b),
    .io_out(FMUL_13_io_out)
  );
  MY_MUL FMUL_14 ( // @[IST3.scala 98:25]
    .clock(FMUL_14_clock),
    .reset(FMUL_14_reset),
    .io_a(FMUL_14_io_a),
    .io_b(FMUL_14_io_b),
    .io_out(FMUL_14_io_out)
  );
  MY_MUL FMUL_15 ( // @[IST3.scala 107:25]
    .clock(FMUL_15_clock),
    .reset(FMUL_15_reset),
    .io_a(FMUL_15_io_a),
    .io_b(FMUL_15_io_b),
    .io_out(FMUL_15_io_out)
  );
  MY_MUL FMUL_16 ( // @[IST3.scala 116:25]
    .clock(FMUL_16_clock),
    .reset(FMUL_16_reset),
    .io_a(FMUL_16_io_a),
    .io_b(FMUL_16_io_b),
    .io_out(FMUL_16_io_out)
  );
  MY_ADD FADD_9 ( // @[IST3.scala 178:24]
    .clock(FADD_9_clock),
    .reset(FADD_9_reset),
    .io_a(FADD_9_io_a),
    .io_b(FADD_9_io_b),
    .io_out(FADD_9_io_out)
  );
  MY_ADD FADD_10 ( // @[IST3.scala 187:25]
    .clock(FADD_10_clock),
    .reset(FADD_10_reset),
    .io_a(FADD_10_io_a),
    .io_b(FADD_10_io_b),
    .io_out(FADD_10_io_out)
  );
  MY_ADD FADD_11 ( // @[IST3.scala 238:25]
    .clock(FADD_11_clock),
    .reset(FADD_11_reset),
    .io_a(FADD_11_io_a),
    .io_b(FADD_11_io_b),
    .io_out(FADD_11_io_out)
  );
  MY_ADD FADD_12 ( // @[IST3.scala 247:25]
    .clock(FADD_12_clock),
    .reset(FADD_12_reset),
    .io_a(FADD_12_io_a),
    .io_b(FADD_12_io_b),
    .io_out(FADD_12_io_out)
  );
  MY_MULADD FADD_MUL_17 ( // @[IST3.scala 299:33]
    .clock(FADD_MUL_17_clock),
    .reset(FADD_MUL_17_reset),
    .io_a(FADD_MUL_17_io_a),
    .io_b(FADD_MUL_17_io_b),
    .io_c(FADD_MUL_17_io_c),
    .io_out(FADD_MUL_17_io_out)
  );
  ValExec_CompareRecF32_lt FCMP_24 ( // @[IST3.scala 350:25]
    .io_a(FCMP_24_io_a),
    .io_b(FCMP_24_io_b),
    .io_actual_out(FCMP_24_io_actual_out)
  );
  MY_ADD FADD_13 ( // @[IST3.scala 364:25]
    .clock(FADD_13_clock),
    .reset(FADD_13_reset),
    .io_a(FADD_13_io_a),
    .io_b(FADD_13_io_b),
    .io_out(FADD_13_io_out)
  );
  ValExec_CompareRecF32_le FCMP_25 ( // @[IST3.scala 398:25]
    .io_a(FCMP_25_io_a),
    .io_b(FCMP_25_io_b),
    .io_actual_out(FCMP_25_io_actual_out)
  );
  assign io_nodeid_ist3_out = nodeid_ist3_temp_5; // @[IST3.scala 397:37]
  assign io_rayid_ist3_out = FCMP_25_io_actual_out & enable_5 & v_cmp_0 & ~break_5 ? rayid_ist3_temp_5 : _GEN_37; // @[IST3.scala 403:98 IST3.scala 407:38]
  assign io_hiT_out = FCMP_25_io_actual_out & enable_5 & v_cmp_0 & ~break_5 ? t_temp_5 : _GEN_34; // @[IST3.scala 403:98 IST3.scala 404:45]
  assign io_hitT_en = FCMP_25_io_actual_out & enable_5 & v_cmp_0 & ~break_5 | _GEN_38; // @[IST3.scala 403:98 IST3.scala 408:45]
  assign io_pop_3 = FCMP_25_io_actual_out & enable_5 & v_cmp_0 & ~break_5 | _GEN_36; // @[IST3.scala 403:98 IST3.scala 406:46]
  assign io_hitIndex = _GEN_41[31:0];
  assign io_break_out = FCMP_25_io_actual_out & enable_5 & v_cmp_0 & ~break_5 ? 1'h0 : _GEN_39; // @[IST3.scala 403:98 IST3.scala 410:41]
  assign io_RAY_AABB_1_out = ray_aabb_1_5; // @[IST3.scala 476:37]
  assign io_RAY_AABB_2_out = ray_aabb_2_5; // @[IST3.scala 477:37]
  assign FADD_MUL_16_clock = clock;
  assign FADD_MUL_16_reset = reset;
  assign FADD_MUL_16_io_a = io_ray_o_in_x; // @[IST3.scala 71:26]
  assign FADD_MUL_16_io_b = io_v22_in_x; // @[IST3.scala 72:26]
  assign FADD_MUL_16_io_c = io_v22_in_w; // @[IST3.scala 73:26]
  assign FMUL_12_clock = clock;
  assign FMUL_12_reset = reset;
  assign FMUL_12_io_a = io_ray_o_in_y; // @[IST3.scala 81:22]
  assign FMUL_12_io_b = io_v22_in_y; // @[IST3.scala 82:22]
  assign FMUL_13_clock = clock;
  assign FMUL_13_reset = reset;
  assign FMUL_13_io_a = io_ray_o_in_z; // @[IST3.scala 90:22]
  assign FMUL_13_io_b = io_v22_in_z; // @[IST3.scala 91:22]
  assign FMUL_14_clock = clock;
  assign FMUL_14_reset = reset;
  assign FMUL_14_io_a = io_ray_d_in_x; // @[IST3.scala 99:22]
  assign FMUL_14_io_b = io_v22_in_x; // @[IST3.scala 100:22]
  assign FMUL_15_clock = clock;
  assign FMUL_15_reset = reset;
  assign FMUL_15_io_a = io_ray_d_in_y; // @[IST3.scala 108:22]
  assign FMUL_15_io_b = io_v22_in_y; // @[IST3.scala 109:22]
  assign FMUL_16_clock = clock;
  assign FMUL_16_reset = reset;
  assign FMUL_16_io_a = io_ray_d_in_z; // @[IST3.scala 117:22]
  assign FMUL_16_io_b = io_v22_in_z; // @[IST3.scala 118:22]
  assign FADD_9_clock = clock;
  assign FADD_9_reset = reset;
  assign FADD_9_io_a = temp_1; // @[IST3.scala 179:21]
  assign FADD_9_io_b = temp_2; // @[IST3.scala 180:21]
  assign FADD_10_clock = clock;
  assign FADD_10_reset = reset;
  assign FADD_10_io_a = temp_3; // @[IST3.scala 188:22]
  assign FADD_10_io_b = temp_4; // @[IST3.scala 189:22]
  assign FADD_11_clock = clock;
  assign FADD_11_reset = reset;
  assign FADD_11_io_a = temp_0_3; // @[IST3.scala 239:22]
  assign FADD_11_io_b = temp_6; // @[IST3.scala 240:22]
  assign FADD_12_clock = clock;
  assign FADD_12_reset = reset;
  assign FADD_12_io_a = temp_5_3; // @[IST3.scala 248:22]
  assign FADD_12_io_b = temp_7; // @[IST3.scala 249:22]
  assign FADD_MUL_17_clock = clock;
  assign FADD_MUL_17_reset = reset;
  assign FADD_MUL_17_io_a = t_temp_3; // @[IST3.scala 300:26]
  assign FADD_MUL_17_io_b = Dy; // @[IST3.scala 301:26]
  assign FADD_MUL_17_io_c = Oy; // @[IST3.scala 302:26]
  assign FCMP_24_io_a = 32'h0; // @[IST3.scala 351:22]
  assign FCMP_24_io_b = temp_v; // @[IST3.scala 352:22]
  assign FADD_13_clock = clock;
  assign FADD_13_reset = reset;
  assign FADD_13_io_a = temp_v; // @[IST3.scala 365:22]
  assign FADD_13_io_b = u_temp_4; // @[IST3.scala 366:22]
  assign FCMP_25_io_a = u_add_v; // @[IST3.scala 399:22]
  assign FCMP_25_io_b = 32'h3f800000; // @[IST3.scala 400:22]
  always @(posedge clock) begin
    if (reset) begin // @[IST3.scala 44:33]
      temp_0 <= 32'h0; // @[IST3.scala 44:33]
    end else begin
      temp_0 <= FADD_MUL_16_io_out; // @[IST3.scala 78:42]
    end
    if (reset) begin // @[IST3.scala 45:33]
      temp_1 <= 32'h0; // @[IST3.scala 45:33]
    end else begin
      temp_1 <= FMUL_12_io_out; // @[IST3.scala 87:42]
    end
    if (reset) begin // @[IST3.scala 46:33]
      temp_2 <= 32'h0; // @[IST3.scala 46:33]
    end else begin
      temp_2 <= FMUL_13_io_out; // @[IST3.scala 96:42]
    end
    if (reset) begin // @[IST3.scala 47:33]
      temp_3 <= 32'h0; // @[IST3.scala 47:33]
    end else begin
      temp_3 <= FMUL_14_io_out; // @[IST3.scala 105:42]
    end
    if (reset) begin // @[IST3.scala 48:33]
      temp_4 <= 32'h0; // @[IST3.scala 48:33]
    end else begin
      temp_4 <= FMUL_15_io_out; // @[IST3.scala 114:42]
    end
    if (reset) begin // @[IST3.scala 49:33]
      temp_5 <= 32'h0; // @[IST3.scala 49:33]
    end else begin
      temp_5 <= FMUL_16_io_out; // @[IST3.scala 123:42]
    end
    if (reset) begin // @[IST3.scala 51:42]
      nodeid_ist3_temp_1_temp <= 32'sh0; // @[IST3.scala 51:42]
    end else begin
      nodeid_ist3_temp_1_temp <= io_nodeid_leaf_3; // @[IST3.scala 60:34]
    end
    if (reset) begin // @[IST3.scala 52:46]
      rayid_ist3_temp_1_temp <= 32'h0; // @[IST3.scala 52:46]
    end else begin
      rayid_ist3_temp_1_temp <= io_rayid_leaf_3; // @[IST3.scala 61:37]
    end
    if (reset) begin // @[IST3.scala 53:56]
      t_temp_1_temp <= 32'h0; // @[IST3.scala 53:56]
    end else begin
      t_temp_1_temp <= io_t_in; // @[IST3.scala 62:47]
    end
    if (reset) begin // @[IST3.scala 54:54]
      u_temp_1_temp <= 32'h0; // @[IST3.scala 54:54]
    end else begin
      u_temp_1_temp <= io_u_in; // @[IST3.scala 63:46]
    end
    if (reset) begin // @[IST3.scala 55:52]
      hitT_temp_1_temp <= 32'h0; // @[IST3.scala 55:52]
    end else begin
      hitT_temp_1_temp <= io_hiT_in; // @[IST3.scala 64:43]
    end
    if (reset) begin // @[IST3.scala 56:55]
      enable_1_temp <= 1'h0; // @[IST3.scala 56:55]
    end else begin
      enable_1_temp <= io_enable_IST3; // @[IST3.scala 65:48]
    end
    if (reset) begin // @[IST3.scala 57:56]
      break_1_temp <= 1'h0; // @[IST3.scala 57:56]
    end else begin
      break_1_temp <= io_break_in; // @[IST3.scala 66:50]
    end
    if (reset) begin // @[IST3.scala 58:51]
      ray_aabb_1_temp <= 1'h0; // @[IST3.scala 58:51]
    end else begin
      ray_aabb_1_temp <= io_RAY_AABB_1; // @[IST3.scala 67:45]
    end
    if (reset) begin // @[IST3.scala 59:51]
      ray_aabb_2_temp <= 1'h0; // @[IST3.scala 59:51]
    end else begin
      ray_aabb_2_temp <= io_RAY_AABB_2; // @[IST3.scala 68:45]
    end
    if (reset) begin // @[IST3.scala 126:37]
      nodeid_ist3_temp_1 <= 32'sh0; // @[IST3.scala 126:37]
    end else begin
      nodeid_ist3_temp_1 <= nodeid_ist3_temp_1_temp; // @[IST3.scala 135:29]
    end
    if (reset) begin // @[IST3.scala 127:41]
      rayid_ist3_temp_1 <= 32'h0; // @[IST3.scala 127:41]
    end else begin
      rayid_ist3_temp_1 <= rayid_ist3_temp_1_temp; // @[IST3.scala 136:32]
    end
    if (reset) begin // @[IST3.scala 128:51]
      t_temp_1 <= 32'h0; // @[IST3.scala 128:51]
    end else begin
      t_temp_1 <= t_temp_1_temp; // @[IST3.scala 137:42]
    end
    if (reset) begin // @[IST3.scala 129:49]
      u_temp_1 <= 32'h0; // @[IST3.scala 129:49]
    end else begin
      u_temp_1 <= u_temp_1_temp; // @[IST3.scala 138:41]
    end
    if (reset) begin // @[IST3.scala 130:47]
      hitT_temp_1 <= 32'h0; // @[IST3.scala 130:47]
    end else begin
      hitT_temp_1 <= hitT_temp_1_temp; // @[IST3.scala 139:38]
    end
    if (reset) begin // @[IST3.scala 131:50]
      enable_1 <= 1'h0; // @[IST3.scala 131:50]
    end else begin
      enable_1 <= enable_1_temp; // @[IST3.scala 140:43]
    end
    if (reset) begin // @[IST3.scala 132:51]
      break_1 <= 1'h0; // @[IST3.scala 132:51]
    end else begin
      break_1 <= break_1_temp; // @[IST3.scala 141:45]
    end
    if (reset) begin // @[IST3.scala 133:46]
      ray_aabb_1 <= 1'h0; // @[IST3.scala 133:46]
    end else begin
      ray_aabb_1 <= ray_aabb_1_temp; // @[IST3.scala 142:40]
    end
    if (reset) begin // @[IST3.scala 134:46]
      ray_aabb_2 <= 1'h0; // @[IST3.scala 134:46]
    end else begin
      ray_aabb_2 <= ray_aabb_2_temp; // @[IST3.scala 143:40]
    end
    if (reset) begin // @[IST3.scala 145:43]
      nodeid_ist3_temp_2_temp <= 32'sh0; // @[IST3.scala 145:43]
    end else begin
      nodeid_ist3_temp_2_temp <= nodeid_ist3_temp_1; // @[IST3.scala 154:34]
    end
    if (reset) begin // @[IST3.scala 146:46]
      rayid_ist3_temp_2_temp <= 32'h0; // @[IST3.scala 146:46]
    end else begin
      rayid_ist3_temp_2_temp <= rayid_ist3_temp_1; // @[IST3.scala 155:37]
    end
    if (reset) begin // @[IST3.scala 147:56]
      t_temp_2_temp <= 32'h0; // @[IST3.scala 147:56]
    end else begin
      t_temp_2_temp <= t_temp_1; // @[IST3.scala 156:46]
    end
    if (reset) begin // @[IST3.scala 148:55]
      u_temp_2_temp <= 32'h0; // @[IST3.scala 148:55]
    end else begin
      u_temp_2_temp <= u_temp_1; // @[IST3.scala 157:45]
    end
    if (reset) begin // @[IST3.scala 149:52]
      hitT_temp_2_temp <= 32'h0; // @[IST3.scala 149:52]
    end else begin
      hitT_temp_2_temp <= hitT_temp_1; // @[IST3.scala 158:43]
    end
    if (reset) begin // @[IST3.scala 150:55]
      enable_2_temp <= 1'h0; // @[IST3.scala 150:55]
    end else begin
      enable_2_temp <= enable_1; // @[IST3.scala 159:47]
    end
    if (reset) begin // @[IST3.scala 151:56]
      break_2_temp <= 1'h0; // @[IST3.scala 151:56]
    end else begin
      break_2_temp <= break_1; // @[IST3.scala 160:48]
    end
    if (reset) begin // @[IST3.scala 152:48]
      ray_aabb_1_2_temp <= 1'h0; // @[IST3.scala 152:48]
    end else begin
      ray_aabb_1_2_temp <= ray_aabb_1; // @[IST3.scala 161:40]
    end
    if (reset) begin // @[IST3.scala 153:48]
      ray_aabb_2_2_temp <= 1'h0; // @[IST3.scala 153:48]
    end else begin
      ray_aabb_2_2_temp <= ray_aabb_2; // @[IST3.scala 162:40]
    end
    if (reset) begin // @[IST3.scala 164:50]
      temp_6 <= 32'h0; // @[IST3.scala 164:50]
    end else begin
      temp_6 <= FADD_9_io_out; // @[IST3.scala 185:26]
    end
    if (reset) begin // @[IST3.scala 165:50]
      temp_7 <= 32'h0; // @[IST3.scala 165:50]
    end else begin
      temp_7 <= FADD_10_io_out; // @[IST3.scala 194:26]
    end
    if (reset) begin // @[IST3.scala 166:47]
      temp_0_2 <= 32'h0; // @[IST3.scala 166:47]
    end else begin
      temp_0_2 <= temp_0; // @[IST3.scala 175:41]
    end
    if (reset) begin // @[IST3.scala 167:47]
      temp_0_3 <= 32'h0; // @[IST3.scala 167:47]
    end else begin
      temp_0_3 <= temp_0_2; // @[IST3.scala 172:41]
    end
    if (reset) begin // @[IST3.scala 168:46]
      temp_5_2 <= 32'h0; // @[IST3.scala 168:46]
    end else begin
      temp_5_2 <= temp_5; // @[IST3.scala 176:41]
    end
    if (reset) begin // @[IST3.scala 169:46]
      temp_5_3 <= 32'h0; // @[IST3.scala 169:46]
    end else begin
      temp_5_3 <= temp_5_2; // @[IST3.scala 174:41]
    end
    if (reset) begin // @[IST3.scala 196:38]
      nodeid_ist3_temp_2 <= 32'sh0; // @[IST3.scala 196:38]
    end else begin
      nodeid_ist3_temp_2 <= nodeid_ist3_temp_2_temp; // @[IST3.scala 205:29]
    end
    if (reset) begin // @[IST3.scala 197:41]
      rayid_ist3_temp_2 <= 32'h0; // @[IST3.scala 197:41]
    end else begin
      rayid_ist3_temp_2 <= rayid_ist3_temp_2_temp; // @[IST3.scala 206:32]
    end
    if (reset) begin // @[IST3.scala 198:51]
      t_temp_2 <= 32'h0; // @[IST3.scala 198:51]
    end else begin
      t_temp_2 <= t_temp_2_temp; // @[IST3.scala 207:41]
    end
    if (reset) begin // @[IST3.scala 199:50]
      u_temp_2 <= 32'h0; // @[IST3.scala 199:50]
    end else begin
      u_temp_2 <= u_temp_2_temp; // @[IST3.scala 208:40]
    end
    if (reset) begin // @[IST3.scala 200:47]
      hitT_temp_2 <= 32'h0; // @[IST3.scala 200:47]
    end else begin
      hitT_temp_2 <= hitT_temp_2_temp; // @[IST3.scala 209:38]
    end
    if (reset) begin // @[IST3.scala 201:50]
      enable_2 <= 1'h0; // @[IST3.scala 201:50]
    end else begin
      enable_2 <= enable_2_temp; // @[IST3.scala 210:42]
    end
    if (reset) begin // @[IST3.scala 202:51]
      break_2 <= 1'h0; // @[IST3.scala 202:51]
    end else begin
      break_2 <= break_2_temp; // @[IST3.scala 211:43]
    end
    if (reset) begin // @[IST3.scala 203:44]
      ray_aabb_1_2 <= 1'h0; // @[IST3.scala 203:44]
    end else begin
      ray_aabb_1_2 <= ray_aabb_1_2_temp; // @[IST3.scala 212:37]
    end
    if (reset) begin // @[IST3.scala 204:43]
      ray_aabb_2_2 <= 1'h0; // @[IST3.scala 204:43]
    end else begin
      ray_aabb_2_2 <= ray_aabb_2_2_temp; // @[IST3.scala 213:37]
    end
    if (reset) begin // @[IST3.scala 217:43]
      nodeid_ist3_temp_3_temp <= 32'sh0; // @[IST3.scala 217:43]
    end else begin
      nodeid_ist3_temp_3_temp <= nodeid_ist3_temp_2; // @[IST3.scala 226:37]
    end
    if (reset) begin // @[IST3.scala 218:46]
      rayid_ist3_temp_3_temp <= 32'h0; // @[IST3.scala 218:46]
    end else begin
      rayid_ist3_temp_3_temp <= rayid_ist3_temp_2; // @[IST3.scala 227:40]
    end
    if (reset) begin // @[IST3.scala 219:56]
      t_temp_3_temp <= 32'h0; // @[IST3.scala 219:56]
    end else begin
      t_temp_3_temp <= t_temp_2; // @[IST3.scala 228:50]
    end
    if (reset) begin // @[IST3.scala 220:55]
      u_temp_3_temp <= 32'h0; // @[IST3.scala 220:55]
    end else begin
      u_temp_3_temp <= u_temp_2; // @[IST3.scala 229:49]
    end
    if (reset) begin // @[IST3.scala 221:52]
      hitT_temp_3_temp <= 32'h0; // @[IST3.scala 221:52]
    end else begin
      hitT_temp_3_temp <= hitT_temp_2; // @[IST3.scala 230:46]
    end
    if (reset) begin // @[IST3.scala 222:55]
      enable_3_temp <= 1'h0; // @[IST3.scala 222:55]
    end else begin
      enable_3_temp <= enable_2; // @[IST3.scala 231:51]
    end
    if (reset) begin // @[IST3.scala 223:56]
      break_3_temp <= 1'h0; // @[IST3.scala 223:56]
    end else begin
      break_3_temp <= break_2; // @[IST3.scala 232:53]
    end
    if (reset) begin // @[IST3.scala 224:48]
      ray_aabb_1_3_temp <= 1'h0; // @[IST3.scala 224:48]
    end else begin
      ray_aabb_1_3_temp <= ray_aabb_1_2; // @[IST3.scala 233:45]
    end
    if (reset) begin // @[IST3.scala 225:48]
      ray_aabb_2_3_temp <= 1'h0; // @[IST3.scala 225:48]
    end else begin
      ray_aabb_2_3_temp <= ray_aabb_2_2; // @[IST3.scala 234:45]
    end
    if (reset) begin // @[IST3.scala 235:58]
      Oy <= 32'h0; // @[IST3.scala 235:58]
    end else begin
      Oy <= FADD_11_io_out; // @[IST3.scala 245:26]
    end
    if (reset) begin // @[IST3.scala 236:58]
      Dy <= 32'h0; // @[IST3.scala 236:58]
    end else begin
      Dy <= FADD_12_io_out; // @[IST3.scala 254:26]
    end
    if (reset) begin // @[IST3.scala 258:38]
      nodeid_ist3_temp_3 <= 32'sh0; // @[IST3.scala 258:38]
    end else begin
      nodeid_ist3_temp_3 <= nodeid_ist3_temp_3_temp; // @[IST3.scala 267:32]
    end
    if (reset) begin // @[IST3.scala 259:41]
      rayid_ist3_temp_3 <= 32'h0; // @[IST3.scala 259:41]
    end else begin
      rayid_ist3_temp_3 <= rayid_ist3_temp_3_temp; // @[IST3.scala 268:35]
    end
    if (reset) begin // @[IST3.scala 260:51]
      t_temp_3 <= 32'h0; // @[IST3.scala 260:51]
    end else begin
      t_temp_3 <= t_temp_3_temp; // @[IST3.scala 269:45]
    end
    if (reset) begin // @[IST3.scala 261:50]
      u_temp_3 <= 32'h0; // @[IST3.scala 261:50]
    end else begin
      u_temp_3 <= u_temp_3_temp; // @[IST3.scala 270:44]
    end
    if (reset) begin // @[IST3.scala 262:47]
      hitT_temp_3 <= 32'h0; // @[IST3.scala 262:47]
    end else begin
      hitT_temp_3 <= hitT_temp_3_temp; // @[IST3.scala 271:41]
    end
    if (reset) begin // @[IST3.scala 263:50]
      enable_3 <= 1'h0; // @[IST3.scala 263:50]
    end else begin
      enable_3 <= enable_3_temp; // @[IST3.scala 272:43]
    end
    if (reset) begin // @[IST3.scala 264:51]
      break_3 <= 1'h0; // @[IST3.scala 264:51]
    end else begin
      break_3 <= break_3_temp; // @[IST3.scala 273:45]
    end
    if (reset) begin // @[IST3.scala 265:43]
      ray_aabb_1_3 <= 1'h0; // @[IST3.scala 265:43]
    end else begin
      ray_aabb_1_3 <= ray_aabb_1_3_temp; // @[IST3.scala 274:37]
    end
    if (reset) begin // @[IST3.scala 266:43]
      ray_aabb_2_3 <= 1'h0; // @[IST3.scala 266:43]
    end else begin
      ray_aabb_2_3 <= ray_aabb_2_3_temp; // @[IST3.scala 275:37]
    end
    if (reset) begin // @[IST3.scala 279:47]
      nodeid_ist3_temp_4_temp <= 32'sh0; // @[IST3.scala 279:47]
    end else begin
      nodeid_ist3_temp_4_temp <= nodeid_ist3_temp_3; // @[IST3.scala 288:41]
    end
    if (reset) begin // @[IST3.scala 280:50]
      rayid_ist3_temp_4_temp <= 32'h0; // @[IST3.scala 280:50]
    end else begin
      rayid_ist3_temp_4_temp <= rayid_ist3_temp_3; // @[IST3.scala 289:44]
    end
    if (reset) begin // @[IST3.scala 281:60]
      t_temp_4_temp <= 32'h0; // @[IST3.scala 281:60]
    end else begin
      t_temp_4_temp <= t_temp_3; // @[IST3.scala 290:54]
    end
    if (reset) begin // @[IST3.scala 282:59]
      u_temp_4_temp <= 32'h0; // @[IST3.scala 282:59]
    end else begin
      u_temp_4_temp <= u_temp_3; // @[IST3.scala 291:53]
    end
    if (reset) begin // @[IST3.scala 283:56]
      hitT_temp_4_temp <= 32'h0; // @[IST3.scala 283:56]
    end else begin
      hitT_temp_4_temp <= hitT_temp_3; // @[IST3.scala 292:50]
    end
    if (reset) begin // @[IST3.scala 284:59]
      enable_4_temp <= 1'h0; // @[IST3.scala 284:59]
    end else begin
      enable_4_temp <= enable_3; // @[IST3.scala 293:55]
    end
    if (reset) begin // @[IST3.scala 285:60]
      break_4_temp <= 1'h0; // @[IST3.scala 285:60]
    end else begin
      break_4_temp <= break_3; // @[IST3.scala 294:56]
    end
    if (reset) begin // @[IST3.scala 286:52]
      ray_aabb_1_4_temp <= 1'h0; // @[IST3.scala 286:52]
    end else begin
      ray_aabb_1_4_temp <= ray_aabb_1_3; // @[IST3.scala 295:48]
    end
    if (reset) begin // @[IST3.scala 287:52]
      ray_aabb_2_4_temp <= 1'h0; // @[IST3.scala 287:52]
    end else begin
      ray_aabb_2_4_temp <= ray_aabb_2_3; // @[IST3.scala 296:48]
    end
    if (reset) begin // @[IST3.scala 297:67]
      temp_v <= 32'h0; // @[IST3.scala 297:67]
    end else begin
      temp_v <= FADD_MUL_17_io_out; // @[IST3.scala 307:42]
    end
    if (reset) begin // @[IST3.scala 309:42]
      nodeid_ist3_temp_4 <= 32'sh0; // @[IST3.scala 309:42]
    end else begin
      nodeid_ist3_temp_4 <= nodeid_ist3_temp_4_temp; // @[IST3.scala 318:36]
    end
    if (reset) begin // @[IST3.scala 310:45]
      rayid_ist3_temp_4 <= 32'h0; // @[IST3.scala 310:45]
    end else begin
      rayid_ist3_temp_4 <= rayid_ist3_temp_4_temp; // @[IST3.scala 319:39]
    end
    if (reset) begin // @[IST3.scala 311:55]
      t_temp_4 <= 32'h0; // @[IST3.scala 311:55]
    end else begin
      t_temp_4 <= t_temp_4_temp; // @[IST3.scala 320:49]
    end
    if (reset) begin // @[IST3.scala 312:54]
      u_temp_4 <= 32'h0; // @[IST3.scala 312:54]
    end else begin
      u_temp_4 <= u_temp_4_temp; // @[IST3.scala 321:48]
    end
    if (reset) begin // @[IST3.scala 313:51]
      hitT_temp_4 <= 32'h0; // @[IST3.scala 313:51]
    end else begin
      hitT_temp_4 <= hitT_temp_4_temp; // @[IST3.scala 322:45]
    end
    if (reset) begin // @[IST3.scala 314:54]
      enable_4 <= 1'h0; // @[IST3.scala 314:54]
    end else begin
      enable_4 <= enable_4_temp; // @[IST3.scala 323:50]
    end
    if (reset) begin // @[IST3.scala 315:55]
      break_4 <= 1'h0; // @[IST3.scala 315:55]
    end else begin
      break_4 <= break_4_temp; // @[IST3.scala 324:51]
    end
    if (reset) begin // @[IST3.scala 316:47]
      ray_aabb_1_4 <= 1'h0; // @[IST3.scala 316:47]
    end else begin
      ray_aabb_1_4 <= ray_aabb_1_4_temp; // @[IST3.scala 325:44]
    end
    if (reset) begin // @[IST3.scala 317:47]
      ray_aabb_2_4 <= 1'h0; // @[IST3.scala 317:47]
    end else begin
      ray_aabb_2_4 <= ray_aabb_2_4_temp; // @[IST3.scala 326:44]
    end
    if (reset) begin // @[IST3.scala 331:52]
      u_add_v <= 32'h0; // @[IST3.scala 331:52]
    end else begin
      u_add_v <= FADD_13_io_out; // @[IST3.scala 371:25]
    end
    if (reset) begin // @[IST3.scala 332:43]
      nodeid_ist3_temp_5_temp <= 32'sh0; // @[IST3.scala 332:43]
    end else begin
      nodeid_ist3_temp_5_temp <= nodeid_ist3_temp_4; // @[IST3.scala 342:37]
    end
    if (reset) begin // @[IST3.scala 333:46]
      rayid_ist3_temp_5_temp <= 32'h0; // @[IST3.scala 333:46]
    end else begin
      rayid_ist3_temp_5_temp <= rayid_ist3_temp_4; // @[IST3.scala 343:40]
    end
    if (reset) begin // @[IST3.scala 334:56]
      t_temp_5_temp <= 32'h0; // @[IST3.scala 334:56]
    end else begin
      t_temp_5_temp <= t_temp_4; // @[IST3.scala 344:50]
    end
    if (reset) begin // @[IST3.scala 335:61]
      v_cmp_0_0 <= 1'h0; // @[IST3.scala 335:61]
    end else begin
      v_cmp_0_0 <= _T;
    end
    if (reset) begin // @[IST3.scala 336:52]
      hitT_temp_5_temp <= 32'h0; // @[IST3.scala 336:52]
    end else begin
      hitT_temp_5_temp <= hitT_temp_4; // @[IST3.scala 345:46]
    end
    if (reset) begin // @[IST3.scala 337:55]
      enable_5_temp <= 1'h0; // @[IST3.scala 337:55]
    end else begin
      enable_5_temp <= enable_4; // @[IST3.scala 346:51]
    end
    if (reset) begin // @[IST3.scala 339:56]
      break_5_temp <= 1'h0; // @[IST3.scala 339:56]
    end else begin
      break_5_temp <= break_4; // @[IST3.scala 347:52]
    end
    if (reset) begin // @[IST3.scala 340:48]
      ray_aabb_1_5_temp <= 1'h0; // @[IST3.scala 340:48]
    end else begin
      ray_aabb_1_5_temp <= ray_aabb_1_4; // @[IST3.scala 348:42]
    end
    if (reset) begin // @[IST3.scala 341:48]
      ray_aabb_2_5_temp <= 1'h0; // @[IST3.scala 341:48]
    end else begin
      ray_aabb_2_5_temp <= ray_aabb_2_4; // @[IST3.scala 349:42]
    end
    if (reset) begin // @[IST3.scala 361:52]
      v_cmp_0 <= 1'h0; // @[IST3.scala 361:52]
    end else begin
      v_cmp_0 <= v_cmp_0_0; // @[IST3.scala 362:45]
    end
    if (reset) begin // @[IST3.scala 377:38]
      nodeid_ist3_temp_5 <= 32'sh0; // @[IST3.scala 377:38]
    end else begin
      nodeid_ist3_temp_5 <= nodeid_ist3_temp_5_temp; // @[IST3.scala 389:32]
    end
    if (reset) begin // @[IST3.scala 378:41]
      rayid_ist3_temp_5 <= 32'h0; // @[IST3.scala 378:41]
    end else begin
      rayid_ist3_temp_5 <= rayid_ist3_temp_5_temp; // @[IST3.scala 390:35]
    end
    if (reset) begin // @[IST3.scala 379:51]
      t_temp_5 <= 32'h0; // @[IST3.scala 379:51]
    end else begin
      t_temp_5 <= t_temp_5_temp; // @[IST3.scala 391:45]
    end
    if (reset) begin // @[IST3.scala 382:47]
      hitT_temp_5 <= 32'h0; // @[IST3.scala 382:47]
    end else begin
      hitT_temp_5 <= hitT_temp_5_temp; // @[IST3.scala 392:41]
    end
    if (reset) begin // @[IST3.scala 383:50]
      enable_5 <= 1'h0; // @[IST3.scala 383:50]
    end else begin
      enable_5 <= enable_5_temp; // @[IST3.scala 393:46]
    end
    if (reset) begin // @[IST3.scala 385:51]
      break_5 <= 1'h0; // @[IST3.scala 385:51]
    end else begin
      break_5 <= break_5_temp; // @[IST3.scala 394:47]
    end
    if (reset) begin // @[IST3.scala 386:43]
      ray_aabb_1_5 <= 1'h0; // @[IST3.scala 386:43]
    end else begin
      ray_aabb_1_5 <= ray_aabb_1_5_temp; // @[IST3.scala 395:40]
    end
    if (reset) begin // @[IST3.scala 387:43]
      ray_aabb_2_5 <= 1'h0; // @[IST3.scala 387:43]
    end else begin
      ray_aabb_2_5 <= ray_aabb_2_5_temp; // @[IST3.scala 396:40]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  temp_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  temp_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  temp_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  temp_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  temp_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  temp_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  nodeid_ist3_temp_1_temp = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  rayid_ist3_temp_1_temp = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  t_temp_1_temp = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  u_temp_1_temp = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  hitT_temp_1_temp = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  enable_1_temp = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  break_1_temp = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  ray_aabb_1_temp = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  ray_aabb_2_temp = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  nodeid_ist3_temp_1 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  rayid_ist3_temp_1 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  t_temp_1 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  u_temp_1 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  hitT_temp_1 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  enable_1 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  break_1 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  ray_aabb_1 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  ray_aabb_2 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  nodeid_ist3_temp_2_temp = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  rayid_ist3_temp_2_temp = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  t_temp_2_temp = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  u_temp_2_temp = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  hitT_temp_2_temp = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  enable_2_temp = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  break_2_temp = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  ray_aabb_1_2_temp = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  ray_aabb_2_2_temp = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  temp_6 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  temp_7 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  temp_0_2 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  temp_0_3 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  temp_5_2 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  temp_5_3 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  nodeid_ist3_temp_2 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  rayid_ist3_temp_2 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  t_temp_2 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  u_temp_2 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  hitT_temp_2 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  enable_2 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  break_2 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  ray_aabb_1_2 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  ray_aabb_2_2 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  nodeid_ist3_temp_3_temp = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  rayid_ist3_temp_3_temp = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  t_temp_3_temp = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  u_temp_3_temp = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  hitT_temp_3_temp = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  enable_3_temp = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  break_3_temp = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  ray_aabb_1_3_temp = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  ray_aabb_2_3_temp = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  Oy = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  Dy = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  nodeid_ist3_temp_3 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  rayid_ist3_temp_3 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  t_temp_3 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  u_temp_3 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  hitT_temp_3 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  enable_3 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  break_3 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  ray_aabb_1_3 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  ray_aabb_2_3 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  nodeid_ist3_temp_4_temp = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  rayid_ist3_temp_4_temp = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  t_temp_4_temp = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  u_temp_4_temp = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  hitT_temp_4_temp = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  enable_4_temp = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  break_4_temp = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  ray_aabb_1_4_temp = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  ray_aabb_2_4_temp = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  temp_v = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  nodeid_ist3_temp_4 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  rayid_ist3_temp_4 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  t_temp_4 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  u_temp_4 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  hitT_temp_4 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  enable_4 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  break_4 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  ray_aabb_1_4 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  ray_aabb_2_4 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  u_add_v = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  nodeid_ist3_temp_5_temp = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  rayid_ist3_temp_5_temp = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  t_temp_5_temp = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  v_cmp_0_0 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  hitT_temp_5_temp = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  enable_5_temp = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  break_5_temp = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  ray_aabb_1_5_temp = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  ray_aabb_2_5_temp = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  v_cmp_0 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  nodeid_ist3_temp_5 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  rayid_ist3_temp_5 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  t_temp_5 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  hitT_temp_5 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  enable_5 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  break_5 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  ray_aabb_1_5 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  ray_aabb_2_5 = _RAND_105[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Triangle(
  input         clock,
  input         reset,
  input         io_To_IST0_enable,
  input  [31:0] io_nodeid_leaf,
  input  [31:0] io_rayid_leaf,
  input  [31:0] io_hiT_in,
  input  [31:0] io_v00_in_x,
  input  [31:0] io_v00_in_y,
  input  [31:0] io_v00_in_z,
  input  [31:0] io_v00_in_w,
  input  [31:0] io_v11_in_x,
  input  [31:0] io_v11_in_y,
  input  [31:0] io_v11_in_z,
  input  [31:0] io_v11_in_w,
  input  [31:0] io_v22_in_x,
  input  [31:0] io_v22_in_y,
  input  [31:0] io_v22_in_z,
  input  [31:0] io_v22_in_w,
  input  [31:0] io_ray_o_in_x,
  input  [31:0] io_ray_o_in_y,
  input  [31:0] io_ray_o_in_z,
  input  [31:0] io_ray_d_in_x,
  input  [31:0] io_ray_d_in_y,
  input  [31:0] io_ray_d_in_z,
  input         io_break_in,
  input         io_RAY_AABB_1,
  input         io_RAY_AABB_2,
  output        io_pop_1,
  output        io_break_1,
  output        io_pop_2,
  output        io_break_2,
  output        io_pop_3,
  output        io_break_3,
  output [31:0] io_hiT_out_1,
  output [31:0] io_hiT_out_2,
  output [31:0] io_hiT_out_3,
  output        io_hitT_en,
  output [31:0] io_hitIndex,
  output [31:0] io_node_id_out_1,
  output [31:0] io_node_id_out_2,
  output [31:0] io_node_id_out_3,
  output [31:0] io_ray_id_ist1,
  output [31:0] io_ray_id_ist2,
  output [31:0] io_ray_id_ist3,
  output [63:0] io_counter_fdiv,
  output        io_RAY_AABB_1_out_IST1,
  output        io_RAY_AABB_2_out_IST1,
  output        io_RAY_AABB_1_out_IST2,
  output        io_RAY_AABB_2_out_IST2,
  output        io_RAY_AABB_1_out_IST3,
  output        io_RAY_AABB_2_out_IST3
);
  wire  IST0_clock; // @[Triangle.scala 52:49]
  wire  IST0_reset; // @[Triangle.scala 52:49]
  wire  IST0_io_enable_IST0; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_nodeid_leaf; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_rayid_leaf; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_hiT_in; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_v00_x; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_v00_y; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_v00_z; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_v00_w; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_v11_in_x; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_v11_in_y; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_v11_in_z; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_v11_in_w; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_v22_in_x; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_v22_in_y; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_v22_in_z; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_v22_in_w; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_ray_o_in_x; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_ray_o_in_y; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_ray_o_in_z; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_ray_d_in_x; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_ray_d_in_y; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_ray_d_in_z; // @[Triangle.scala 52:49]
  wire  IST0_io_RAY_AABB_1; // @[Triangle.scala 52:49]
  wire  IST0_io_RAY_AABB_2; // @[Triangle.scala 52:49]
  wire  IST0_io_break_in; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_Oz; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_invDz_div; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_nodeid_ist0_out; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_rayid_ist0_out; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_hiT_out; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_v11_out_x; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_v11_out_y; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_v11_out_z; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_v11_out_w; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_v22_out_x; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_v22_out_y; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_v22_out_z; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_v22_out_w; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_ray_o_out_x; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_ray_o_out_y; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_ray_o_out_z; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_ray_d_out_x; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_ray_d_out_y; // @[Triangle.scala 52:49]
  wire [31:0] IST0_io_ray_d_out_z; // @[Triangle.scala 52:49]
  wire  IST0_io_enable_SU_out; // @[Triangle.scala 52:49]
  wire  IST0_io_break_out; // @[Triangle.scala 52:49]
  wire  IST0_io_RAY_AABB_1_out; // @[Triangle.scala 52:49]
  wire  IST0_io_RAY_AABB_2_out; // @[Triangle.scala 52:49]
  wire  SU_clock; // @[Triangle.scala 53:50]
  wire  SU_reset; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_invDz_div; // @[Triangle.scala 53:50]
  wire  SU_io_valid_in; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_v11_x; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_v11_y; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_v11_z; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_v11_w; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_v22_x; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_v22_y; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_v22_z; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_v22_w; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_ray_in; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_Oz; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_ray_o_in_x; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_ray_o_in_y; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_ray_o_in_z; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_ray_d_in_x; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_ray_d_in_y; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_ray_d_in_z; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_node_id_in; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_hitT_in; // @[Triangle.scala 53:50]
  wire  SU_io_break_in; // @[Triangle.scala 53:50]
  wire  SU_io_RAY_AABB_1; // @[Triangle.scala 53:50]
  wire  SU_io_RAY_AABB_2; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_fdiv_out; // @[Triangle.scala 53:50]
  wire  SU_io_valid_out; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_v11_out_x; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_v11_out_y; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_v11_out_z; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_v11_out_w; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_v22_out_x; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_v22_out_y; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_v22_out_z; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_v22_out_w; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_ray_out; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_Oz_out; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_ray_o_out_x; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_ray_o_out_y; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_ray_o_out_z; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_ray_d_out_x; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_ray_d_out_y; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_ray_d_out_z; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_node_id_out; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_hitT_out; // @[Triangle.scala 53:50]
  wire [31:0] SU_io_counter_fdiv; // @[Triangle.scala 53:50]
  wire  SU_io_break_out; // @[Triangle.scala 53:50]
  wire  SU_io_RAY_AABB_1_out; // @[Triangle.scala 53:50]
  wire  SU_io_RAY_AABB_2_out; // @[Triangle.scala 53:50]
  wire  IST1_clock; // @[Triangle.scala 54:49]
  wire  IST1_reset; // @[Triangle.scala 54:49]
  wire  IST1_io_enable_IST1; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_nodeid_leaf_1; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_rayid_leaf_1; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_hiT_in; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_Oz; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_invDz; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_v11_in_x; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_v11_in_y; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_v11_in_z; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_v11_in_w; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_v22_in_x; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_v22_in_y; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_v22_in_z; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_v22_in_w; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_ray_o_in_x; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_ray_o_in_y; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_ray_o_in_z; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_ray_d_in_x; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_ray_d_in_y; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_ray_d_in_z; // @[Triangle.scala 54:49]
  wire  IST1_io_break_in; // @[Triangle.scala 54:49]
  wire  IST1_io_RAY_AABB_1; // @[Triangle.scala 54:49]
  wire  IST1_io_RAY_AABB_2; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_nodeid_ist1_out; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_rayid_ist1_out; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_hiT_out; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_t; // @[Triangle.scala 54:49]
  wire  IST1_io_pop_1; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_v11_out_x; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_v11_out_y; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_v11_out_z; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_v11_out_w; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_v22_out_x; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_v22_out_y; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_v22_out_z; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_v22_out_w; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_ray_o_out_x; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_ray_o_out_y; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_ray_o_out_z; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_ray_d_out_x; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_ray_d_out_y; // @[Triangle.scala 54:49]
  wire [31:0] IST1_io_ray_d_out_z; // @[Triangle.scala 54:49]
  wire  IST1_io_enable_IST2; // @[Triangle.scala 54:49]
  wire  IST1_io_break_out; // @[Triangle.scala 54:49]
  wire  IST1_io_break_ist1; // @[Triangle.scala 54:49]
  wire  IST1_io_RAY_AABB_1_out; // @[Triangle.scala 54:49]
  wire  IST1_io_RAY_AABB_2_out; // @[Triangle.scala 54:49]
  wire  IST2_clock; // @[Triangle.scala 55:49]
  wire  IST2_reset; // @[Triangle.scala 55:49]
  wire  IST2_io_enable_IST2; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_nodeid_leaf_2; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_rayid_leaf_2; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_hiT_in; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_v11_in_x; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_v11_in_y; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_v11_in_z; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_v11_in_w; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_v22_in_x; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_v22_in_y; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_v22_in_z; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_v22_in_w; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_ray_o_in_x; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_ray_o_in_y; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_ray_o_in_z; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_ray_d_in_x; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_ray_d_in_y; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_ray_d_in_z; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_t; // @[Triangle.scala 55:49]
  wire  IST2_io_break_in; // @[Triangle.scala 55:49]
  wire  IST2_io_RAY_AABB_1; // @[Triangle.scala 55:49]
  wire  IST2_io_RAY_AABB_2; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_nodeid_ist2_out; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_rayid_ist2_out; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_hiT_out; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_u; // @[Triangle.scala 55:49]
  wire  IST2_io_pop_2; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_t_out; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_v22_out_x; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_v22_out_y; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_v22_out_z; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_v22_out_w; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_ray_o_out_x; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_ray_o_out_y; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_ray_o_out_z; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_ray_d_out_x; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_ray_d_out_y; // @[Triangle.scala 55:49]
  wire [31:0] IST2_io_ray_d_out_z; // @[Triangle.scala 55:49]
  wire  IST2_io_enable_IST3; // @[Triangle.scala 55:49]
  wire  IST2_io_break_ist2; // @[Triangle.scala 55:49]
  wire  IST2_io_break_out; // @[Triangle.scala 55:49]
  wire  IST2_io_RAY_AABB_1_out; // @[Triangle.scala 55:49]
  wire  IST2_io_RAY_AABB_2_out; // @[Triangle.scala 55:49]
  wire  IST3_clock; // @[Triangle.scala 56:49]
  wire  IST3_reset; // @[Triangle.scala 56:49]
  wire  IST3_io_enable_IST3; // @[Triangle.scala 56:49]
  wire [31:0] IST3_io_nodeid_leaf_3; // @[Triangle.scala 56:49]
  wire [31:0] IST3_io_rayid_leaf_3; // @[Triangle.scala 56:49]
  wire [31:0] IST3_io_hiT_in; // @[Triangle.scala 56:49]
  wire [31:0] IST3_io_t_in; // @[Triangle.scala 56:49]
  wire [31:0] IST3_io_v22_in_x; // @[Triangle.scala 56:49]
  wire [31:0] IST3_io_v22_in_y; // @[Triangle.scala 56:49]
  wire [31:0] IST3_io_v22_in_z; // @[Triangle.scala 56:49]
  wire [31:0] IST3_io_v22_in_w; // @[Triangle.scala 56:49]
  wire [31:0] IST3_io_ray_o_in_x; // @[Triangle.scala 56:49]
  wire [31:0] IST3_io_ray_o_in_y; // @[Triangle.scala 56:49]
  wire [31:0] IST3_io_ray_o_in_z; // @[Triangle.scala 56:49]
  wire [31:0] IST3_io_ray_d_in_x; // @[Triangle.scala 56:49]
  wire [31:0] IST3_io_ray_d_in_y; // @[Triangle.scala 56:49]
  wire [31:0] IST3_io_ray_d_in_z; // @[Triangle.scala 56:49]
  wire [31:0] IST3_io_u_in; // @[Triangle.scala 56:49]
  wire  IST3_io_break_in; // @[Triangle.scala 56:49]
  wire  IST3_io_RAY_AABB_1; // @[Triangle.scala 56:49]
  wire  IST3_io_RAY_AABB_2; // @[Triangle.scala 56:49]
  wire [31:0] IST3_io_nodeid_ist3_out; // @[Triangle.scala 56:49]
  wire [31:0] IST3_io_rayid_ist3_out; // @[Triangle.scala 56:49]
  wire [31:0] IST3_io_hiT_out; // @[Triangle.scala 56:49]
  wire  IST3_io_hitT_en; // @[Triangle.scala 56:49]
  wire  IST3_io_pop_3; // @[Triangle.scala 56:49]
  wire [31:0] IST3_io_hitIndex; // @[Triangle.scala 56:49]
  wire  IST3_io_break_out; // @[Triangle.scala 56:49]
  wire  IST3_io_RAY_AABB_1_out; // @[Triangle.scala 56:49]
  wire  IST3_io_RAY_AABB_2_out; // @[Triangle.scala 56:49]
  IST0 IST0 ( // @[Triangle.scala 52:49]
    .clock(IST0_clock),
    .reset(IST0_reset),
    .io_enable_IST0(IST0_io_enable_IST0),
    .io_nodeid_leaf(IST0_io_nodeid_leaf),
    .io_rayid_leaf(IST0_io_rayid_leaf),
    .io_hiT_in(IST0_io_hiT_in),
    .io_v00_x(IST0_io_v00_x),
    .io_v00_y(IST0_io_v00_y),
    .io_v00_z(IST0_io_v00_z),
    .io_v00_w(IST0_io_v00_w),
    .io_v11_in_x(IST0_io_v11_in_x),
    .io_v11_in_y(IST0_io_v11_in_y),
    .io_v11_in_z(IST0_io_v11_in_z),
    .io_v11_in_w(IST0_io_v11_in_w),
    .io_v22_in_x(IST0_io_v22_in_x),
    .io_v22_in_y(IST0_io_v22_in_y),
    .io_v22_in_z(IST0_io_v22_in_z),
    .io_v22_in_w(IST0_io_v22_in_w),
    .io_ray_o_in_x(IST0_io_ray_o_in_x),
    .io_ray_o_in_y(IST0_io_ray_o_in_y),
    .io_ray_o_in_z(IST0_io_ray_o_in_z),
    .io_ray_d_in_x(IST0_io_ray_d_in_x),
    .io_ray_d_in_y(IST0_io_ray_d_in_y),
    .io_ray_d_in_z(IST0_io_ray_d_in_z),
    .io_RAY_AABB_1(IST0_io_RAY_AABB_1),
    .io_RAY_AABB_2(IST0_io_RAY_AABB_2),
    .io_break_in(IST0_io_break_in),
    .io_Oz(IST0_io_Oz),
    .io_invDz_div(IST0_io_invDz_div),
    .io_nodeid_ist0_out(IST0_io_nodeid_ist0_out),
    .io_rayid_ist0_out(IST0_io_rayid_ist0_out),
    .io_hiT_out(IST0_io_hiT_out),
    .io_v11_out_x(IST0_io_v11_out_x),
    .io_v11_out_y(IST0_io_v11_out_y),
    .io_v11_out_z(IST0_io_v11_out_z),
    .io_v11_out_w(IST0_io_v11_out_w),
    .io_v22_out_x(IST0_io_v22_out_x),
    .io_v22_out_y(IST0_io_v22_out_y),
    .io_v22_out_z(IST0_io_v22_out_z),
    .io_v22_out_w(IST0_io_v22_out_w),
    .io_ray_o_out_x(IST0_io_ray_o_out_x),
    .io_ray_o_out_y(IST0_io_ray_o_out_y),
    .io_ray_o_out_z(IST0_io_ray_o_out_z),
    .io_ray_d_out_x(IST0_io_ray_d_out_x),
    .io_ray_d_out_y(IST0_io_ray_d_out_y),
    .io_ray_d_out_z(IST0_io_ray_d_out_z),
    .io_enable_SU_out(IST0_io_enable_SU_out),
    .io_break_out(IST0_io_break_out),
    .io_RAY_AABB_1_out(IST0_io_RAY_AABB_1_out),
    .io_RAY_AABB_2_out(IST0_io_RAY_AABB_2_out)
  );
  Schedule_unit SU ( // @[Triangle.scala 53:50]
    .clock(SU_clock),
    .reset(SU_reset),
    .io_invDz_div(SU_io_invDz_div),
    .io_valid_in(SU_io_valid_in),
    .io_v11_x(SU_io_v11_x),
    .io_v11_y(SU_io_v11_y),
    .io_v11_z(SU_io_v11_z),
    .io_v11_w(SU_io_v11_w),
    .io_v22_x(SU_io_v22_x),
    .io_v22_y(SU_io_v22_y),
    .io_v22_z(SU_io_v22_z),
    .io_v22_w(SU_io_v22_w),
    .io_ray_in(SU_io_ray_in),
    .io_Oz(SU_io_Oz),
    .io_ray_o_in_x(SU_io_ray_o_in_x),
    .io_ray_o_in_y(SU_io_ray_o_in_y),
    .io_ray_o_in_z(SU_io_ray_o_in_z),
    .io_ray_d_in_x(SU_io_ray_d_in_x),
    .io_ray_d_in_y(SU_io_ray_d_in_y),
    .io_ray_d_in_z(SU_io_ray_d_in_z),
    .io_node_id_in(SU_io_node_id_in),
    .io_hitT_in(SU_io_hitT_in),
    .io_break_in(SU_io_break_in),
    .io_RAY_AABB_1(SU_io_RAY_AABB_1),
    .io_RAY_AABB_2(SU_io_RAY_AABB_2),
    .io_fdiv_out(SU_io_fdiv_out),
    .io_valid_out(SU_io_valid_out),
    .io_v11_out_x(SU_io_v11_out_x),
    .io_v11_out_y(SU_io_v11_out_y),
    .io_v11_out_z(SU_io_v11_out_z),
    .io_v11_out_w(SU_io_v11_out_w),
    .io_v22_out_x(SU_io_v22_out_x),
    .io_v22_out_y(SU_io_v22_out_y),
    .io_v22_out_z(SU_io_v22_out_z),
    .io_v22_out_w(SU_io_v22_out_w),
    .io_ray_out(SU_io_ray_out),
    .io_Oz_out(SU_io_Oz_out),
    .io_ray_o_out_x(SU_io_ray_o_out_x),
    .io_ray_o_out_y(SU_io_ray_o_out_y),
    .io_ray_o_out_z(SU_io_ray_o_out_z),
    .io_ray_d_out_x(SU_io_ray_d_out_x),
    .io_ray_d_out_y(SU_io_ray_d_out_y),
    .io_ray_d_out_z(SU_io_ray_d_out_z),
    .io_node_id_out(SU_io_node_id_out),
    .io_hitT_out(SU_io_hitT_out),
    .io_counter_fdiv(SU_io_counter_fdiv),
    .io_break_out(SU_io_break_out),
    .io_RAY_AABB_1_out(SU_io_RAY_AABB_1_out),
    .io_RAY_AABB_2_out(SU_io_RAY_AABB_2_out)
  );
  IST1 IST1 ( // @[Triangle.scala 54:49]
    .clock(IST1_clock),
    .reset(IST1_reset),
    .io_enable_IST1(IST1_io_enable_IST1),
    .io_nodeid_leaf_1(IST1_io_nodeid_leaf_1),
    .io_rayid_leaf_1(IST1_io_rayid_leaf_1),
    .io_hiT_in(IST1_io_hiT_in),
    .io_Oz(IST1_io_Oz),
    .io_invDz(IST1_io_invDz),
    .io_v11_in_x(IST1_io_v11_in_x),
    .io_v11_in_y(IST1_io_v11_in_y),
    .io_v11_in_z(IST1_io_v11_in_z),
    .io_v11_in_w(IST1_io_v11_in_w),
    .io_v22_in_x(IST1_io_v22_in_x),
    .io_v22_in_y(IST1_io_v22_in_y),
    .io_v22_in_z(IST1_io_v22_in_z),
    .io_v22_in_w(IST1_io_v22_in_w),
    .io_ray_o_in_x(IST1_io_ray_o_in_x),
    .io_ray_o_in_y(IST1_io_ray_o_in_y),
    .io_ray_o_in_z(IST1_io_ray_o_in_z),
    .io_ray_d_in_x(IST1_io_ray_d_in_x),
    .io_ray_d_in_y(IST1_io_ray_d_in_y),
    .io_ray_d_in_z(IST1_io_ray_d_in_z),
    .io_break_in(IST1_io_break_in),
    .io_RAY_AABB_1(IST1_io_RAY_AABB_1),
    .io_RAY_AABB_2(IST1_io_RAY_AABB_2),
    .io_nodeid_ist1_out(IST1_io_nodeid_ist1_out),
    .io_rayid_ist1_out(IST1_io_rayid_ist1_out),
    .io_hiT_out(IST1_io_hiT_out),
    .io_t(IST1_io_t),
    .io_pop_1(IST1_io_pop_1),
    .io_v11_out_x(IST1_io_v11_out_x),
    .io_v11_out_y(IST1_io_v11_out_y),
    .io_v11_out_z(IST1_io_v11_out_z),
    .io_v11_out_w(IST1_io_v11_out_w),
    .io_v22_out_x(IST1_io_v22_out_x),
    .io_v22_out_y(IST1_io_v22_out_y),
    .io_v22_out_z(IST1_io_v22_out_z),
    .io_v22_out_w(IST1_io_v22_out_w),
    .io_ray_o_out_x(IST1_io_ray_o_out_x),
    .io_ray_o_out_y(IST1_io_ray_o_out_y),
    .io_ray_o_out_z(IST1_io_ray_o_out_z),
    .io_ray_d_out_x(IST1_io_ray_d_out_x),
    .io_ray_d_out_y(IST1_io_ray_d_out_y),
    .io_ray_d_out_z(IST1_io_ray_d_out_z),
    .io_enable_IST2(IST1_io_enable_IST2),
    .io_break_out(IST1_io_break_out),
    .io_break_ist1(IST1_io_break_ist1),
    .io_RAY_AABB_1_out(IST1_io_RAY_AABB_1_out),
    .io_RAY_AABB_2_out(IST1_io_RAY_AABB_2_out)
  );
  IST2 IST2 ( // @[Triangle.scala 55:49]
    .clock(IST2_clock),
    .reset(IST2_reset),
    .io_enable_IST2(IST2_io_enable_IST2),
    .io_nodeid_leaf_2(IST2_io_nodeid_leaf_2),
    .io_rayid_leaf_2(IST2_io_rayid_leaf_2),
    .io_hiT_in(IST2_io_hiT_in),
    .io_v11_in_x(IST2_io_v11_in_x),
    .io_v11_in_y(IST2_io_v11_in_y),
    .io_v11_in_z(IST2_io_v11_in_z),
    .io_v11_in_w(IST2_io_v11_in_w),
    .io_v22_in_x(IST2_io_v22_in_x),
    .io_v22_in_y(IST2_io_v22_in_y),
    .io_v22_in_z(IST2_io_v22_in_z),
    .io_v22_in_w(IST2_io_v22_in_w),
    .io_ray_o_in_x(IST2_io_ray_o_in_x),
    .io_ray_o_in_y(IST2_io_ray_o_in_y),
    .io_ray_o_in_z(IST2_io_ray_o_in_z),
    .io_ray_d_in_x(IST2_io_ray_d_in_x),
    .io_ray_d_in_y(IST2_io_ray_d_in_y),
    .io_ray_d_in_z(IST2_io_ray_d_in_z),
    .io_t(IST2_io_t),
    .io_break_in(IST2_io_break_in),
    .io_RAY_AABB_1(IST2_io_RAY_AABB_1),
    .io_RAY_AABB_2(IST2_io_RAY_AABB_2),
    .io_nodeid_ist2_out(IST2_io_nodeid_ist2_out),
    .io_rayid_ist2_out(IST2_io_rayid_ist2_out),
    .io_hiT_out(IST2_io_hiT_out),
    .io_u(IST2_io_u),
    .io_pop_2(IST2_io_pop_2),
    .io_t_out(IST2_io_t_out),
    .io_v22_out_x(IST2_io_v22_out_x),
    .io_v22_out_y(IST2_io_v22_out_y),
    .io_v22_out_z(IST2_io_v22_out_z),
    .io_v22_out_w(IST2_io_v22_out_w),
    .io_ray_o_out_x(IST2_io_ray_o_out_x),
    .io_ray_o_out_y(IST2_io_ray_o_out_y),
    .io_ray_o_out_z(IST2_io_ray_o_out_z),
    .io_ray_d_out_x(IST2_io_ray_d_out_x),
    .io_ray_d_out_y(IST2_io_ray_d_out_y),
    .io_ray_d_out_z(IST2_io_ray_d_out_z),
    .io_enable_IST3(IST2_io_enable_IST3),
    .io_break_ist2(IST2_io_break_ist2),
    .io_break_out(IST2_io_break_out),
    .io_RAY_AABB_1_out(IST2_io_RAY_AABB_1_out),
    .io_RAY_AABB_2_out(IST2_io_RAY_AABB_2_out)
  );
  IST3 IST3 ( // @[Triangle.scala 56:49]
    .clock(IST3_clock),
    .reset(IST3_reset),
    .io_enable_IST3(IST3_io_enable_IST3),
    .io_nodeid_leaf_3(IST3_io_nodeid_leaf_3),
    .io_rayid_leaf_3(IST3_io_rayid_leaf_3),
    .io_hiT_in(IST3_io_hiT_in),
    .io_t_in(IST3_io_t_in),
    .io_v22_in_x(IST3_io_v22_in_x),
    .io_v22_in_y(IST3_io_v22_in_y),
    .io_v22_in_z(IST3_io_v22_in_z),
    .io_v22_in_w(IST3_io_v22_in_w),
    .io_ray_o_in_x(IST3_io_ray_o_in_x),
    .io_ray_o_in_y(IST3_io_ray_o_in_y),
    .io_ray_o_in_z(IST3_io_ray_o_in_z),
    .io_ray_d_in_x(IST3_io_ray_d_in_x),
    .io_ray_d_in_y(IST3_io_ray_d_in_y),
    .io_ray_d_in_z(IST3_io_ray_d_in_z),
    .io_u_in(IST3_io_u_in),
    .io_break_in(IST3_io_break_in),
    .io_RAY_AABB_1(IST3_io_RAY_AABB_1),
    .io_RAY_AABB_2(IST3_io_RAY_AABB_2),
    .io_nodeid_ist3_out(IST3_io_nodeid_ist3_out),
    .io_rayid_ist3_out(IST3_io_rayid_ist3_out),
    .io_hiT_out(IST3_io_hiT_out),
    .io_hitT_en(IST3_io_hitT_en),
    .io_pop_3(IST3_io_pop_3),
    .io_hitIndex(IST3_io_hitIndex),
    .io_break_out(IST3_io_break_out),
    .io_RAY_AABB_1_out(IST3_io_RAY_AABB_1_out),
    .io_RAY_AABB_2_out(IST3_io_RAY_AABB_2_out)
  );
  assign io_pop_1 = IST1_io_pop_1; // @[Triangle.scala 129:41]
  assign io_break_1 = IST1_io_break_out; // @[Triangle.scala 132:39]
  assign io_pop_2 = IST2_io_pop_2; // @[Triangle.scala 133:41]
  assign io_break_2 = IST2_io_break_out; // @[Triangle.scala 136:39]
  assign io_pop_3 = IST3_io_pop_3; // @[Triangle.scala 137:41]
  assign io_break_3 = IST3_io_break_out; // @[Triangle.scala 140:39]
  assign io_hiT_out_1 = IST1_io_hiT_out; // @[Triangle.scala 141:37]
  assign io_hiT_out_2 = IST2_io_hiT_out; // @[Triangle.scala 142:37]
  assign io_hiT_out_3 = IST3_io_hiT_out; // @[Triangle.scala 143:37]
  assign io_hitT_en = IST3_io_hitT_en; // @[Triangle.scala 144:40]
  assign io_hitIndex = IST3_io_hitIndex; // @[Triangle.scala 146:40]
  assign io_node_id_out_1 = IST1_io_nodeid_ist1_out; // @[Triangle.scala 131:30]
  assign io_node_id_out_2 = IST2_io_nodeid_ist2_out; // @[Triangle.scala 135:30]
  assign io_node_id_out_3 = IST3_io_nodeid_ist3_out; // @[Triangle.scala 139:30]
  assign io_ray_id_ist1 = IST1_io_rayid_ist1_out; // @[Triangle.scala 130:37]
  assign io_ray_id_ist2 = IST2_io_rayid_ist2_out; // @[Triangle.scala 134:37]
  assign io_ray_id_ist3 = IST3_io_rayid_ist3_out; // @[Triangle.scala 138:37]
  assign io_counter_fdiv = {{32'd0}, SU_io_counter_fdiv}; // @[Triangle.scala 85:37]
  assign io_RAY_AABB_1_out_IST1 = IST1_io_RAY_AABB_1_out; // @[Triangle.scala 148:33]
  assign io_RAY_AABB_2_out_IST1 = IST1_io_RAY_AABB_2_out; // @[Triangle.scala 149:33]
  assign io_RAY_AABB_1_out_IST2 = IST2_io_RAY_AABB_1_out; // @[Triangle.scala 150:33]
  assign io_RAY_AABB_2_out_IST2 = IST2_io_RAY_AABB_2_out; // @[Triangle.scala 151:33]
  assign io_RAY_AABB_1_out_IST3 = IST3_io_RAY_AABB_1_out; // @[Triangle.scala 152:33]
  assign io_RAY_AABB_2_out_IST3 = IST3_io_RAY_AABB_2_out; // @[Triangle.scala 153:33]
  assign IST0_clock = clock;
  assign IST0_reset = reset;
  assign IST0_io_enable_IST0 = io_To_IST0_enable; // @[Triangle.scala 61:32]
  assign IST0_io_nodeid_leaf = io_nodeid_leaf; // @[Triangle.scala 62:33]
  assign IST0_io_rayid_leaf = io_rayid_leaf; // @[Triangle.scala 63:36]
  assign IST0_io_hiT_in = io_hiT_in; // @[Triangle.scala 64:40]
  assign IST0_io_v00_x = io_v00_in_x; // @[Triangle.scala 65:43]
  assign IST0_io_v00_y = io_v00_in_y; // @[Triangle.scala 65:43]
  assign IST0_io_v00_z = io_v00_in_z; // @[Triangle.scala 65:43]
  assign IST0_io_v00_w = io_v00_in_w; // @[Triangle.scala 65:43]
  assign IST0_io_v11_in_x = io_v11_in_x; // @[Triangle.scala 66:40]
  assign IST0_io_v11_in_y = io_v11_in_y; // @[Triangle.scala 66:40]
  assign IST0_io_v11_in_z = io_v11_in_z; // @[Triangle.scala 66:40]
  assign IST0_io_v11_in_w = io_v11_in_w; // @[Triangle.scala 66:40]
  assign IST0_io_v22_in_x = io_v22_in_x; // @[Triangle.scala 67:40]
  assign IST0_io_v22_in_y = io_v22_in_y; // @[Triangle.scala 67:40]
  assign IST0_io_v22_in_z = io_v22_in_z; // @[Triangle.scala 67:40]
  assign IST0_io_v22_in_w = io_v22_in_w; // @[Triangle.scala 67:40]
  assign IST0_io_ray_o_in_x = io_ray_o_in_x; // @[Triangle.scala 68:37]
  assign IST0_io_ray_o_in_y = io_ray_o_in_y; // @[Triangle.scala 68:37]
  assign IST0_io_ray_o_in_z = io_ray_o_in_z; // @[Triangle.scala 68:37]
  assign IST0_io_ray_d_in_x = io_ray_d_in_x; // @[Triangle.scala 69:37]
  assign IST0_io_ray_d_in_y = io_ray_d_in_y; // @[Triangle.scala 69:37]
  assign IST0_io_ray_d_in_z = io_ray_d_in_z; // @[Triangle.scala 69:37]
  assign IST0_io_RAY_AABB_1 = io_RAY_AABB_1; // @[Triangle.scala 59:31]
  assign IST0_io_RAY_AABB_2 = io_RAY_AABB_2; // @[Triangle.scala 60:31]
  assign IST0_io_break_in = io_break_in; // @[Triangle.scala 70:37]
  assign SU_clock = clock;
  assign SU_reset = reset;
  assign SU_io_invDz_div = IST0_io_invDz_div; // @[Triangle.scala 77:36]
  assign SU_io_valid_in = IST0_io_enable_SU_out; // @[Triangle.scala 75:39]
  assign SU_io_v11_x = IST0_io_v11_out_x; // @[Triangle.scala 81:43]
  assign SU_io_v11_y = IST0_io_v11_out_y; // @[Triangle.scala 81:43]
  assign SU_io_v11_z = IST0_io_v11_out_z; // @[Triangle.scala 81:43]
  assign SU_io_v11_w = IST0_io_v11_out_w; // @[Triangle.scala 81:43]
  assign SU_io_v22_x = IST0_io_v22_out_x; // @[Triangle.scala 82:43]
  assign SU_io_v22_y = IST0_io_v22_out_y; // @[Triangle.scala 82:43]
  assign SU_io_v22_z = IST0_io_v22_out_z; // @[Triangle.scala 82:43]
  assign SU_io_v22_w = IST0_io_v22_out_w; // @[Triangle.scala 82:43]
  assign SU_io_ray_in = IST0_io_rayid_ist0_out; // @[Triangle.scala 79:40]
  assign SU_io_Oz = IST0_io_Oz; // @[Triangle.scala 76:44]
  assign SU_io_ray_o_in_x = IST0_io_ray_o_out_x; // @[Triangle.scala 83:37]
  assign SU_io_ray_o_in_y = IST0_io_ray_o_out_y; // @[Triangle.scala 83:37]
  assign SU_io_ray_o_in_z = IST0_io_ray_o_out_z; // @[Triangle.scala 83:37]
  assign SU_io_ray_d_in_x = IST0_io_ray_d_out_x; // @[Triangle.scala 84:37]
  assign SU_io_ray_d_in_y = IST0_io_ray_d_out_y; // @[Triangle.scala 84:37]
  assign SU_io_ray_d_in_z = IST0_io_ray_d_out_z; // @[Triangle.scala 84:37]
  assign SU_io_node_id_in = IST0_io_nodeid_ist0_out; // @[Triangle.scala 78:33]
  assign SU_io_hitT_in = IST0_io_hiT_out; // @[Triangle.scala 80:39]
  assign SU_io_break_in = IST0_io_break_out; // @[Triangle.scala 74:37]
  assign SU_io_RAY_AABB_1 = IST0_io_RAY_AABB_1_out; // @[Triangle.scala 72:31]
  assign SU_io_RAY_AABB_2 = IST0_io_RAY_AABB_2_out; // @[Triangle.scala 73:31]
  assign IST1_clock = clock;
  assign IST1_reset = reset;
  assign IST1_io_enable_IST1 = SU_io_valid_out; // @[Triangle.scala 90:32]
  assign IST1_io_nodeid_leaf_1 = SU_io_node_id_out; // @[Triangle.scala 91:30]
  assign IST1_io_rayid_leaf_1 = SU_io_ray_out; // @[Triangle.scala 92:33]
  assign IST1_io_hiT_in = SU_io_hitT_out; // @[Triangle.scala 93:40]
  assign IST1_io_Oz = SU_io_Oz_out; // @[Triangle.scala 94:44]
  assign IST1_io_invDz = SU_io_fdiv_out; // @[Triangle.scala 95:41]
  assign IST1_io_v11_in_x = SU_io_v11_out_x; // @[Triangle.scala 96:40]
  assign IST1_io_v11_in_y = SU_io_v11_out_y; // @[Triangle.scala 96:40]
  assign IST1_io_v11_in_z = SU_io_v11_out_z; // @[Triangle.scala 96:40]
  assign IST1_io_v11_in_w = SU_io_v11_out_w; // @[Triangle.scala 96:40]
  assign IST1_io_v22_in_x = SU_io_v22_out_x; // @[Triangle.scala 97:40]
  assign IST1_io_v22_in_y = SU_io_v22_out_y; // @[Triangle.scala 97:40]
  assign IST1_io_v22_in_z = SU_io_v22_out_z; // @[Triangle.scala 97:40]
  assign IST1_io_v22_in_w = SU_io_v22_out_w; // @[Triangle.scala 97:40]
  assign IST1_io_ray_o_in_x = SU_io_ray_o_out_x; // @[Triangle.scala 98:37]
  assign IST1_io_ray_o_in_y = SU_io_ray_o_out_y; // @[Triangle.scala 98:37]
  assign IST1_io_ray_o_in_z = SU_io_ray_o_out_z; // @[Triangle.scala 98:37]
  assign IST1_io_ray_d_in_x = SU_io_ray_d_out_x; // @[Triangle.scala 99:37]
  assign IST1_io_ray_d_in_y = SU_io_ray_d_out_y; // @[Triangle.scala 99:37]
  assign IST1_io_ray_d_in_z = SU_io_ray_d_out_z; // @[Triangle.scala 99:37]
  assign IST1_io_break_in = SU_io_break_out; // @[Triangle.scala 89:36]
  assign IST1_io_RAY_AABB_1 = SU_io_RAY_AABB_1_out; // @[Triangle.scala 87:30]
  assign IST1_io_RAY_AABB_2 = SU_io_RAY_AABB_2_out; // @[Triangle.scala 88:30]
  assign IST2_clock = clock;
  assign IST2_reset = reset;
  assign IST2_io_enable_IST2 = IST1_io_enable_IST2; // @[Triangle.scala 105:35]
  assign IST2_io_nodeid_leaf_2 = IST1_io_nodeid_ist1_out; // @[Triangle.scala 106:33]
  assign IST2_io_rayid_leaf_2 = IST1_io_rayid_ist1_out; // @[Triangle.scala 107:36]
  assign IST2_io_hiT_in = IST1_io_hiT_out; // @[Triangle.scala 108:42]
  assign IST2_io_v11_in_x = IST1_io_v11_out_x; // @[Triangle.scala 109:42]
  assign IST2_io_v11_in_y = IST1_io_v11_out_y; // @[Triangle.scala 109:42]
  assign IST2_io_v11_in_z = IST1_io_v11_out_z; // @[Triangle.scala 109:42]
  assign IST2_io_v11_in_w = IST1_io_v11_out_w; // @[Triangle.scala 109:42]
  assign IST2_io_v22_in_x = IST1_io_v22_out_x; // @[Triangle.scala 110:42]
  assign IST2_io_v22_in_y = IST1_io_v22_out_y; // @[Triangle.scala 110:42]
  assign IST2_io_v22_in_z = IST1_io_v22_out_z; // @[Triangle.scala 110:42]
  assign IST2_io_v22_in_w = IST1_io_v22_out_w; // @[Triangle.scala 110:42]
  assign IST2_io_ray_o_in_x = IST1_io_ray_o_out_x; // @[Triangle.scala 111:40]
  assign IST2_io_ray_o_in_y = IST1_io_ray_o_out_y; // @[Triangle.scala 111:40]
  assign IST2_io_ray_o_in_z = IST1_io_ray_o_out_z; // @[Triangle.scala 111:40]
  assign IST2_io_ray_d_in_x = IST1_io_ray_d_out_x; // @[Triangle.scala 112:40]
  assign IST2_io_ray_d_in_y = IST1_io_ray_d_out_y; // @[Triangle.scala 112:40]
  assign IST2_io_ray_d_in_z = IST1_io_ray_d_out_z; // @[Triangle.scala 112:40]
  assign IST2_io_t = IST1_io_t; // @[Triangle.scala 113:49]
  assign IST2_io_break_in = IST1_io_break_ist1; // @[Triangle.scala 103:39]
  assign IST2_io_RAY_AABB_1 = IST1_io_RAY_AABB_1_out; // @[Triangle.scala 101:33]
  assign IST2_io_RAY_AABB_2 = IST1_io_RAY_AABB_2_out; // @[Triangle.scala 102:33]
  assign IST3_clock = clock;
  assign IST3_reset = reset;
  assign IST3_io_enable_IST3 = IST2_io_enable_IST3; // @[Triangle.scala 118:38]
  assign IST3_io_nodeid_leaf_3 = IST2_io_nodeid_ist2_out; // @[Triangle.scala 119:36]
  assign IST3_io_rayid_leaf_3 = IST2_io_rayid_ist2_out; // @[Triangle.scala 120:39]
  assign IST3_io_hiT_in = IST2_io_hiT_out; // @[Triangle.scala 121:45]
  assign IST3_io_t_in = IST2_io_t_out; // @[Triangle.scala 122:48]
  assign IST3_io_v22_in_x = IST2_io_v22_out_x; // @[Triangle.scala 123:45]
  assign IST3_io_v22_in_y = IST2_io_v22_out_y; // @[Triangle.scala 123:45]
  assign IST3_io_v22_in_z = IST2_io_v22_out_z; // @[Triangle.scala 123:45]
  assign IST3_io_v22_in_w = IST2_io_v22_out_w; // @[Triangle.scala 123:45]
  assign IST3_io_ray_o_in_x = IST2_io_ray_o_out_x; // @[Triangle.scala 124:41]
  assign IST3_io_ray_o_in_y = IST2_io_ray_o_out_y; // @[Triangle.scala 124:41]
  assign IST3_io_ray_o_in_z = IST2_io_ray_o_out_z; // @[Triangle.scala 124:41]
  assign IST3_io_ray_d_in_x = IST2_io_ray_d_out_x; // @[Triangle.scala 125:41]
  assign IST3_io_ray_d_in_y = IST2_io_ray_d_out_y; // @[Triangle.scala 125:41]
  assign IST3_io_ray_d_in_z = IST2_io_ray_d_out_z; // @[Triangle.scala 125:41]
  assign IST3_io_u_in = IST2_io_u; // @[Triangle.scala 126:47]
  assign IST3_io_break_in = IST2_io_break_ist2; // @[Triangle.scala 117:42]
  assign IST3_io_RAY_AABB_1 = IST2_io_RAY_AABB_1_out; // @[Triangle.scala 115:35]
  assign IST3_io_RAY_AABB_2 = IST2_io_RAY_AABB_2_out; // @[Triangle.scala 116:35]
endmodule
module TOP_1(
  input         clock,
  input         reset,
  output [31:0] io_hitT,
  output [31:0] io_hitIndex,
  output        io_rtp_finish,
  output [31:0] io_ray_id_triangle,
  output [63:0] io_counter_fdiv,
  output [63:0] io_TRV_1_valid,
  output [63:0] io_TRV_2_valid,
  output [63:0] io_IST_1_valid,
  output [63:0] io_clock_count
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [63:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  wire  Ray_Dispatch_clock; // @[Top_1.scala 24:44]
  wire  Ray_Dispatch_reset; // @[Top_1.scala 24:44]
  wire  Ray_Dispatch_io_dispatch; // @[Top_1.scala 24:44]
  wire  Ray_Dispatch_io_dispatch_2; // @[Top_1.scala 24:44]
  wire [31:0] Ray_Dispatch_io_rayid_id; // @[Top_1.scala 24:44]
  wire [31:0] Ray_Dispatch_io_rayid_id_2; // @[Top_1.scala 24:44]
  wire  Ray_Dispatch_io_ray_out; // @[Top_1.scala 24:44]
  wire  Ray_Dispatch_io_ray_out_2; // @[Top_1.scala 24:44]
  wire  Ray_Dispatch_io_ray_finish; // @[Top_1.scala 24:44]
  wire  Ray_origx_clock; // @[Top_1.scala 25:48]
  wire [31:0] Ray_origx_io_Ray_id; // @[Top_1.scala 25:48]
  wire [31:0] Ray_origx_io_Ray_id_2; // @[Top_1.scala 25:48]
  wire [31:0] Ray_origx_io_Ray_out; // @[Top_1.scala 25:48]
  wire [31:0] Ray_origx_io_Ray_out_2; // @[Top_1.scala 25:48]
  wire  Ray_origy_clock; // @[Top_1.scala 26:48]
  wire [31:0] Ray_origy_io_Ray_id; // @[Top_1.scala 26:48]
  wire [31:0] Ray_origy_io_Ray_id_2; // @[Top_1.scala 26:48]
  wire [31:0] Ray_origy_io_Ray_out; // @[Top_1.scala 26:48]
  wire [31:0] Ray_origy_io_Ray_out_2; // @[Top_1.scala 26:48]
  wire  Ray_origz_clock; // @[Top_1.scala 27:48]
  wire [31:0] Ray_origz_io_Ray_id; // @[Top_1.scala 27:48]
  wire [31:0] Ray_origz_io_Ray_id_2; // @[Top_1.scala 27:48]
  wire [31:0] Ray_origz_io_Ray_out; // @[Top_1.scala 27:48]
  wire [31:0] Ray_origz_io_Ray_out_2; // @[Top_1.scala 27:48]
  wire  Ray_dirx_clock; // @[Top_1.scala 30:50]
  wire [31:0] Ray_dirx_io_Ray_id; // @[Top_1.scala 30:50]
  wire [31:0] Ray_dirx_io_Ray_id_2; // @[Top_1.scala 30:50]
  wire [31:0] Ray_dirx_io_Ray_out; // @[Top_1.scala 30:50]
  wire [31:0] Ray_dirx_io_Ray_out_2; // @[Top_1.scala 30:50]
  wire  Ray_diry_clock; // @[Top_1.scala 31:49]
  wire [31:0] Ray_diry_io_Ray_id; // @[Top_1.scala 31:49]
  wire [31:0] Ray_diry_io_Ray_id_2; // @[Top_1.scala 31:49]
  wire [31:0] Ray_diry_io_Ray_out; // @[Top_1.scala 31:49]
  wire [31:0] Ray_diry_io_Ray_out_2; // @[Top_1.scala 31:49]
  wire  Ray_dirz_clock; // @[Top_1.scala 32:49]
  wire [31:0] Ray_dirz_io_Ray_id; // @[Top_1.scala 32:49]
  wire [31:0] Ray_dirz_io_Ray_id_2; // @[Top_1.scala 32:49]
  wire [31:0] Ray_dirz_io_Ray_out; // @[Top_1.scala 32:49]
  wire [31:0] Ray_dirz_io_Ray_out_2; // @[Top_1.scala 32:49]
  wire  Ray_hitT_clock; // @[Top_1.scala 33:49]
  wire [31:0] Ray_hitT_io_Ray_id; // @[Top_1.scala 33:49]
  wire [31:0] Ray_hitT_io_Ray_id_2; // @[Top_1.scala 33:49]
  wire [31:0] Ray_hitT_io_Ray_out; // @[Top_1.scala 33:49]
  wire [31:0] Ray_hitT_io_Ray_out_2; // @[Top_1.scala 33:49]
  wire  Ray_idirx_clock; // @[Top_1.scala 35:49]
  wire [31:0] Ray_idirx_io_Ray_id; // @[Top_1.scala 35:49]
  wire [31:0] Ray_idirx_io_Ray_id_2; // @[Top_1.scala 35:49]
  wire [31:0] Ray_idirx_io_Ray_out; // @[Top_1.scala 35:49]
  wire [31:0] Ray_idirx_io_Ray_out_2; // @[Top_1.scala 35:49]
  wire  Ray_idiry_clock; // @[Top_1.scala 36:49]
  wire [31:0] Ray_idiry_io_Ray_id; // @[Top_1.scala 36:49]
  wire [31:0] Ray_idiry_io_Ray_id_2; // @[Top_1.scala 36:49]
  wire [31:0] Ray_idiry_io_Ray_out; // @[Top_1.scala 36:49]
  wire [31:0] Ray_idiry_io_Ray_out_2; // @[Top_1.scala 36:49]
  wire  Ray_idirz_clock; // @[Top_1.scala 37:49]
  wire [31:0] Ray_idirz_io_Ray_id; // @[Top_1.scala 37:49]
  wire [31:0] Ray_idirz_io_Ray_id_2; // @[Top_1.scala 37:49]
  wire [31:0] Ray_idirz_io_Ray_out; // @[Top_1.scala 37:49]
  wire [31:0] Ray_idirz_io_Ray_out_2; // @[Top_1.scala 37:49]
  wire  Ray_oodx_clock; // @[Top_1.scala 39:48]
  wire [31:0] Ray_oodx_io_Ray_id; // @[Top_1.scala 39:48]
  wire [31:0] Ray_oodx_io_Ray_id_2; // @[Top_1.scala 39:48]
  wire [31:0] Ray_oodx_io_Ray_out; // @[Top_1.scala 39:48]
  wire [31:0] Ray_oodx_io_Ray_out_2; // @[Top_1.scala 39:48]
  wire  Ray_oody_clock; // @[Top_1.scala 40:48]
  wire [31:0] Ray_oody_io_Ray_id; // @[Top_1.scala 40:48]
  wire [31:0] Ray_oody_io_Ray_id_2; // @[Top_1.scala 40:48]
  wire [31:0] Ray_oody_io_Ray_out; // @[Top_1.scala 40:48]
  wire [31:0] Ray_oody_io_Ray_out_2; // @[Top_1.scala 40:48]
  wire  Ray_oodz_clock; // @[Top_1.scala 41:48]
  wire [31:0] Ray_oodz_io_Ray_id; // @[Top_1.scala 41:48]
  wire [31:0] Ray_oodz_io_Ray_id_2; // @[Top_1.scala 41:48]
  wire [31:0] Ray_oodz_io_Ray_out; // @[Top_1.scala 41:48]
  wire [31:0] Ray_oodz_io_Ray_out_2; // @[Top_1.scala 41:48]
  wire  BVH_RAM_0_x_clock; // @[Top_1.scala 43:41]
  wire [31:0] BVH_RAM_0_x_io_BVH_id; // @[Top_1.scala 43:41]
  wire [31:0] BVH_RAM_0_x_io_BVH_id_2; // @[Top_1.scala 43:41]
  wire [31:0] BVH_RAM_0_x_io_BVH_out; // @[Top_1.scala 43:41]
  wire [31:0] BVH_RAM_0_x_io_BVH_out_2; // @[Top_1.scala 43:41]
  wire  BVH_RAM_0_y_clock; // @[Top_1.scala 44:41]
  wire [31:0] BVH_RAM_0_y_io_BVH_id; // @[Top_1.scala 44:41]
  wire [31:0] BVH_RAM_0_y_io_BVH_id_2; // @[Top_1.scala 44:41]
  wire [31:0] BVH_RAM_0_y_io_BVH_out; // @[Top_1.scala 44:41]
  wire [31:0] BVH_RAM_0_y_io_BVH_out_2; // @[Top_1.scala 44:41]
  wire  BVH_RAM_0_z_clock; // @[Top_1.scala 45:41]
  wire [31:0] BVH_RAM_0_z_io_BVH_id; // @[Top_1.scala 45:41]
  wire [31:0] BVH_RAM_0_z_io_BVH_id_2; // @[Top_1.scala 45:41]
  wire [31:0] BVH_RAM_0_z_io_BVH_out; // @[Top_1.scala 45:41]
  wire [31:0] BVH_RAM_0_z_io_BVH_out_2; // @[Top_1.scala 45:41]
  wire  BVH_RAM_0_w_clock; // @[Top_1.scala 46:40]
  wire [31:0] BVH_RAM_0_w_io_BVH_id; // @[Top_1.scala 46:40]
  wire [31:0] BVH_RAM_0_w_io_BVH_id_2; // @[Top_1.scala 46:40]
  wire [31:0] BVH_RAM_0_w_io_BVH_out; // @[Top_1.scala 46:40]
  wire [31:0] BVH_RAM_0_w_io_BVH_out_2; // @[Top_1.scala 46:40]
  wire  BVH_RAM_1_x_clock; // @[Top_1.scala 48:41]
  wire [31:0] BVH_RAM_1_x_io_BVH_id; // @[Top_1.scala 48:41]
  wire [31:0] BVH_RAM_1_x_io_BVH_id_2; // @[Top_1.scala 48:41]
  wire [31:0] BVH_RAM_1_x_io_BVH_out; // @[Top_1.scala 48:41]
  wire [31:0] BVH_RAM_1_x_io_BVH_out_2; // @[Top_1.scala 48:41]
  wire  BVH_RAM_1_y_clock; // @[Top_1.scala 49:41]
  wire [31:0] BVH_RAM_1_y_io_BVH_id; // @[Top_1.scala 49:41]
  wire [31:0] BVH_RAM_1_y_io_BVH_id_2; // @[Top_1.scala 49:41]
  wire [31:0] BVH_RAM_1_y_io_BVH_out; // @[Top_1.scala 49:41]
  wire [31:0] BVH_RAM_1_y_io_BVH_out_2; // @[Top_1.scala 49:41]
  wire  BVH_RAM_1_z_clock; // @[Top_1.scala 50:41]
  wire [31:0] BVH_RAM_1_z_io_BVH_id; // @[Top_1.scala 50:41]
  wire [31:0] BVH_RAM_1_z_io_BVH_id_2; // @[Top_1.scala 50:41]
  wire [31:0] BVH_RAM_1_z_io_BVH_out; // @[Top_1.scala 50:41]
  wire [31:0] BVH_RAM_1_z_io_BVH_out_2; // @[Top_1.scala 50:41]
  wire  BVH_RAM_1_w_clock; // @[Top_1.scala 51:40]
  wire [31:0] BVH_RAM_1_w_io_BVH_id; // @[Top_1.scala 51:40]
  wire [31:0] BVH_RAM_1_w_io_BVH_id_2; // @[Top_1.scala 51:40]
  wire [31:0] BVH_RAM_1_w_io_BVH_out; // @[Top_1.scala 51:40]
  wire [31:0] BVH_RAM_1_w_io_BVH_out_2; // @[Top_1.scala 51:40]
  wire  BVH_RAM_z_x_clock; // @[Top_1.scala 53:41]
  wire [31:0] BVH_RAM_z_x_io_BVH_id; // @[Top_1.scala 53:41]
  wire [31:0] BVH_RAM_z_x_io_BVH_id_2; // @[Top_1.scala 53:41]
  wire [31:0] BVH_RAM_z_x_io_BVH_out; // @[Top_1.scala 53:41]
  wire [31:0] BVH_RAM_z_x_io_BVH_out_2; // @[Top_1.scala 53:41]
  wire  BVH_RAM_z_y_clock; // @[Top_1.scala 54:41]
  wire [31:0] BVH_RAM_z_y_io_BVH_id; // @[Top_1.scala 54:41]
  wire [31:0] BVH_RAM_z_y_io_BVH_id_2; // @[Top_1.scala 54:41]
  wire [31:0] BVH_RAM_z_y_io_BVH_out; // @[Top_1.scala 54:41]
  wire [31:0] BVH_RAM_z_y_io_BVH_out_2; // @[Top_1.scala 54:41]
  wire  BVH_RAM_z_z_clock; // @[Top_1.scala 55:41]
  wire [31:0] BVH_RAM_z_z_io_BVH_id; // @[Top_1.scala 55:41]
  wire [31:0] BVH_RAM_z_z_io_BVH_id_2; // @[Top_1.scala 55:41]
  wire [31:0] BVH_RAM_z_z_io_BVH_out; // @[Top_1.scala 55:41]
  wire [31:0] BVH_RAM_z_z_io_BVH_out_2; // @[Top_1.scala 55:41]
  wire  BVH_RAM_z_w_clock; // @[Top_1.scala 56:40]
  wire [31:0] BVH_RAM_z_w_io_BVH_id; // @[Top_1.scala 56:40]
  wire [31:0] BVH_RAM_z_w_io_BVH_id_2; // @[Top_1.scala 56:40]
  wire [31:0] BVH_RAM_z_w_io_BVH_out; // @[Top_1.scala 56:40]
  wire [31:0] BVH_RAM_z_w_io_BVH_out_2; // @[Top_1.scala 56:40]
  wire  BVH_RAM_tmp_x_clock; // @[Top_1.scala 58:37]
  wire [31:0] BVH_RAM_tmp_x_io_BVH_id; // @[Top_1.scala 58:37]
  wire [31:0] BVH_RAM_tmp_x_io_BVH_id_2; // @[Top_1.scala 58:37]
  wire [31:0] BVH_RAM_tmp_x_io_BVH_out; // @[Top_1.scala 58:37]
  wire [31:0] BVH_RAM_tmp_x_io_BVH_out_2; // @[Top_1.scala 58:37]
  wire  BVH_RAM_tmp_y_clock; // @[Top_1.scala 59:37]
  wire [31:0] BVH_RAM_tmp_y_io_BVH_id; // @[Top_1.scala 59:37]
  wire [31:0] BVH_RAM_tmp_y_io_BVH_id_2; // @[Top_1.scala 59:37]
  wire [31:0] BVH_RAM_tmp_y_io_BVH_out; // @[Top_1.scala 59:37]
  wire [31:0] BVH_RAM_tmp_y_io_BVH_out_2; // @[Top_1.scala 59:37]
  wire  TRI_RAM_x_clock; // @[Top_1.scala 61:50]
  wire [31:0] TRI_RAM_x_io_Triangle_id; // @[Top_1.scala 61:50]
  wire [31:0] TRI_RAM_x_io_v00_out; // @[Top_1.scala 61:50]
  wire [31:0] TRI_RAM_x_io_v11_out; // @[Top_1.scala 61:50]
  wire [31:0] TRI_RAM_x_io_v22_out; // @[Top_1.scala 61:50]
  wire [31:0] TRI_RAM_x_io_valid; // @[Top_1.scala 61:50]
  wire  TRI_RAM_y_clock; // @[Top_1.scala 62:50]
  wire [31:0] TRI_RAM_y_io_Triangle_id; // @[Top_1.scala 62:50]
  wire [31:0] TRI_RAM_y_io_v00_out; // @[Top_1.scala 62:50]
  wire [31:0] TRI_RAM_y_io_v11_out; // @[Top_1.scala 62:50]
  wire [31:0] TRI_RAM_y_io_v22_out; // @[Top_1.scala 62:50]
  wire  TRI_RAM_z_clock; // @[Top_1.scala 63:50]
  wire [31:0] TRI_RAM_z_io_Triangle_id; // @[Top_1.scala 63:50]
  wire [31:0] TRI_RAM_z_io_v00_out; // @[Top_1.scala 63:50]
  wire [31:0] TRI_RAM_z_io_v11_out; // @[Top_1.scala 63:50]
  wire [31:0] TRI_RAM_z_io_v22_out; // @[Top_1.scala 63:50]
  wire  TRI_RAM_w_clock; // @[Top_1.scala 64:49]
  wire [31:0] TRI_RAM_w_io_Triangle_id; // @[Top_1.scala 64:49]
  wire [31:0] TRI_RAM_w_io_v00_out; // @[Top_1.scala 64:49]
  wire [31:0] TRI_RAM_w_io_v11_out; // @[Top_1.scala 64:49]
  wire [31:0] TRI_RAM_w_io_v22_out; // @[Top_1.scala 64:49]
  wire  RAY_AABB_clock; // @[Top_1.scala 65:46]
  wire  RAY_AABB_reset; // @[Top_1.scala 65:46]
  wire [31:0] RAY_AABB_io_ray_idir_x; // @[Top_1.scala 65:46]
  wire [31:0] RAY_AABB_io_ray_idir_y; // @[Top_1.scala 65:46]
  wire [31:0] RAY_AABB_io_ray_idir_z; // @[Top_1.scala 65:46]
  wire [31:0] RAY_AABB_io_ray_ood_x; // @[Top_1.scala 65:46]
  wire [31:0] RAY_AABB_io_ray_ood_y; // @[Top_1.scala 65:46]
  wire [31:0] RAY_AABB_io_ray_ood_z; // @[Top_1.scala 65:46]
  wire [31:0] RAY_AABB_io_ray_hitT; // @[Top_1.scala 65:46]
  wire [31:0] RAY_AABB_io_bvh_n0xy_x; // @[Top_1.scala 65:46]
  wire [31:0] RAY_AABB_io_bvh_n0xy_y; // @[Top_1.scala 65:46]
  wire [31:0] RAY_AABB_io_bvh_n0xy_z; // @[Top_1.scala 65:46]
  wire [31:0] RAY_AABB_io_bvh_n0xy_w; // @[Top_1.scala 65:46]
  wire [31:0] RAY_AABB_io_bvh_n1xy_x; // @[Top_1.scala 65:46]
  wire [31:0] RAY_AABB_io_bvh_n1xy_y; // @[Top_1.scala 65:46]
  wire [31:0] RAY_AABB_io_bvh_n1xy_z; // @[Top_1.scala 65:46]
  wire [31:0] RAY_AABB_io_bvh_n1xy_w; // @[Top_1.scala 65:46]
  wire [31:0] RAY_AABB_io_bvh_nz_x; // @[Top_1.scala 65:46]
  wire [31:0] RAY_AABB_io_bvh_nz_y; // @[Top_1.scala 65:46]
  wire [31:0] RAY_AABB_io_bvh_nz_z; // @[Top_1.scala 65:46]
  wire [31:0] RAY_AABB_io_bvh_nz_w; // @[Top_1.scala 65:46]
  wire [31:0] RAY_AABB_io_bvh_temp_x; // @[Top_1.scala 65:46]
  wire [31:0] RAY_AABB_io_bvh_temp_y; // @[Top_1.scala 65:46]
  wire [31:0] RAY_AABB_io_rayid; // @[Top_1.scala 65:46]
  wire  RAY_AABB_io_valid_en; // @[Top_1.scala 65:46]
  wire [31:0] RAY_AABB_io_rayid_out; // @[Top_1.scala 65:46]
  wire [31:0] RAY_AABB_io_nodeIdx_0; // @[Top_1.scala 65:46]
  wire [31:0] RAY_AABB_io_nodeIdx_1; // @[Top_1.scala 65:46]
  wire [31:0] RAY_AABB_io_nodeIdx_2; // @[Top_1.scala 65:46]
  wire  RAY_AABB_io_push; // @[Top_1.scala 65:46]
  wire  RAY_AABB_io_pop; // @[Top_1.scala 65:46]
  wire  RAY_AABB_io_leaf; // @[Top_1.scala 65:46]
  wire  RAY_AABB_io_back; // @[Top_1.scala 65:46]
  wire [31:0] RAY_AABB_io_hitT_out; // @[Top_1.scala 65:46]
  wire  RAY_AABB_io_valid_out; // @[Top_1.scala 65:46]
  wire  RAY_AABB_2_clock; // @[Top_1.scala 66:48]
  wire  RAY_AABB_2_reset; // @[Top_1.scala 66:48]
  wire [31:0] RAY_AABB_2_io_ray_idir_x; // @[Top_1.scala 66:48]
  wire [31:0] RAY_AABB_2_io_ray_idir_y; // @[Top_1.scala 66:48]
  wire [31:0] RAY_AABB_2_io_ray_idir_z; // @[Top_1.scala 66:48]
  wire [31:0] RAY_AABB_2_io_ray_ood_x; // @[Top_1.scala 66:48]
  wire [31:0] RAY_AABB_2_io_ray_ood_y; // @[Top_1.scala 66:48]
  wire [31:0] RAY_AABB_2_io_ray_ood_z; // @[Top_1.scala 66:48]
  wire [31:0] RAY_AABB_2_io_ray_hitT; // @[Top_1.scala 66:48]
  wire [31:0] RAY_AABB_2_io_bvh_n0xy_x; // @[Top_1.scala 66:48]
  wire [31:0] RAY_AABB_2_io_bvh_n0xy_y; // @[Top_1.scala 66:48]
  wire [31:0] RAY_AABB_2_io_bvh_n0xy_z; // @[Top_1.scala 66:48]
  wire [31:0] RAY_AABB_2_io_bvh_n0xy_w; // @[Top_1.scala 66:48]
  wire [31:0] RAY_AABB_2_io_bvh_n1xy_x; // @[Top_1.scala 66:48]
  wire [31:0] RAY_AABB_2_io_bvh_n1xy_y; // @[Top_1.scala 66:48]
  wire [31:0] RAY_AABB_2_io_bvh_n1xy_z; // @[Top_1.scala 66:48]
  wire [31:0] RAY_AABB_2_io_bvh_n1xy_w; // @[Top_1.scala 66:48]
  wire [31:0] RAY_AABB_2_io_bvh_nz_x; // @[Top_1.scala 66:48]
  wire [31:0] RAY_AABB_2_io_bvh_nz_y; // @[Top_1.scala 66:48]
  wire [31:0] RAY_AABB_2_io_bvh_nz_z; // @[Top_1.scala 66:48]
  wire [31:0] RAY_AABB_2_io_bvh_nz_w; // @[Top_1.scala 66:48]
  wire [31:0] RAY_AABB_2_io_bvh_temp_x; // @[Top_1.scala 66:48]
  wire [31:0] RAY_AABB_2_io_bvh_temp_y; // @[Top_1.scala 66:48]
  wire [31:0] RAY_AABB_2_io_rayid; // @[Top_1.scala 66:48]
  wire  RAY_AABB_2_io_valid_en; // @[Top_1.scala 66:48]
  wire [31:0] RAY_AABB_2_io_rayid_out; // @[Top_1.scala 66:48]
  wire [31:0] RAY_AABB_2_io_nodeIdx_0; // @[Top_1.scala 66:48]
  wire [31:0] RAY_AABB_2_io_nodeIdx_1; // @[Top_1.scala 66:48]
  wire [31:0] RAY_AABB_2_io_nodeIdx_2; // @[Top_1.scala 66:48]
  wire  RAY_AABB_2_io_push; // @[Top_1.scala 66:48]
  wire  RAY_AABB_2_io_pop; // @[Top_1.scala 66:48]
  wire  RAY_AABB_2_io_leaf; // @[Top_1.scala 66:48]
  wire  RAY_AABB_2_io_back; // @[Top_1.scala 66:48]
  wire [31:0] RAY_AABB_2_io_hitT_out; // @[Top_1.scala 66:48]
  wire  RAY_AABB_2_io_valid_out; // @[Top_1.scala 66:48]
  wire  Arbitration_1_clock; // @[Top_1.scala 67:50]
  wire  Arbitration_1_reset; // @[Top_1.scala 67:50]
  wire [31:0] Arbitration_1_io_node_id_0; // @[Top_1.scala 67:50]
  wire [63:0] Arbitration_1_io_ray_id_0; // @[Top_1.scala 67:50]
  wire [31:0] Arbitration_1_io_hit_0; // @[Top_1.scala 67:50]
  wire  Arbitration_1_io_valid_0; // @[Top_1.scala 67:50]
  wire [31:0] Arbitration_1_io_node_id_1; // @[Top_1.scala 67:50]
  wire [31:0] Arbitration_1_io_ray_id_1; // @[Top_1.scala 67:50]
  wire  Arbitration_1_io_valid_1; // @[Top_1.scala 67:50]
  wire [31:0] Arbitration_1_io_ray_id_2; // @[Top_1.scala 67:50]
  wire  Arbitration_1_io_valid_2; // @[Top_1.scala 67:50]
  wire [31:0] Arbitration_1_io_node_id_out; // @[Top_1.scala 67:50]
  wire [31:0] Arbitration_1_io_ray_id_out; // @[Top_1.scala 67:50]
  wire [31:0] Arbitration_1_io_hit_out; // @[Top_1.scala 67:50]
  wire  Arbitration_1_io_valid_out; // @[Top_1.scala 67:50]
  wire  Arbitration_1_2_clock; // @[Top_1.scala 68:47]
  wire  Arbitration_1_2_reset; // @[Top_1.scala 68:47]
  wire [31:0] Arbitration_1_2_io_node_id_0; // @[Top_1.scala 68:47]
  wire [63:0] Arbitration_1_2_io_ray_id_0; // @[Top_1.scala 68:47]
  wire [31:0] Arbitration_1_2_io_hit_0; // @[Top_1.scala 68:47]
  wire  Arbitration_1_2_io_valid_0; // @[Top_1.scala 68:47]
  wire [31:0] Arbitration_1_2_io_node_id_1; // @[Top_1.scala 68:47]
  wire [31:0] Arbitration_1_2_io_ray_id_1; // @[Top_1.scala 68:47]
  wire  Arbitration_1_2_io_valid_1; // @[Top_1.scala 68:47]
  wire [31:0] Arbitration_1_2_io_ray_id_2; // @[Top_1.scala 68:47]
  wire  Arbitration_1_2_io_valid_2; // @[Top_1.scala 68:47]
  wire [31:0] Arbitration_1_2_io_node_id_out; // @[Top_1.scala 68:47]
  wire [31:0] Arbitration_1_2_io_ray_id_out; // @[Top_1.scala 68:47]
  wire [31:0] Arbitration_1_2_io_hit_out; // @[Top_1.scala 68:47]
  wire  Arbitration_1_2_io_valid_out; // @[Top_1.scala 68:47]
  wire  Arbitration_2_clock; // @[Top_1.scala 70:45]
  wire  Arbitration_2_reset; // @[Top_1.scala 70:45]
  wire [31:0] Arbitration_2_io_ray_id_2_0; // @[Top_1.scala 70:45]
  wire [31:0] Arbitration_2_io_hit_2_0; // @[Top_1.scala 70:45]
  wire  Arbitration_2_io_valid_2_0; // @[Top_1.scala 70:45]
  wire [31:0] Arbitration_2_io_ray_id_2_1; // @[Top_1.scala 70:45]
  wire [31:0] Arbitration_2_io_hit_2_1; // @[Top_1.scala 70:45]
  wire  Arbitration_2_io_valid_2_1; // @[Top_1.scala 70:45]
  wire [31:0] Arbitration_2_io_ray_id_2_2; // @[Top_1.scala 70:45]
  wire [31:0] Arbitration_2_io_hit_2_2; // @[Top_1.scala 70:45]
  wire  Arbitration_2_io_valid_2_2; // @[Top_1.scala 70:45]
  wire [31:0] Arbitration_2_io_ray_id_2_3; // @[Top_1.scala 70:45]
  wire [31:0] Arbitration_2_io_hit_2_3; // @[Top_1.scala 70:45]
  wire  Arbitration_2_io_valid_2_3; // @[Top_1.scala 70:45]
  wire [31:0] Arbitration_2_io_ray_id_out; // @[Top_1.scala 70:45]
  wire [31:0] Arbitration_2_io_hit_out; // @[Top_1.scala 70:45]
  wire  Arbitration_2_io_valid_out; // @[Top_1.scala 70:45]
  wire  Arbitration_2_2_clock; // @[Top_1.scala 71:42]
  wire  Arbitration_2_2_reset; // @[Top_1.scala 71:42]
  wire [31:0] Arbitration_2_2_io_ray_id_2_0; // @[Top_1.scala 71:42]
  wire [31:0] Arbitration_2_2_io_hit_2_0; // @[Top_1.scala 71:42]
  wire  Arbitration_2_2_io_valid_2_0; // @[Top_1.scala 71:42]
  wire [31:0] Arbitration_2_2_io_ray_id_2_1; // @[Top_1.scala 71:42]
  wire [31:0] Arbitration_2_2_io_hit_2_1; // @[Top_1.scala 71:42]
  wire  Arbitration_2_2_io_valid_2_1; // @[Top_1.scala 71:42]
  wire [31:0] Arbitration_2_2_io_ray_id_2_2; // @[Top_1.scala 71:42]
  wire [31:0] Arbitration_2_2_io_hit_2_2; // @[Top_1.scala 71:42]
  wire  Arbitration_2_2_io_valid_2_2; // @[Top_1.scala 71:42]
  wire [31:0] Arbitration_2_2_io_ray_id_2_3; // @[Top_1.scala 71:42]
  wire [31:0] Arbitration_2_2_io_hit_2_3; // @[Top_1.scala 71:42]
  wire  Arbitration_2_2_io_valid_2_3; // @[Top_1.scala 71:42]
  wire [31:0] Arbitration_2_2_io_ray_id_out; // @[Top_1.scala 71:42]
  wire [31:0] Arbitration_2_2_io_hit_out; // @[Top_1.scala 71:42]
  wire  Arbitration_2_2_io_valid_out; // @[Top_1.scala 71:42]
  wire  Arbitration_3_clock; // @[Top_1.scala 72:45]
  wire  Arbitration_3_reset; // @[Top_1.scala 72:45]
  wire [31:0] Arbitration_3_io_node_id_3_0; // @[Top_1.scala 72:45]
  wire [31:0] Arbitration_3_io_ray_id_3_0; // @[Top_1.scala 72:45]
  wire [31:0] Arbitration_3_io_hit_3_0; // @[Top_1.scala 72:45]
  wire  Arbitration_3_io_valid_3_0; // @[Top_1.scala 72:45]
  wire [31:0] Arbitration_3_io_node_id_3_1; // @[Top_1.scala 72:45]
  wire [31:0] Arbitration_3_io_ray_id_3_1; // @[Top_1.scala 72:45]
  wire [31:0] Arbitration_3_io_hit_3_1; // @[Top_1.scala 72:45]
  wire  Arbitration_3_io_valid_3_1; // @[Top_1.scala 72:45]
  wire [31:0] Arbitration_3_io_node_id_3_2; // @[Top_1.scala 72:45]
  wire [31:0] Arbitration_3_io_ray_id_3_2; // @[Top_1.scala 72:45]
  wire [31:0] Arbitration_3_io_hit_3_2; // @[Top_1.scala 72:45]
  wire  Arbitration_3_io_valid_3_2; // @[Top_1.scala 72:45]
  wire [31:0] Arbitration_3_io_node_id_3_3; // @[Top_1.scala 72:45]
  wire [31:0] Arbitration_3_io_ray_id_3_3; // @[Top_1.scala 72:45]
  wire [31:0] Arbitration_3_io_hit_3_3; // @[Top_1.scala 72:45]
  wire  Arbitration_3_io_valid_3_3; // @[Top_1.scala 72:45]
  wire [31:0] Arbitration_3_io_node_id_3_4; // @[Top_1.scala 72:45]
  wire [31:0] Arbitration_3_io_ray_id_3_4; // @[Top_1.scala 72:45]
  wire [31:0] Arbitration_3_io_hit_3_4; // @[Top_1.scala 72:45]
  wire  Arbitration_3_io_valid_3_4; // @[Top_1.scala 72:45]
  wire [31:0] Arbitration_3_io_node_id_out; // @[Top_1.scala 72:45]
  wire [31:0] Arbitration_3_io_ray_id_out; // @[Top_1.scala 72:45]
  wire [31:0] Arbitration_3_io_hit_out; // @[Top_1.scala 72:45]
  wire  Arbitration_3_io_valid_out; // @[Top_1.scala 72:45]
  wire  Arbitration_3_2_clock; // @[Top_1.scala 73:42]
  wire  Arbitration_3_2_reset; // @[Top_1.scala 73:42]
  wire [31:0] Arbitration_3_2_io_node_id_3_0; // @[Top_1.scala 73:42]
  wire [31:0] Arbitration_3_2_io_ray_id_3_0; // @[Top_1.scala 73:42]
  wire [31:0] Arbitration_3_2_io_hit_3_0; // @[Top_1.scala 73:42]
  wire  Arbitration_3_2_io_valid_3_0; // @[Top_1.scala 73:42]
  wire [31:0] Arbitration_3_2_io_node_id_3_1; // @[Top_1.scala 73:42]
  wire [31:0] Arbitration_3_2_io_ray_id_3_1; // @[Top_1.scala 73:42]
  wire [31:0] Arbitration_3_2_io_hit_3_1; // @[Top_1.scala 73:42]
  wire  Arbitration_3_2_io_valid_3_1; // @[Top_1.scala 73:42]
  wire [31:0] Arbitration_3_2_io_node_id_3_2; // @[Top_1.scala 73:42]
  wire [31:0] Arbitration_3_2_io_ray_id_3_2; // @[Top_1.scala 73:42]
  wire [31:0] Arbitration_3_2_io_hit_3_2; // @[Top_1.scala 73:42]
  wire  Arbitration_3_2_io_valid_3_2; // @[Top_1.scala 73:42]
  wire [31:0] Arbitration_3_2_io_node_id_3_3; // @[Top_1.scala 73:42]
  wire [31:0] Arbitration_3_2_io_ray_id_3_3; // @[Top_1.scala 73:42]
  wire [31:0] Arbitration_3_2_io_hit_3_3; // @[Top_1.scala 73:42]
  wire  Arbitration_3_2_io_valid_3_3; // @[Top_1.scala 73:42]
  wire [31:0] Arbitration_3_2_io_node_id_3_4; // @[Top_1.scala 73:42]
  wire [31:0] Arbitration_3_2_io_ray_id_3_4; // @[Top_1.scala 73:42]
  wire [31:0] Arbitration_3_2_io_hit_3_4; // @[Top_1.scala 73:42]
  wire  Arbitration_3_2_io_valid_3_4; // @[Top_1.scala 73:42]
  wire [31:0] Arbitration_3_2_io_node_id_out; // @[Top_1.scala 73:42]
  wire [31:0] Arbitration_3_2_io_ray_id_out; // @[Top_1.scala 73:42]
  wire [31:0] Arbitration_3_2_io_hit_out; // @[Top_1.scala 73:42]
  wire  Arbitration_3_2_io_valid_out; // @[Top_1.scala 73:42]
  wire  Arbitration_4_clock; // @[Top_1.scala 74:45]
  wire  Arbitration_4_reset; // @[Top_1.scala 74:45]
  wire [31:0] Arbitration_4_io_node_id_4_0; // @[Top_1.scala 74:45]
  wire [31:0] Arbitration_4_io_ray_id_4_0; // @[Top_1.scala 74:45]
  wire [31:0] Arbitration_4_io_hit_4_0; // @[Top_1.scala 74:45]
  wire  Arbitration_4_io_valid_4_0; // @[Top_1.scala 74:45]
  wire [31:0] Arbitration_4_io_node_id_4_1; // @[Top_1.scala 74:45]
  wire [31:0] Arbitration_4_io_ray_id_4_1; // @[Top_1.scala 74:45]
  wire [31:0] Arbitration_4_io_hit_4_1; // @[Top_1.scala 74:45]
  wire  Arbitration_4_io_valid_4_1; // @[Top_1.scala 74:45]
  wire [31:0] Arbitration_4_io_node_id_out; // @[Top_1.scala 74:45]
  wire [31:0] Arbitration_4_io_ray_id_out; // @[Top_1.scala 74:45]
  wire [31:0] Arbitration_4_io_hit_out; // @[Top_1.scala 74:45]
  wire  Arbitration_4_io_RAY_AABB_out; // @[Top_1.scala 74:45]
  wire  Arbitration_4_io_RAY_AABB_2_out; // @[Top_1.scala 74:45]
  wire  Arbitration_4_io_valid_out; // @[Top_1.scala 74:45]
  wire  Stack_manage_clock; // @[Top_1.scala 75:41]
  wire  Stack_manage_reset; // @[Top_1.scala 75:41]
  wire  Stack_manage_io_push; // @[Top_1.scala 75:41]
  wire  Stack_manage_io_push_en; // @[Top_1.scala 75:41]
  wire  Stack_manage_io_pop; // @[Top_1.scala 75:41]
  wire  Stack_manage_io_pop_en; // @[Top_1.scala 75:41]
  wire [31:0] Stack_manage_io_ray_id_push; // @[Top_1.scala 75:41]
  wire [31:0] Stack_manage_io_ray_id_pop; // @[Top_1.scala 75:41]
  wire [31:0] Stack_manage_io_node_id_push_in; // @[Top_1.scala 75:41]
  wire [31:0] Stack_manage_io_hitT_in; // @[Top_1.scala 75:41]
  wire [31:0] Stack_manage_io_hitT_out; // @[Top_1.scala 75:41]
  wire [31:0] Stack_manage_io_node_id_out; // @[Top_1.scala 75:41]
  wire [31:0] Stack_manage_io_ray_id_out; // @[Top_1.scala 75:41]
  wire  Stack_manage_io_pop_valid; // @[Top_1.scala 75:41]
  wire  Stack_manage_io_Dis_en; // @[Top_1.scala 75:41]
  wire  Stack_manage_io_Finish; // @[Top_1.scala 75:41]
  wire  Stack_manage_2_clock; // @[Top_1.scala 76:38]
  wire  Stack_manage_2_reset; // @[Top_1.scala 76:38]
  wire  Stack_manage_2_io_push; // @[Top_1.scala 76:38]
  wire  Stack_manage_2_io_push_en; // @[Top_1.scala 76:38]
  wire  Stack_manage_2_io_pop; // @[Top_1.scala 76:38]
  wire  Stack_manage_2_io_pop_en; // @[Top_1.scala 76:38]
  wire [31:0] Stack_manage_2_io_ray_id_push; // @[Top_1.scala 76:38]
  wire [31:0] Stack_manage_2_io_ray_id_pop; // @[Top_1.scala 76:38]
  wire [31:0] Stack_manage_2_io_node_id_push_in; // @[Top_1.scala 76:38]
  wire [31:0] Stack_manage_2_io_hitT_in; // @[Top_1.scala 76:38]
  wire [31:0] Stack_manage_2_io_hitT_out; // @[Top_1.scala 76:38]
  wire [31:0] Stack_manage_2_io_node_id_out; // @[Top_1.scala 76:38]
  wire [31:0] Stack_manage_2_io_ray_id_out; // @[Top_1.scala 76:38]
  wire  Stack_manage_2_io_pop_valid; // @[Top_1.scala 76:38]
  wire  Stack_manage_2_io_Dis_en; // @[Top_1.scala 76:38]
  wire  Stack_manage_2_io_Finish; // @[Top_1.scala 76:38]
  wire  Triangle_clock; // @[Top_1.scala 77:51]
  wire  Triangle_reset; // @[Top_1.scala 77:51]
  wire  Triangle_io_To_IST0_enable; // @[Top_1.scala 77:51]
  wire [31:0] Triangle_io_nodeid_leaf; // @[Top_1.scala 77:51]
  wire [31:0] Triangle_io_rayid_leaf; // @[Top_1.scala 77:51]
  wire [31:0] Triangle_io_hiT_in; // @[Top_1.scala 77:51]
  wire [31:0] Triangle_io_v00_in_x; // @[Top_1.scala 77:51]
  wire [31:0] Triangle_io_v00_in_y; // @[Top_1.scala 77:51]
  wire [31:0] Triangle_io_v00_in_z; // @[Top_1.scala 77:51]
  wire [31:0] Triangle_io_v00_in_w; // @[Top_1.scala 77:51]
  wire [31:0] Triangle_io_v11_in_x; // @[Top_1.scala 77:51]
  wire [31:0] Triangle_io_v11_in_y; // @[Top_1.scala 77:51]
  wire [31:0] Triangle_io_v11_in_z; // @[Top_1.scala 77:51]
  wire [31:0] Triangle_io_v11_in_w; // @[Top_1.scala 77:51]
  wire [31:0] Triangle_io_v22_in_x; // @[Top_1.scala 77:51]
  wire [31:0] Triangle_io_v22_in_y; // @[Top_1.scala 77:51]
  wire [31:0] Triangle_io_v22_in_z; // @[Top_1.scala 77:51]
  wire [31:0] Triangle_io_v22_in_w; // @[Top_1.scala 77:51]
  wire [31:0] Triangle_io_ray_o_in_x; // @[Top_1.scala 77:51]
  wire [31:0] Triangle_io_ray_o_in_y; // @[Top_1.scala 77:51]
  wire [31:0] Triangle_io_ray_o_in_z; // @[Top_1.scala 77:51]
  wire [31:0] Triangle_io_ray_d_in_x; // @[Top_1.scala 77:51]
  wire [31:0] Triangle_io_ray_d_in_y; // @[Top_1.scala 77:51]
  wire [31:0] Triangle_io_ray_d_in_z; // @[Top_1.scala 77:51]
  wire  Triangle_io_break_in; // @[Top_1.scala 77:51]
  wire  Triangle_io_RAY_AABB_1; // @[Top_1.scala 77:51]
  wire  Triangle_io_RAY_AABB_2; // @[Top_1.scala 77:51]
  wire  Triangle_io_pop_1; // @[Top_1.scala 77:51]
  wire  Triangle_io_break_1; // @[Top_1.scala 77:51]
  wire  Triangle_io_pop_2; // @[Top_1.scala 77:51]
  wire  Triangle_io_break_2; // @[Top_1.scala 77:51]
  wire  Triangle_io_pop_3; // @[Top_1.scala 77:51]
  wire  Triangle_io_break_3; // @[Top_1.scala 77:51]
  wire [31:0] Triangle_io_hiT_out_1; // @[Top_1.scala 77:51]
  wire [31:0] Triangle_io_hiT_out_2; // @[Top_1.scala 77:51]
  wire [31:0] Triangle_io_hiT_out_3; // @[Top_1.scala 77:51]
  wire  Triangle_io_hitT_en; // @[Top_1.scala 77:51]
  wire [31:0] Triangle_io_hitIndex; // @[Top_1.scala 77:51]
  wire [31:0] Triangle_io_node_id_out_1; // @[Top_1.scala 77:51]
  wire [31:0] Triangle_io_node_id_out_2; // @[Top_1.scala 77:51]
  wire [31:0] Triangle_io_node_id_out_3; // @[Top_1.scala 77:51]
  wire [31:0] Triangle_io_ray_id_ist1; // @[Top_1.scala 77:51]
  wire [31:0] Triangle_io_ray_id_ist2; // @[Top_1.scala 77:51]
  wire [31:0] Triangle_io_ray_id_ist3; // @[Top_1.scala 77:51]
  wire [63:0] Triangle_io_counter_fdiv; // @[Top_1.scala 77:51]
  wire  Triangle_io_RAY_AABB_1_out_IST1; // @[Top_1.scala 77:51]
  wire  Triangle_io_RAY_AABB_2_out_IST1; // @[Top_1.scala 77:51]
  wire  Triangle_io_RAY_AABB_1_out_IST2; // @[Top_1.scala 77:51]
  wire  Triangle_io_RAY_AABB_2_out_IST2; // @[Top_1.scala 77:51]
  wire  Triangle_io_RAY_AABB_1_out_IST3; // @[Top_1.scala 77:51]
  wire  Triangle_io_RAY_AABB_2_out_IST3; // @[Top_1.scala 77:51]
  reg [63:0] clock_counter; // @[Top_1.scala 79:42]
  wire [63:0] _T_1 = clock_counter + 64'h1; // @[Top_1.scala 80:53]
  reg  memory_valid; // @[Top_1.scala 129:54]
  reg [31:0] hit_temp; // @[Top_1.scala 130:61]
  reg [31:0] ray_id_temp; // @[Top_1.scala 131:57]
  reg  hit_from_arb; // @[Top_1.scala 132:57]
  reg [63:0] TRV_1; // @[Top_1.scala 133:64]
  wire  _T_8 = Arbitration_1_io_valid_out & Arbitration_1_io_hit_out != 32'h0; // @[Top_1.scala 134:36]
  wire [32:0] _T_9 = $signed(Arbitration_1_io_node_id_out) / 32'sh4; // @[Top_1.scala 143:75]
  wire  _T_24 = Arbitration_1_io_valid_out & Arbitration_1_io_hit_out == 32'h0; // @[Top_1.scala 159:42]
  wire [31:0] _GEN_13 = Arbitration_1_io_ray_id_out; // @[Top_1.scala 159:76 Top_1.scala 161:53]
  wire  _GEN_31 = Arbitration_1_io_valid_out & Arbitration_1_io_hit_out != 32'h0 | _T_24; // @[Top_1.scala 134:70 Top_1.scala 135:51]
  wire [32:0] _GEN_34 = Arbitration_1_io_valid_out & Arbitration_1_io_hit_out != 32'h0 ? $signed(_T_9) : $signed(_T_9); // @[Top_1.scala 134:70 Top_1.scala 143:44]
  wire [31:0] _GEN_51 = hit_from_arb ? hit_temp : Ray_hitT_io_Ray_out; // @[Top_1.scala 198:33 Top_1.scala 199:53 Top_1.scala 201:53]
  wire [63:0] _T_42 = TRV_1 + 64'h1; // @[Top_1.scala 222:79]
  reg  memory_valid_2; // @[Top_1.scala 264:56]
  reg [31:0] hit_temp_2; // @[Top_1.scala 265:63]
  reg [31:0] ray_id_temp_2; // @[Top_1.scala 266:59]
  reg  hit_from_arb_2; // @[Top_1.scala 267:59]
  reg [63:0] TRV_2; // @[Top_1.scala 268:70]
  wire  _T_45 = Arbitration_1_2_io_valid_out & Arbitration_1_2_io_hit_out != 32'h0; // @[Top_1.scala 269:38]
  wire [32:0] _T_46 = $signed(Arbitration_1_2_io_node_id_out) / 32'sh4; // @[Top_1.scala 280:79]
  wire  _T_61 = Arbitration_1_2_io_valid_out & Arbitration_1_2_io_hit_out == 32'h0; // @[Top_1.scala 296:44]
  wire [31:0] _GEN_81 = Arbitration_1_2_io_ray_id_out; // @[Top_1.scala 296:80 Top_1.scala 300:54]
  wire  _GEN_98 = Arbitration_1_2_io_valid_out & Arbitration_1_2_io_hit_out != 32'h0 | _T_61; // @[Top_1.scala 269:74 Top_1.scala 270:58]
  wire [32:0] _GEN_101 = Arbitration_1_2_io_valid_out & Arbitration_1_2_io_hit_out != 32'h0 ? $signed(_T_46) : $signed(
    _T_46); // @[Top_1.scala 269:74 Top_1.scala 280:46]
  wire [31:0] _GEN_118 = hit_from_arb_2 ? hit_temp_2 : Ray_hitT_io_Ray_out_2; // @[Top_1.scala 337:35 Top_1.scala 338:55 Top_1.scala 340:55]
  wire [63:0] _T_79 = TRV_2 + 64'h1; // @[Top_1.scala 358:85]
  wire  hi = ~RAY_AABB_io_nodeIdx_2[31]; // @[common.scala 128:29]
  wire [30:0] lo = ~RAY_AABB_io_nodeIdx_2[30:0]; // @[common.scala 128:45]
  wire [31:0] _T_88 = {hi,lo}; // @[common.scala 128:56]
  wire  hi_1 = ~RAY_AABB_2_io_nodeIdx_2[31]; // @[common.scala 128:29]
  wire [30:0] lo_1 = ~RAY_AABB_2_io_nodeIdx_2[30:0]; // @[common.scala 128:45]
  wire [31:0] _T_94 = {hi_1,lo_1}; // @[common.scala 128:56]
  wire  _T_96 = ~Stack_manage_io_node_id_out[31]; // @[common.scala 100:25]
  wire [30:0] lo_2 = ~Stack_manage_io_node_id_out[30:0]; // @[common.scala 128:45]
  wire [31:0] _T_109 = {_T_96,lo_2}; // @[common.scala 128:56]
  wire [31:0] _GEN_168 = _T_96 & Stack_manage_io_pop_valid ? Stack_manage_io_ray_id_out : 32'h0; // @[Top_1.scala 451:81 Top_1.scala 453:50]
  wire  _T_111 = ~Stack_manage_2_io_node_id_out[31]; // @[common.scala 100:25]
  wire [30:0] lo_3 = ~Stack_manage_2_io_node_id_out[30:0]; // @[common.scala 128:45]
  wire [31:0] _T_124 = {_T_111,lo_3}; // @[common.scala 128:56]
  wire [31:0] _GEN_182 = _T_111 & Stack_manage_2_io_pop_valid ? Stack_manage_2_io_ray_id_out : 32'h0; // @[Top_1.scala 471:85 Top_1.scala 473:52]
  wire [31:0] _T_128 = $signed(Triangle_io_node_id_out_1) + 32'sh3; // @[Top_1.scala 517:71]
  wire [31:0] _T_136 = $signed(Triangle_io_node_id_out_2) + 32'sh3; // @[Top_1.scala 542:71]
  wire [31:0] _T_144 = $signed(Triangle_io_node_id_out_3) + 32'sh3; // @[Top_1.scala 566:71]
  reg  leaf_memory_valid; // @[Top_1.scala 666:58]
  reg [31:0] hitT_temp; // @[Top_1.scala 667:68]
  reg [31:0] ray_leaf_temp; // @[Top_1.scala 668:64]
  reg [31:0] leaf_node_id_temp; // @[Top_1.scala 669:57]
  reg  ray_aabb; // @[Top_1.scala 670:69]
  reg  ray_aabb_2; // @[Top_1.scala 671:71]
  reg [63:0] IST_1; // @[Top_1.scala 672:75]
  wire  _GEN_239 = Arbitration_4_io_valid_out; // @[Top_1.scala 673:37 Top_1.scala 674:50 Top_1.scala 691:50]
  wire  _GEN_245 = Arbitration_4_io_valid_out & Arbitration_4_io_RAY_AABB_out; // @[Top_1.scala 673:37 Top_1.scala 688:64 Top_1.scala 695:64]
  wire  _GEN_246 = Arbitration_4_io_valid_out & Arbitration_4_io_RAY_AABB_2_out; // @[Top_1.scala 673:37 Top_1.scala 689:61 Top_1.scala 696:61]
  wire [63:0] _T_159 = IST_1 + 64'h1; // @[Top_1.scala 724:76]
  ray_dispatch Ray_Dispatch ( // @[Top_1.scala 24:44]
    .clock(Ray_Dispatch_clock),
    .reset(Ray_Dispatch_reset),
    .io_dispatch(Ray_Dispatch_io_dispatch),
    .io_dispatch_2(Ray_Dispatch_io_dispatch_2),
    .io_rayid_id(Ray_Dispatch_io_rayid_id),
    .io_rayid_id_2(Ray_Dispatch_io_rayid_id_2),
    .io_ray_out(Ray_Dispatch_io_ray_out),
    .io_ray_out_2(Ray_Dispatch_io_ray_out_2),
    .io_ray_finish(Ray_Dispatch_io_ray_finish)
  );
  ray_memory Ray_origx ( // @[Top_1.scala 25:48]
    .clock(Ray_origx_clock),
    .io_Ray_id(Ray_origx_io_Ray_id),
    .io_Ray_id_2(Ray_origx_io_Ray_id_2),
    .io_Ray_out(Ray_origx_io_Ray_out),
    .io_Ray_out_2(Ray_origx_io_Ray_out_2)
  );
  ray_memory Ray_origy ( // @[Top_1.scala 26:48]
    .clock(Ray_origy_clock),
    .io_Ray_id(Ray_origy_io_Ray_id),
    .io_Ray_id_2(Ray_origy_io_Ray_id_2),
    .io_Ray_out(Ray_origy_io_Ray_out),
    .io_Ray_out_2(Ray_origy_io_Ray_out_2)
  );
  ray_memory Ray_origz ( // @[Top_1.scala 27:48]
    .clock(Ray_origz_clock),
    .io_Ray_id(Ray_origz_io_Ray_id),
    .io_Ray_id_2(Ray_origz_io_Ray_id_2),
    .io_Ray_out(Ray_origz_io_Ray_out),
    .io_Ray_out_2(Ray_origz_io_Ray_out_2)
  );
  ray_memory Ray_dirx ( // @[Top_1.scala 30:50]
    .clock(Ray_dirx_clock),
    .io_Ray_id(Ray_dirx_io_Ray_id),
    .io_Ray_id_2(Ray_dirx_io_Ray_id_2),
    .io_Ray_out(Ray_dirx_io_Ray_out),
    .io_Ray_out_2(Ray_dirx_io_Ray_out_2)
  );
  ray_memory Ray_diry ( // @[Top_1.scala 31:49]
    .clock(Ray_diry_clock),
    .io_Ray_id(Ray_diry_io_Ray_id),
    .io_Ray_id_2(Ray_diry_io_Ray_id_2),
    .io_Ray_out(Ray_diry_io_Ray_out),
    .io_Ray_out_2(Ray_diry_io_Ray_out_2)
  );
  ray_memory Ray_dirz ( // @[Top_1.scala 32:49]
    .clock(Ray_dirz_clock),
    .io_Ray_id(Ray_dirz_io_Ray_id),
    .io_Ray_id_2(Ray_dirz_io_Ray_id_2),
    .io_Ray_out(Ray_dirz_io_Ray_out),
    .io_Ray_out_2(Ray_dirz_io_Ray_out_2)
  );
  ray_memory Ray_hitT ( // @[Top_1.scala 33:49]
    .clock(Ray_hitT_clock),
    .io_Ray_id(Ray_hitT_io_Ray_id),
    .io_Ray_id_2(Ray_hitT_io_Ray_id_2),
    .io_Ray_out(Ray_hitT_io_Ray_out),
    .io_Ray_out_2(Ray_hitT_io_Ray_out_2)
  );
  ray_memory Ray_idirx ( // @[Top_1.scala 35:49]
    .clock(Ray_idirx_clock),
    .io_Ray_id(Ray_idirx_io_Ray_id),
    .io_Ray_id_2(Ray_idirx_io_Ray_id_2),
    .io_Ray_out(Ray_idirx_io_Ray_out),
    .io_Ray_out_2(Ray_idirx_io_Ray_out_2)
  );
  ray_memory Ray_idiry ( // @[Top_1.scala 36:49]
    .clock(Ray_idiry_clock),
    .io_Ray_id(Ray_idiry_io_Ray_id),
    .io_Ray_id_2(Ray_idiry_io_Ray_id_2),
    .io_Ray_out(Ray_idiry_io_Ray_out),
    .io_Ray_out_2(Ray_idiry_io_Ray_out_2)
  );
  ray_memory Ray_idirz ( // @[Top_1.scala 37:49]
    .clock(Ray_idirz_clock),
    .io_Ray_id(Ray_idirz_io_Ray_id),
    .io_Ray_id_2(Ray_idirz_io_Ray_id_2),
    .io_Ray_out(Ray_idirz_io_Ray_out),
    .io_Ray_out_2(Ray_idirz_io_Ray_out_2)
  );
  ray_memory Ray_oodx ( // @[Top_1.scala 39:48]
    .clock(Ray_oodx_clock),
    .io_Ray_id(Ray_oodx_io_Ray_id),
    .io_Ray_id_2(Ray_oodx_io_Ray_id_2),
    .io_Ray_out(Ray_oodx_io_Ray_out),
    .io_Ray_out_2(Ray_oodx_io_Ray_out_2)
  );
  ray_memory Ray_oody ( // @[Top_1.scala 40:48]
    .clock(Ray_oody_clock),
    .io_Ray_id(Ray_oody_io_Ray_id),
    .io_Ray_id_2(Ray_oody_io_Ray_id_2),
    .io_Ray_out(Ray_oody_io_Ray_out),
    .io_Ray_out_2(Ray_oody_io_Ray_out_2)
  );
  ray_memory Ray_oodz ( // @[Top_1.scala 41:48]
    .clock(Ray_oodz_clock),
    .io_Ray_id(Ray_oodz_io_Ray_id),
    .io_Ray_id_2(Ray_oodz_io_Ray_id_2),
    .io_Ray_out(Ray_oodz_io_Ray_out),
    .io_Ray_out_2(Ray_oodz_io_Ray_out_2)
  );
  BVH_memory BVH_RAM_0_x ( // @[Top_1.scala 43:41]
    .clock(BVH_RAM_0_x_clock),
    .io_BVH_id(BVH_RAM_0_x_io_BVH_id),
    .io_BVH_id_2(BVH_RAM_0_x_io_BVH_id_2),
    .io_BVH_out(BVH_RAM_0_x_io_BVH_out),
    .io_BVH_out_2(BVH_RAM_0_x_io_BVH_out_2)
  );
  BVH_memory BVH_RAM_0_y ( // @[Top_1.scala 44:41]
    .clock(BVH_RAM_0_y_clock),
    .io_BVH_id(BVH_RAM_0_y_io_BVH_id),
    .io_BVH_id_2(BVH_RAM_0_y_io_BVH_id_2),
    .io_BVH_out(BVH_RAM_0_y_io_BVH_out),
    .io_BVH_out_2(BVH_RAM_0_y_io_BVH_out_2)
  );
  BVH_memory BVH_RAM_0_z ( // @[Top_1.scala 45:41]
    .clock(BVH_RAM_0_z_clock),
    .io_BVH_id(BVH_RAM_0_z_io_BVH_id),
    .io_BVH_id_2(BVH_RAM_0_z_io_BVH_id_2),
    .io_BVH_out(BVH_RAM_0_z_io_BVH_out),
    .io_BVH_out_2(BVH_RAM_0_z_io_BVH_out_2)
  );
  BVH_memory BVH_RAM_0_w ( // @[Top_1.scala 46:40]
    .clock(BVH_RAM_0_w_clock),
    .io_BVH_id(BVH_RAM_0_w_io_BVH_id),
    .io_BVH_id_2(BVH_RAM_0_w_io_BVH_id_2),
    .io_BVH_out(BVH_RAM_0_w_io_BVH_out),
    .io_BVH_out_2(BVH_RAM_0_w_io_BVH_out_2)
  );
  BVH_memory BVH_RAM_1_x ( // @[Top_1.scala 48:41]
    .clock(BVH_RAM_1_x_clock),
    .io_BVH_id(BVH_RAM_1_x_io_BVH_id),
    .io_BVH_id_2(BVH_RAM_1_x_io_BVH_id_2),
    .io_BVH_out(BVH_RAM_1_x_io_BVH_out),
    .io_BVH_out_2(BVH_RAM_1_x_io_BVH_out_2)
  );
  BVH_memory BVH_RAM_1_y ( // @[Top_1.scala 49:41]
    .clock(BVH_RAM_1_y_clock),
    .io_BVH_id(BVH_RAM_1_y_io_BVH_id),
    .io_BVH_id_2(BVH_RAM_1_y_io_BVH_id_2),
    .io_BVH_out(BVH_RAM_1_y_io_BVH_out),
    .io_BVH_out_2(BVH_RAM_1_y_io_BVH_out_2)
  );
  BVH_memory BVH_RAM_1_z ( // @[Top_1.scala 50:41]
    .clock(BVH_RAM_1_z_clock),
    .io_BVH_id(BVH_RAM_1_z_io_BVH_id),
    .io_BVH_id_2(BVH_RAM_1_z_io_BVH_id_2),
    .io_BVH_out(BVH_RAM_1_z_io_BVH_out),
    .io_BVH_out_2(BVH_RAM_1_z_io_BVH_out_2)
  );
  BVH_memory BVH_RAM_1_w ( // @[Top_1.scala 51:40]
    .clock(BVH_RAM_1_w_clock),
    .io_BVH_id(BVH_RAM_1_w_io_BVH_id),
    .io_BVH_id_2(BVH_RAM_1_w_io_BVH_id_2),
    .io_BVH_out(BVH_RAM_1_w_io_BVH_out),
    .io_BVH_out_2(BVH_RAM_1_w_io_BVH_out_2)
  );
  BVH_memory BVH_RAM_z_x ( // @[Top_1.scala 53:41]
    .clock(BVH_RAM_z_x_clock),
    .io_BVH_id(BVH_RAM_z_x_io_BVH_id),
    .io_BVH_id_2(BVH_RAM_z_x_io_BVH_id_2),
    .io_BVH_out(BVH_RAM_z_x_io_BVH_out),
    .io_BVH_out_2(BVH_RAM_z_x_io_BVH_out_2)
  );
  BVH_memory BVH_RAM_z_y ( // @[Top_1.scala 54:41]
    .clock(BVH_RAM_z_y_clock),
    .io_BVH_id(BVH_RAM_z_y_io_BVH_id),
    .io_BVH_id_2(BVH_RAM_z_y_io_BVH_id_2),
    .io_BVH_out(BVH_RAM_z_y_io_BVH_out),
    .io_BVH_out_2(BVH_RAM_z_y_io_BVH_out_2)
  );
  BVH_memory BVH_RAM_z_z ( // @[Top_1.scala 55:41]
    .clock(BVH_RAM_z_z_clock),
    .io_BVH_id(BVH_RAM_z_z_io_BVH_id),
    .io_BVH_id_2(BVH_RAM_z_z_io_BVH_id_2),
    .io_BVH_out(BVH_RAM_z_z_io_BVH_out),
    .io_BVH_out_2(BVH_RAM_z_z_io_BVH_out_2)
  );
  BVH_memory BVH_RAM_z_w ( // @[Top_1.scala 56:40]
    .clock(BVH_RAM_z_w_clock),
    .io_BVH_id(BVH_RAM_z_w_io_BVH_id),
    .io_BVH_id_2(BVH_RAM_z_w_io_BVH_id_2),
    .io_BVH_out(BVH_RAM_z_w_io_BVH_out),
    .io_BVH_out_2(BVH_RAM_z_w_io_BVH_out_2)
  );
  BVH_memory_0 BVH_RAM_tmp_x ( // @[Top_1.scala 58:37]
    .clock(BVH_RAM_tmp_x_clock),
    .io_BVH_id(BVH_RAM_tmp_x_io_BVH_id),
    .io_BVH_id_2(BVH_RAM_tmp_x_io_BVH_id_2),
    .io_BVH_out(BVH_RAM_tmp_x_io_BVH_out),
    .io_BVH_out_2(BVH_RAM_tmp_x_io_BVH_out_2)
  );
  BVH_memory_0 BVH_RAM_tmp_y ( // @[Top_1.scala 59:37]
    .clock(BVH_RAM_tmp_y_clock),
    .io_BVH_id(BVH_RAM_tmp_y_io_BVH_id),
    .io_BVH_id_2(BVH_RAM_tmp_y_io_BVH_id_2),
    .io_BVH_out(BVH_RAM_tmp_y_io_BVH_out),
    .io_BVH_out_2(BVH_RAM_tmp_y_io_BVH_out_2)
  );
  Triangle_memory_valid TRI_RAM_x ( // @[Top_1.scala 61:50]
    .clock(TRI_RAM_x_clock),
    .io_Triangle_id(TRI_RAM_x_io_Triangle_id),
    .io_v00_out(TRI_RAM_x_io_v00_out),
    .io_v11_out(TRI_RAM_x_io_v11_out),
    .io_v22_out(TRI_RAM_x_io_v22_out),
    .io_valid(TRI_RAM_x_io_valid)
  );
  Triangle_memory TRI_RAM_y ( // @[Top_1.scala 62:50]
    .clock(TRI_RAM_y_clock),
    .io_Triangle_id(TRI_RAM_y_io_Triangle_id),
    .io_v00_out(TRI_RAM_y_io_v00_out),
    .io_v11_out(TRI_RAM_y_io_v11_out),
    .io_v22_out(TRI_RAM_y_io_v22_out)
  );
  Triangle_memory TRI_RAM_z ( // @[Top_1.scala 63:50]
    .clock(TRI_RAM_z_clock),
    .io_Triangle_id(TRI_RAM_z_io_Triangle_id),
    .io_v00_out(TRI_RAM_z_io_v00_out),
    .io_v11_out(TRI_RAM_z_io_v11_out),
    .io_v22_out(TRI_RAM_z_io_v22_out)
  );
  Triangle_memory TRI_RAM_w ( // @[Top_1.scala 64:49]
    .clock(TRI_RAM_w_clock),
    .io_Triangle_id(TRI_RAM_w_io_Triangle_id),
    .io_v00_out(TRI_RAM_w_io_v00_out),
    .io_v11_out(TRI_RAM_w_io_v11_out),
    .io_v22_out(TRI_RAM_w_io_v22_out)
  );
  ray_AABB_1 RAY_AABB ( // @[Top_1.scala 65:46]
    .clock(RAY_AABB_clock),
    .reset(RAY_AABB_reset),
    .io_ray_idir_x(RAY_AABB_io_ray_idir_x),
    .io_ray_idir_y(RAY_AABB_io_ray_idir_y),
    .io_ray_idir_z(RAY_AABB_io_ray_idir_z),
    .io_ray_ood_x(RAY_AABB_io_ray_ood_x),
    .io_ray_ood_y(RAY_AABB_io_ray_ood_y),
    .io_ray_ood_z(RAY_AABB_io_ray_ood_z),
    .io_ray_hitT(RAY_AABB_io_ray_hitT),
    .io_bvh_n0xy_x(RAY_AABB_io_bvh_n0xy_x),
    .io_bvh_n0xy_y(RAY_AABB_io_bvh_n0xy_y),
    .io_bvh_n0xy_z(RAY_AABB_io_bvh_n0xy_z),
    .io_bvh_n0xy_w(RAY_AABB_io_bvh_n0xy_w),
    .io_bvh_n1xy_x(RAY_AABB_io_bvh_n1xy_x),
    .io_bvh_n1xy_y(RAY_AABB_io_bvh_n1xy_y),
    .io_bvh_n1xy_z(RAY_AABB_io_bvh_n1xy_z),
    .io_bvh_n1xy_w(RAY_AABB_io_bvh_n1xy_w),
    .io_bvh_nz_x(RAY_AABB_io_bvh_nz_x),
    .io_bvh_nz_y(RAY_AABB_io_bvh_nz_y),
    .io_bvh_nz_z(RAY_AABB_io_bvh_nz_z),
    .io_bvh_nz_w(RAY_AABB_io_bvh_nz_w),
    .io_bvh_temp_x(RAY_AABB_io_bvh_temp_x),
    .io_bvh_temp_y(RAY_AABB_io_bvh_temp_y),
    .io_rayid(RAY_AABB_io_rayid),
    .io_valid_en(RAY_AABB_io_valid_en),
    .io_rayid_out(RAY_AABB_io_rayid_out),
    .io_nodeIdx_0(RAY_AABB_io_nodeIdx_0),
    .io_nodeIdx_1(RAY_AABB_io_nodeIdx_1),
    .io_nodeIdx_2(RAY_AABB_io_nodeIdx_2),
    .io_push(RAY_AABB_io_push),
    .io_pop(RAY_AABB_io_pop),
    .io_leaf(RAY_AABB_io_leaf),
    .io_back(RAY_AABB_io_back),
    .io_hitT_out(RAY_AABB_io_hitT_out),
    .io_valid_out(RAY_AABB_io_valid_out)
  );
  ray_AABB_1 RAY_AABB_2 ( // @[Top_1.scala 66:48]
    .clock(RAY_AABB_2_clock),
    .reset(RAY_AABB_2_reset),
    .io_ray_idir_x(RAY_AABB_2_io_ray_idir_x),
    .io_ray_idir_y(RAY_AABB_2_io_ray_idir_y),
    .io_ray_idir_z(RAY_AABB_2_io_ray_idir_z),
    .io_ray_ood_x(RAY_AABB_2_io_ray_ood_x),
    .io_ray_ood_y(RAY_AABB_2_io_ray_ood_y),
    .io_ray_ood_z(RAY_AABB_2_io_ray_ood_z),
    .io_ray_hitT(RAY_AABB_2_io_ray_hitT),
    .io_bvh_n0xy_x(RAY_AABB_2_io_bvh_n0xy_x),
    .io_bvh_n0xy_y(RAY_AABB_2_io_bvh_n0xy_y),
    .io_bvh_n0xy_z(RAY_AABB_2_io_bvh_n0xy_z),
    .io_bvh_n0xy_w(RAY_AABB_2_io_bvh_n0xy_w),
    .io_bvh_n1xy_x(RAY_AABB_2_io_bvh_n1xy_x),
    .io_bvh_n1xy_y(RAY_AABB_2_io_bvh_n1xy_y),
    .io_bvh_n1xy_z(RAY_AABB_2_io_bvh_n1xy_z),
    .io_bvh_n1xy_w(RAY_AABB_2_io_bvh_n1xy_w),
    .io_bvh_nz_x(RAY_AABB_2_io_bvh_nz_x),
    .io_bvh_nz_y(RAY_AABB_2_io_bvh_nz_y),
    .io_bvh_nz_z(RAY_AABB_2_io_bvh_nz_z),
    .io_bvh_nz_w(RAY_AABB_2_io_bvh_nz_w),
    .io_bvh_temp_x(RAY_AABB_2_io_bvh_temp_x),
    .io_bvh_temp_y(RAY_AABB_2_io_bvh_temp_y),
    .io_rayid(RAY_AABB_2_io_rayid),
    .io_valid_en(RAY_AABB_2_io_valid_en),
    .io_rayid_out(RAY_AABB_2_io_rayid_out),
    .io_nodeIdx_0(RAY_AABB_2_io_nodeIdx_0),
    .io_nodeIdx_1(RAY_AABB_2_io_nodeIdx_1),
    .io_nodeIdx_2(RAY_AABB_2_io_nodeIdx_2),
    .io_push(RAY_AABB_2_io_push),
    .io_pop(RAY_AABB_2_io_pop),
    .io_leaf(RAY_AABB_2_io_leaf),
    .io_back(RAY_AABB_2_io_back),
    .io_hitT_out(RAY_AABB_2_io_hitT_out),
    .io_valid_out(RAY_AABB_2_io_valid_out)
  );
  Arbitration_1 Arbitration_1 ( // @[Top_1.scala 67:50]
    .clock(Arbitration_1_clock),
    .reset(Arbitration_1_reset),
    .io_node_id_0(Arbitration_1_io_node_id_0),
    .io_ray_id_0(Arbitration_1_io_ray_id_0),
    .io_hit_0(Arbitration_1_io_hit_0),
    .io_valid_0(Arbitration_1_io_valid_0),
    .io_node_id_1(Arbitration_1_io_node_id_1),
    .io_ray_id_1(Arbitration_1_io_ray_id_1),
    .io_valid_1(Arbitration_1_io_valid_1),
    .io_ray_id_2(Arbitration_1_io_ray_id_2),
    .io_valid_2(Arbitration_1_io_valid_2),
    .io_node_id_out(Arbitration_1_io_node_id_out),
    .io_ray_id_out(Arbitration_1_io_ray_id_out),
    .io_hit_out(Arbitration_1_io_hit_out),
    .io_valid_out(Arbitration_1_io_valid_out)
  );
  Arbitration_1 Arbitration_1_2 ( // @[Top_1.scala 68:47]
    .clock(Arbitration_1_2_clock),
    .reset(Arbitration_1_2_reset),
    .io_node_id_0(Arbitration_1_2_io_node_id_0),
    .io_ray_id_0(Arbitration_1_2_io_ray_id_0),
    .io_hit_0(Arbitration_1_2_io_hit_0),
    .io_valid_0(Arbitration_1_2_io_valid_0),
    .io_node_id_1(Arbitration_1_2_io_node_id_1),
    .io_ray_id_1(Arbitration_1_2_io_ray_id_1),
    .io_valid_1(Arbitration_1_2_io_valid_1),
    .io_ray_id_2(Arbitration_1_2_io_ray_id_2),
    .io_valid_2(Arbitration_1_2_io_valid_2),
    .io_node_id_out(Arbitration_1_2_io_node_id_out),
    .io_ray_id_out(Arbitration_1_2_io_ray_id_out),
    .io_hit_out(Arbitration_1_2_io_hit_out),
    .io_valid_out(Arbitration_1_2_io_valid_out)
  );
  Arbitration_2_1 Arbitration_2 ( // @[Top_1.scala 70:45]
    .clock(Arbitration_2_clock),
    .reset(Arbitration_2_reset),
    .io_ray_id_2_0(Arbitration_2_io_ray_id_2_0),
    .io_hit_2_0(Arbitration_2_io_hit_2_0),
    .io_valid_2_0(Arbitration_2_io_valid_2_0),
    .io_ray_id_2_1(Arbitration_2_io_ray_id_2_1),
    .io_hit_2_1(Arbitration_2_io_hit_2_1),
    .io_valid_2_1(Arbitration_2_io_valid_2_1),
    .io_ray_id_2_2(Arbitration_2_io_ray_id_2_2),
    .io_hit_2_2(Arbitration_2_io_hit_2_2),
    .io_valid_2_2(Arbitration_2_io_valid_2_2),
    .io_ray_id_2_3(Arbitration_2_io_ray_id_2_3),
    .io_hit_2_3(Arbitration_2_io_hit_2_3),
    .io_valid_2_3(Arbitration_2_io_valid_2_3),
    .io_ray_id_out(Arbitration_2_io_ray_id_out),
    .io_hit_out(Arbitration_2_io_hit_out),
    .io_valid_out(Arbitration_2_io_valid_out)
  );
  Arbitration_2_1 Arbitration_2_2 ( // @[Top_1.scala 71:42]
    .clock(Arbitration_2_2_clock),
    .reset(Arbitration_2_2_reset),
    .io_ray_id_2_0(Arbitration_2_2_io_ray_id_2_0),
    .io_hit_2_0(Arbitration_2_2_io_hit_2_0),
    .io_valid_2_0(Arbitration_2_2_io_valid_2_0),
    .io_ray_id_2_1(Arbitration_2_2_io_ray_id_2_1),
    .io_hit_2_1(Arbitration_2_2_io_hit_2_1),
    .io_valid_2_1(Arbitration_2_2_io_valid_2_1),
    .io_ray_id_2_2(Arbitration_2_2_io_ray_id_2_2),
    .io_hit_2_2(Arbitration_2_2_io_hit_2_2),
    .io_valid_2_2(Arbitration_2_2_io_valid_2_2),
    .io_ray_id_2_3(Arbitration_2_2_io_ray_id_2_3),
    .io_hit_2_3(Arbitration_2_2_io_hit_2_3),
    .io_valid_2_3(Arbitration_2_2_io_valid_2_3),
    .io_ray_id_out(Arbitration_2_2_io_ray_id_out),
    .io_hit_out(Arbitration_2_2_io_hit_out),
    .io_valid_out(Arbitration_2_2_io_valid_out)
  );
  Arbitration_3 Arbitration_3 ( // @[Top_1.scala 72:45]
    .clock(Arbitration_3_clock),
    .reset(Arbitration_3_reset),
    .io_node_id_3_0(Arbitration_3_io_node_id_3_0),
    .io_ray_id_3_0(Arbitration_3_io_ray_id_3_0),
    .io_hit_3_0(Arbitration_3_io_hit_3_0),
    .io_valid_3_0(Arbitration_3_io_valid_3_0),
    .io_node_id_3_1(Arbitration_3_io_node_id_3_1),
    .io_ray_id_3_1(Arbitration_3_io_ray_id_3_1),
    .io_hit_3_1(Arbitration_3_io_hit_3_1),
    .io_valid_3_1(Arbitration_3_io_valid_3_1),
    .io_node_id_3_2(Arbitration_3_io_node_id_3_2),
    .io_ray_id_3_2(Arbitration_3_io_ray_id_3_2),
    .io_hit_3_2(Arbitration_3_io_hit_3_2),
    .io_valid_3_2(Arbitration_3_io_valid_3_2),
    .io_node_id_3_3(Arbitration_3_io_node_id_3_3),
    .io_ray_id_3_3(Arbitration_3_io_ray_id_3_3),
    .io_hit_3_3(Arbitration_3_io_hit_3_3),
    .io_valid_3_3(Arbitration_3_io_valid_3_3),
    .io_node_id_3_4(Arbitration_3_io_node_id_3_4),
    .io_ray_id_3_4(Arbitration_3_io_ray_id_3_4),
    .io_hit_3_4(Arbitration_3_io_hit_3_4),
    .io_valid_3_4(Arbitration_3_io_valid_3_4),
    .io_node_id_out(Arbitration_3_io_node_id_out),
    .io_ray_id_out(Arbitration_3_io_ray_id_out),
    .io_hit_out(Arbitration_3_io_hit_out),
    .io_valid_out(Arbitration_3_io_valid_out)
  );
  Arbitration_3 Arbitration_3_2 ( // @[Top_1.scala 73:42]
    .clock(Arbitration_3_2_clock),
    .reset(Arbitration_3_2_reset),
    .io_node_id_3_0(Arbitration_3_2_io_node_id_3_0),
    .io_ray_id_3_0(Arbitration_3_2_io_ray_id_3_0),
    .io_hit_3_0(Arbitration_3_2_io_hit_3_0),
    .io_valid_3_0(Arbitration_3_2_io_valid_3_0),
    .io_node_id_3_1(Arbitration_3_2_io_node_id_3_1),
    .io_ray_id_3_1(Arbitration_3_2_io_ray_id_3_1),
    .io_hit_3_1(Arbitration_3_2_io_hit_3_1),
    .io_valid_3_1(Arbitration_3_2_io_valid_3_1),
    .io_node_id_3_2(Arbitration_3_2_io_node_id_3_2),
    .io_ray_id_3_2(Arbitration_3_2_io_ray_id_3_2),
    .io_hit_3_2(Arbitration_3_2_io_hit_3_2),
    .io_valid_3_2(Arbitration_3_2_io_valid_3_2),
    .io_node_id_3_3(Arbitration_3_2_io_node_id_3_3),
    .io_ray_id_3_3(Arbitration_3_2_io_ray_id_3_3),
    .io_hit_3_3(Arbitration_3_2_io_hit_3_3),
    .io_valid_3_3(Arbitration_3_2_io_valid_3_3),
    .io_node_id_3_4(Arbitration_3_2_io_node_id_3_4),
    .io_ray_id_3_4(Arbitration_3_2_io_ray_id_3_4),
    .io_hit_3_4(Arbitration_3_2_io_hit_3_4),
    .io_valid_3_4(Arbitration_3_2_io_valid_3_4),
    .io_node_id_out(Arbitration_3_2_io_node_id_out),
    .io_ray_id_out(Arbitration_3_2_io_ray_id_out),
    .io_hit_out(Arbitration_3_2_io_hit_out),
    .io_valid_out(Arbitration_3_2_io_valid_out)
  );
  Arbitration_4 Arbitration_4 ( // @[Top_1.scala 74:45]
    .clock(Arbitration_4_clock),
    .reset(Arbitration_4_reset),
    .io_node_id_4_0(Arbitration_4_io_node_id_4_0),
    .io_ray_id_4_0(Arbitration_4_io_ray_id_4_0),
    .io_hit_4_0(Arbitration_4_io_hit_4_0),
    .io_valid_4_0(Arbitration_4_io_valid_4_0),
    .io_node_id_4_1(Arbitration_4_io_node_id_4_1),
    .io_ray_id_4_1(Arbitration_4_io_ray_id_4_1),
    .io_hit_4_1(Arbitration_4_io_hit_4_1),
    .io_valid_4_1(Arbitration_4_io_valid_4_1),
    .io_node_id_out(Arbitration_4_io_node_id_out),
    .io_ray_id_out(Arbitration_4_io_ray_id_out),
    .io_hit_out(Arbitration_4_io_hit_out),
    .io_RAY_AABB_out(Arbitration_4_io_RAY_AABB_out),
    .io_RAY_AABB_2_out(Arbitration_4_io_RAY_AABB_2_out),
    .io_valid_out(Arbitration_4_io_valid_out)
  );
  Stackmanage Stack_manage ( // @[Top_1.scala 75:41]
    .clock(Stack_manage_clock),
    .reset(Stack_manage_reset),
    .io_push(Stack_manage_io_push),
    .io_push_en(Stack_manage_io_push_en),
    .io_pop(Stack_manage_io_pop),
    .io_pop_en(Stack_manage_io_pop_en),
    .io_ray_id_push(Stack_manage_io_ray_id_push),
    .io_ray_id_pop(Stack_manage_io_ray_id_pop),
    .io_node_id_push_in(Stack_manage_io_node_id_push_in),
    .io_hitT_in(Stack_manage_io_hitT_in),
    .io_hitT_out(Stack_manage_io_hitT_out),
    .io_node_id_out(Stack_manage_io_node_id_out),
    .io_ray_id_out(Stack_manage_io_ray_id_out),
    .io_pop_valid(Stack_manage_io_pop_valid),
    .io_Dis_en(Stack_manage_io_Dis_en),
    .io_Finish(Stack_manage_io_Finish)
  );
  Stackmanage Stack_manage_2 ( // @[Top_1.scala 76:38]
    .clock(Stack_manage_2_clock),
    .reset(Stack_manage_2_reset),
    .io_push(Stack_manage_2_io_push),
    .io_push_en(Stack_manage_2_io_push_en),
    .io_pop(Stack_manage_2_io_pop),
    .io_pop_en(Stack_manage_2_io_pop_en),
    .io_ray_id_push(Stack_manage_2_io_ray_id_push),
    .io_ray_id_pop(Stack_manage_2_io_ray_id_pop),
    .io_node_id_push_in(Stack_manage_2_io_node_id_push_in),
    .io_hitT_in(Stack_manage_2_io_hitT_in),
    .io_hitT_out(Stack_manage_2_io_hitT_out),
    .io_node_id_out(Stack_manage_2_io_node_id_out),
    .io_ray_id_out(Stack_manage_2_io_ray_id_out),
    .io_pop_valid(Stack_manage_2_io_pop_valid),
    .io_Dis_en(Stack_manage_2_io_Dis_en),
    .io_Finish(Stack_manage_2_io_Finish)
  );
  Triangle Triangle ( // @[Top_1.scala 77:51]
    .clock(Triangle_clock),
    .reset(Triangle_reset),
    .io_To_IST0_enable(Triangle_io_To_IST0_enable),
    .io_nodeid_leaf(Triangle_io_nodeid_leaf),
    .io_rayid_leaf(Triangle_io_rayid_leaf),
    .io_hiT_in(Triangle_io_hiT_in),
    .io_v00_in_x(Triangle_io_v00_in_x),
    .io_v00_in_y(Triangle_io_v00_in_y),
    .io_v00_in_z(Triangle_io_v00_in_z),
    .io_v00_in_w(Triangle_io_v00_in_w),
    .io_v11_in_x(Triangle_io_v11_in_x),
    .io_v11_in_y(Triangle_io_v11_in_y),
    .io_v11_in_z(Triangle_io_v11_in_z),
    .io_v11_in_w(Triangle_io_v11_in_w),
    .io_v22_in_x(Triangle_io_v22_in_x),
    .io_v22_in_y(Triangle_io_v22_in_y),
    .io_v22_in_z(Triangle_io_v22_in_z),
    .io_v22_in_w(Triangle_io_v22_in_w),
    .io_ray_o_in_x(Triangle_io_ray_o_in_x),
    .io_ray_o_in_y(Triangle_io_ray_o_in_y),
    .io_ray_o_in_z(Triangle_io_ray_o_in_z),
    .io_ray_d_in_x(Triangle_io_ray_d_in_x),
    .io_ray_d_in_y(Triangle_io_ray_d_in_y),
    .io_ray_d_in_z(Triangle_io_ray_d_in_z),
    .io_break_in(Triangle_io_break_in),
    .io_RAY_AABB_1(Triangle_io_RAY_AABB_1),
    .io_RAY_AABB_2(Triangle_io_RAY_AABB_2),
    .io_pop_1(Triangle_io_pop_1),
    .io_break_1(Triangle_io_break_1),
    .io_pop_2(Triangle_io_pop_2),
    .io_break_2(Triangle_io_break_2),
    .io_pop_3(Triangle_io_pop_3),
    .io_break_3(Triangle_io_break_3),
    .io_hiT_out_1(Triangle_io_hiT_out_1),
    .io_hiT_out_2(Triangle_io_hiT_out_2),
    .io_hiT_out_3(Triangle_io_hiT_out_3),
    .io_hitT_en(Triangle_io_hitT_en),
    .io_hitIndex(Triangle_io_hitIndex),
    .io_node_id_out_1(Triangle_io_node_id_out_1),
    .io_node_id_out_2(Triangle_io_node_id_out_2),
    .io_node_id_out_3(Triangle_io_node_id_out_3),
    .io_ray_id_ist1(Triangle_io_ray_id_ist1),
    .io_ray_id_ist2(Triangle_io_ray_id_ist2),
    .io_ray_id_ist3(Triangle_io_ray_id_ist3),
    .io_counter_fdiv(Triangle_io_counter_fdiv),
    .io_RAY_AABB_1_out_IST1(Triangle_io_RAY_AABB_1_out_IST1),
    .io_RAY_AABB_2_out_IST1(Triangle_io_RAY_AABB_2_out_IST1),
    .io_RAY_AABB_1_out_IST2(Triangle_io_RAY_AABB_1_out_IST2),
    .io_RAY_AABB_2_out_IST2(Triangle_io_RAY_AABB_2_out_IST2),
    .io_RAY_AABB_1_out_IST3(Triangle_io_RAY_AABB_1_out_IST3),
    .io_RAY_AABB_2_out_IST3(Triangle_io_RAY_AABB_2_out_IST3)
  );
  assign io_hitT = Triangle_io_hitT_en ? Triangle_io_hiT_out_3 : 32'h0; // @[Top_1.scala 764:30 Top_1.scala 765:70 Top_1.scala 769:70]
  assign io_hitIndex = Triangle_io_hitT_en ? $signed(Triangle_io_hitIndex) : $signed(32'sh0); // @[Top_1.scala 764:30 Top_1.scala 766:65 Top_1.scala 770:65]
  assign io_rtp_finish = Ray_Dispatch_io_ray_finish & Stack_manage_io_Finish; // @[Top_1.scala 107:87]
  assign io_ray_id_triangle = Triangle_io_hitT_en ? Triangle_io_ray_id_ist3 : 32'h0; // @[Top_1.scala 764:30 Top_1.scala 767:57 Top_1.scala 771:57]
  assign io_counter_fdiv = Triangle_io_counter_fdiv; // @[Top_1.scala 759:57]
  assign io_TRV_1_valid = TRV_1; // @[Top_1.scala 250:61]
  assign io_TRV_2_valid = TRV_2; // @[Top_1.scala 396:66]
  assign io_IST_1_valid = IST_1; // @[Top_1.scala 753:59]
  assign io_clock_count = clock_counter; // @[Top_1.scala 81:37]
  assign Ray_Dispatch_clock = clock;
  assign Ray_Dispatch_reset = reset;
  assign Ray_Dispatch_io_dispatch = Stack_manage_io_Dis_en; // @[Top_1.scala 84:53]
  assign Ray_Dispatch_io_dispatch_2 = Stack_manage_2_io_Dis_en; // @[Top_1.scala 85:50]
  assign Ray_origx_clock = clock;
  assign Ray_origx_io_Ray_id = Arbitration_4_io_ray_id_out; // @[Top_1.scala 673:37 Top_1.scala 679:54]
  assign Ray_origx_io_Ray_id_2 = 32'h0;
  assign Ray_origy_clock = clock;
  assign Ray_origy_io_Ray_id = Arbitration_4_io_ray_id_out; // @[Top_1.scala 673:37 Top_1.scala 679:54]
  assign Ray_origy_io_Ray_id_2 = 32'h0;
  assign Ray_origz_clock = clock;
  assign Ray_origz_io_Ray_id = Arbitration_4_io_ray_id_out; // @[Top_1.scala 673:37 Top_1.scala 679:54]
  assign Ray_origz_io_Ray_id_2 = 32'h0;
  assign Ray_dirx_clock = clock;
  assign Ray_dirx_io_Ray_id = Arbitration_4_io_ray_id_out; // @[Top_1.scala 673:37 Top_1.scala 679:54]
  assign Ray_dirx_io_Ray_id_2 = 32'h0;
  assign Ray_diry_clock = clock;
  assign Ray_diry_io_Ray_id = Arbitration_4_io_ray_id_out; // @[Top_1.scala 673:37 Top_1.scala 679:54]
  assign Ray_diry_io_Ray_id_2 = 32'h0;
  assign Ray_dirz_clock = clock;
  assign Ray_dirz_io_Ray_id = Arbitration_4_io_ray_id_out; // @[Top_1.scala 673:37 Top_1.scala 679:54]
  assign Ray_dirz_io_Ray_id_2 = 32'h0;
  assign Ray_hitT_clock = clock;
  assign Ray_hitT_io_Ray_id = Arbitration_1_io_hit_out; // @[Top_1.scala 159:76 Top_1.scala 182:53]
  assign Ray_hitT_io_Ray_id_2 = Arbitration_1_2_io_ray_id_out; // @[Top_1.scala 296:80 Top_1.scala 300:54]
  assign Ray_idirx_clock = clock;
  assign Ray_idirx_io_Ray_id = Arbitration_1_io_valid_out & Arbitration_1_io_hit_out != 32'h0 ?
    Arbitration_1_io_ray_id_out : _GEN_13; // @[Top_1.scala 134:70 Top_1.scala 136:51]
  assign Ray_idirx_io_Ray_id_2 = Arbitration_1_2_io_valid_out & Arbitration_1_2_io_hit_out != 32'h0 ?
    Arbitration_1_2_io_ray_id_out : _GEN_81; // @[Top_1.scala 269:74 Top_1.scala 273:55]
  assign Ray_idiry_clock = clock;
  assign Ray_idiry_io_Ray_id = Arbitration_1_io_valid_out & Arbitration_1_io_hit_out != 32'h0 ?
    Arbitration_1_io_ray_id_out : _GEN_13; // @[Top_1.scala 134:70 Top_1.scala 136:51]
  assign Ray_idiry_io_Ray_id_2 = Arbitration_1_2_io_valid_out & Arbitration_1_2_io_hit_out != 32'h0 ?
    Arbitration_1_2_io_ray_id_out : _GEN_81; // @[Top_1.scala 269:74 Top_1.scala 273:55]
  assign Ray_idirz_clock = clock;
  assign Ray_idirz_io_Ray_id = Arbitration_1_io_valid_out & Arbitration_1_io_hit_out != 32'h0 ?
    Arbitration_1_io_ray_id_out : _GEN_13; // @[Top_1.scala 134:70 Top_1.scala 136:51]
  assign Ray_idirz_io_Ray_id_2 = Arbitration_1_2_io_valid_out & Arbitration_1_2_io_hit_out != 32'h0 ?
    Arbitration_1_2_io_ray_id_out : _GEN_81; // @[Top_1.scala 269:74 Top_1.scala 273:55]
  assign Ray_oodx_clock = clock;
  assign Ray_oodx_io_Ray_id = Arbitration_1_io_valid_out & Arbitration_1_io_hit_out != 32'h0 ?
    Arbitration_1_io_ray_id_out : _GEN_13; // @[Top_1.scala 134:70 Top_1.scala 136:51]
  assign Ray_oodx_io_Ray_id_2 = Arbitration_1_2_io_valid_out & Arbitration_1_2_io_hit_out != 32'h0 ?
    Arbitration_1_2_io_ray_id_out : _GEN_81; // @[Top_1.scala 269:74 Top_1.scala 273:55]
  assign Ray_oody_clock = clock;
  assign Ray_oody_io_Ray_id = Arbitration_1_io_valid_out & Arbitration_1_io_hit_out != 32'h0 ?
    Arbitration_1_io_ray_id_out : _GEN_13; // @[Top_1.scala 134:70 Top_1.scala 136:51]
  assign Ray_oody_io_Ray_id_2 = Arbitration_1_2_io_valid_out & Arbitration_1_2_io_hit_out != 32'h0 ?
    Arbitration_1_2_io_ray_id_out : _GEN_81; // @[Top_1.scala 269:74 Top_1.scala 273:55]
  assign Ray_oodz_clock = clock;
  assign Ray_oodz_io_Ray_id = Arbitration_1_io_valid_out & Arbitration_1_io_hit_out != 32'h0 ?
    Arbitration_1_io_ray_id_out : _GEN_13; // @[Top_1.scala 134:70 Top_1.scala 136:51]
  assign Ray_oodz_io_Ray_id_2 = Arbitration_1_2_io_valid_out & Arbitration_1_2_io_hit_out != 32'h0 ?
    Arbitration_1_2_io_ray_id_out : _GEN_81; // @[Top_1.scala 269:74 Top_1.scala 273:55]
  assign BVH_RAM_0_x_clock = clock;
  assign BVH_RAM_0_x_io_BVH_id = _GEN_34[31:0];
  assign BVH_RAM_0_x_io_BVH_id_2 = _GEN_101[31:0];
  assign BVH_RAM_0_y_clock = clock;
  assign BVH_RAM_0_y_io_BVH_id = _GEN_34[31:0];
  assign BVH_RAM_0_y_io_BVH_id_2 = _GEN_101[31:0];
  assign BVH_RAM_0_z_clock = clock;
  assign BVH_RAM_0_z_io_BVH_id = _GEN_34[31:0];
  assign BVH_RAM_0_z_io_BVH_id_2 = _GEN_101[31:0];
  assign BVH_RAM_0_w_clock = clock;
  assign BVH_RAM_0_w_io_BVH_id = _GEN_34[31:0];
  assign BVH_RAM_0_w_io_BVH_id_2 = _GEN_101[31:0];
  assign BVH_RAM_1_x_clock = clock;
  assign BVH_RAM_1_x_io_BVH_id = _GEN_34[31:0];
  assign BVH_RAM_1_x_io_BVH_id_2 = _GEN_101[31:0];
  assign BVH_RAM_1_y_clock = clock;
  assign BVH_RAM_1_y_io_BVH_id = _GEN_34[31:0];
  assign BVH_RAM_1_y_io_BVH_id_2 = _GEN_101[31:0];
  assign BVH_RAM_1_z_clock = clock;
  assign BVH_RAM_1_z_io_BVH_id = _GEN_34[31:0];
  assign BVH_RAM_1_z_io_BVH_id_2 = _GEN_101[31:0];
  assign BVH_RAM_1_w_clock = clock;
  assign BVH_RAM_1_w_io_BVH_id = _GEN_34[31:0];
  assign BVH_RAM_1_w_io_BVH_id_2 = _GEN_101[31:0];
  assign BVH_RAM_z_x_clock = clock;
  assign BVH_RAM_z_x_io_BVH_id = _GEN_34[31:0];
  assign BVH_RAM_z_x_io_BVH_id_2 = _GEN_101[31:0];
  assign BVH_RAM_z_y_clock = clock;
  assign BVH_RAM_z_y_io_BVH_id = _GEN_34[31:0];
  assign BVH_RAM_z_y_io_BVH_id_2 = _GEN_101[31:0];
  assign BVH_RAM_z_z_clock = clock;
  assign BVH_RAM_z_z_io_BVH_id = _GEN_34[31:0];
  assign BVH_RAM_z_z_io_BVH_id_2 = _GEN_101[31:0];
  assign BVH_RAM_z_w_clock = clock;
  assign BVH_RAM_z_w_io_BVH_id = _GEN_34[31:0];
  assign BVH_RAM_z_w_io_BVH_id_2 = _GEN_101[31:0];
  assign BVH_RAM_tmp_x_clock = clock;
  assign BVH_RAM_tmp_x_io_BVH_id = _GEN_34[31:0];
  assign BVH_RAM_tmp_x_io_BVH_id_2 = _GEN_101[31:0];
  assign BVH_RAM_tmp_y_clock = clock;
  assign BVH_RAM_tmp_y_io_BVH_id = _GEN_34[31:0];
  assign BVH_RAM_tmp_y_io_BVH_id_2 = _GEN_101[31:0];
  assign TRI_RAM_x_clock = clock;
  assign TRI_RAM_x_io_Triangle_id = Arbitration_4_io_node_id_out; // @[Top_1.scala 673:37 Top_1.scala 675:47]
  assign TRI_RAM_y_clock = clock;
  assign TRI_RAM_y_io_Triangle_id = Arbitration_4_io_node_id_out; // @[Top_1.scala 673:37 Top_1.scala 675:47]
  assign TRI_RAM_z_clock = clock;
  assign TRI_RAM_z_io_Triangle_id = Arbitration_4_io_node_id_out; // @[Top_1.scala 673:37 Top_1.scala 675:47]
  assign TRI_RAM_w_clock = clock;
  assign TRI_RAM_w_io_Triangle_id = Arbitration_4_io_node_id_out; // @[Top_1.scala 673:37 Top_1.scala 675:47]
  assign RAY_AABB_clock = clock;
  assign RAY_AABB_reset = reset;
  assign RAY_AABB_io_ray_idir_x = memory_valid ? Ray_idirx_io_Ray_out : 32'h0; // @[Top_1.scala 190:29 Top_1.scala 191:53 Top_1.scala 224:53]
  assign RAY_AABB_io_ray_idir_y = memory_valid ? Ray_idiry_io_Ray_out : 32'h0; // @[Top_1.scala 190:29 Top_1.scala 192:53 Top_1.scala 225:53]
  assign RAY_AABB_io_ray_idir_z = memory_valid ? Ray_idirz_io_Ray_out : 32'h0; // @[Top_1.scala 190:29 Top_1.scala 193:53 Top_1.scala 226:53]
  assign RAY_AABB_io_ray_ood_x = memory_valid ? Ray_oodx_io_Ray_out : 32'h0; // @[Top_1.scala 190:29 Top_1.scala 194:51 Top_1.scala 227:51]
  assign RAY_AABB_io_ray_ood_y = memory_valid ? Ray_oody_io_Ray_out : 32'h0; // @[Top_1.scala 190:29 Top_1.scala 195:51 Top_1.scala 228:51]
  assign RAY_AABB_io_ray_ood_z = memory_valid ? Ray_oodz_io_Ray_out : 32'h0; // @[Top_1.scala 190:29 Top_1.scala 196:51 Top_1.scala 229:51]
  assign RAY_AABB_io_ray_hitT = memory_valid ? _GEN_51 : 32'h0; // @[Top_1.scala 190:29 Top_1.scala 230:53]
  assign RAY_AABB_io_bvh_n0xy_x = memory_valid ? BVH_RAM_0_x_io_BVH_out : 32'h0; // @[Top_1.scala 190:29 Top_1.scala 203:49 Top_1.scala 232:49]
  assign RAY_AABB_io_bvh_n0xy_y = memory_valid ? BVH_RAM_0_y_io_BVH_out : 32'h0; // @[Top_1.scala 190:29 Top_1.scala 204:49 Top_1.scala 233:49]
  assign RAY_AABB_io_bvh_n0xy_z = memory_valid ? BVH_RAM_0_z_io_BVH_out : 32'h0; // @[Top_1.scala 190:29 Top_1.scala 205:49 Top_1.scala 234:49]
  assign RAY_AABB_io_bvh_n0xy_w = memory_valid ? BVH_RAM_0_w_io_BVH_out : 32'h0; // @[Top_1.scala 190:29 Top_1.scala 206:48 Top_1.scala 235:48]
  assign RAY_AABB_io_bvh_n1xy_x = memory_valid ? BVH_RAM_1_x_io_BVH_out : 32'h0; // @[Top_1.scala 190:29 Top_1.scala 208:49 Top_1.scala 236:49]
  assign RAY_AABB_io_bvh_n1xy_y = memory_valid ? BVH_RAM_1_y_io_BVH_out : 32'h0; // @[Top_1.scala 190:29 Top_1.scala 209:49 Top_1.scala 237:49]
  assign RAY_AABB_io_bvh_n1xy_z = memory_valid ? BVH_RAM_1_z_io_BVH_out : 32'h0; // @[Top_1.scala 190:29 Top_1.scala 210:49 Top_1.scala 238:49]
  assign RAY_AABB_io_bvh_n1xy_w = memory_valid ? BVH_RAM_1_w_io_BVH_out : 32'h0; // @[Top_1.scala 190:29 Top_1.scala 211:48 Top_1.scala 239:48]
  assign RAY_AABB_io_bvh_nz_x = memory_valid ? BVH_RAM_z_x_io_BVH_out : 32'h0; // @[Top_1.scala 190:29 Top_1.scala 213:51 Top_1.scala 240:51]
  assign RAY_AABB_io_bvh_nz_y = memory_valid ? BVH_RAM_z_y_io_BVH_out : 32'h0; // @[Top_1.scala 190:29 Top_1.scala 214:51 Top_1.scala 241:51]
  assign RAY_AABB_io_bvh_nz_z = memory_valid ? BVH_RAM_z_z_io_BVH_out : 32'h0; // @[Top_1.scala 190:29 Top_1.scala 215:51 Top_1.scala 242:51]
  assign RAY_AABB_io_bvh_nz_w = memory_valid ? BVH_RAM_z_w_io_BVH_out : 32'h0; // @[Top_1.scala 190:29 Top_1.scala 216:50 Top_1.scala 243:49]
  assign RAY_AABB_io_bvh_temp_x = memory_valid ? $signed(BVH_RAM_tmp_x_io_BVH_out) : $signed(32'sh0); // @[Top_1.scala 190:29 Top_1.scala 218:48 Top_1.scala 244:48]
  assign RAY_AABB_io_bvh_temp_y = memory_valid ? $signed(BVH_RAM_tmp_y_io_BVH_out) : $signed(32'sh0); // @[Top_1.scala 190:29 Top_1.scala 219:48 Top_1.scala 245:48]
  assign RAY_AABB_io_rayid = memory_valid ? ray_id_temp : 32'h0; // @[Top_1.scala 190:29 Top_1.scala 220:57 Top_1.scala 246:57]
  assign RAY_AABB_io_valid_en = memory_valid; // @[Top_1.scala 190:29 Top_1.scala 221:53 Top_1.scala 247:53]
  assign RAY_AABB_2_clock = clock;
  assign RAY_AABB_2_reset = reset;
  assign RAY_AABB_2_io_ray_idir_x = memory_valid_2 ? Ray_idirx_io_Ray_out_2 : 32'h0; // @[Top_1.scala 329:31 Top_1.scala 330:55 Top_1.scala 360:55]
  assign RAY_AABB_2_io_ray_idir_y = memory_valid_2 ? Ray_idiry_io_Ray_out_2 : 32'h0; // @[Top_1.scala 329:31 Top_1.scala 331:55 Top_1.scala 361:55]
  assign RAY_AABB_2_io_ray_idir_z = memory_valid_2 ? Ray_idirz_io_Ray_out_2 : 32'h0; // @[Top_1.scala 329:31 Top_1.scala 332:55 Top_1.scala 362:55]
  assign RAY_AABB_2_io_ray_ood_x = memory_valid_2 ? Ray_oodx_io_Ray_out_2 : 32'h0; // @[Top_1.scala 329:31 Top_1.scala 333:53 Top_1.scala 363:53]
  assign RAY_AABB_2_io_ray_ood_y = memory_valid_2 ? Ray_oody_io_Ray_out_2 : 32'h0; // @[Top_1.scala 329:31 Top_1.scala 334:53 Top_1.scala 364:53]
  assign RAY_AABB_2_io_ray_ood_z = memory_valid_2 ? Ray_oodz_io_Ray_out_2 : 32'h0; // @[Top_1.scala 329:31 Top_1.scala 335:53 Top_1.scala 365:53]
  assign RAY_AABB_2_io_ray_hitT = memory_valid_2 ? _GEN_118 : 32'h0; // @[Top_1.scala 329:31 Top_1.scala 366:55]
  assign RAY_AABB_2_io_bvh_n0xy_x = memory_valid_2 ? BVH_RAM_0_x_io_BVH_out_2 : 32'h0; // @[Top_1.scala 329:31 Top_1.scala 342:51 Top_1.scala 368:51]
  assign RAY_AABB_2_io_bvh_n0xy_y = memory_valid_2 ? BVH_RAM_0_y_io_BVH_out_2 : 32'h0; // @[Top_1.scala 329:31 Top_1.scala 343:51 Top_1.scala 369:51]
  assign RAY_AABB_2_io_bvh_n0xy_z = memory_valid_2 ? BVH_RAM_0_z_io_BVH_out_2 : 32'h0; // @[Top_1.scala 329:31 Top_1.scala 344:51 Top_1.scala 370:51]
  assign RAY_AABB_2_io_bvh_n0xy_w = memory_valid_2 ? BVH_RAM_0_w_io_BVH_out_2 : 32'h0; // @[Top_1.scala 329:31 Top_1.scala 345:50 Top_1.scala 371:50]
  assign RAY_AABB_2_io_bvh_n1xy_x = memory_valid_2 ? BVH_RAM_1_x_io_BVH_out_2 : 32'h0; // @[Top_1.scala 329:31 Top_1.scala 346:51 Top_1.scala 372:51]
  assign RAY_AABB_2_io_bvh_n1xy_y = memory_valid_2 ? BVH_RAM_1_y_io_BVH_out_2 : 32'h0; // @[Top_1.scala 329:31 Top_1.scala 347:51 Top_1.scala 373:51]
  assign RAY_AABB_2_io_bvh_n1xy_z = memory_valid_2 ? BVH_RAM_1_z_io_BVH_out_2 : 32'h0; // @[Top_1.scala 329:31 Top_1.scala 348:51 Top_1.scala 374:51]
  assign RAY_AABB_2_io_bvh_n1xy_w = memory_valid_2 ? BVH_RAM_1_w_io_BVH_out_2 : 32'h0; // @[Top_1.scala 329:31 Top_1.scala 349:50 Top_1.scala 375:50]
  assign RAY_AABB_2_io_bvh_nz_x = memory_valid_2 ? BVH_RAM_z_x_io_BVH_out_2 : 32'h0; // @[Top_1.scala 329:31 Top_1.scala 350:53 Top_1.scala 376:53]
  assign RAY_AABB_2_io_bvh_nz_y = memory_valid_2 ? BVH_RAM_z_y_io_BVH_out_2 : 32'h0; // @[Top_1.scala 329:31 Top_1.scala 351:53 Top_1.scala 377:53]
  assign RAY_AABB_2_io_bvh_nz_z = memory_valid_2 ? BVH_RAM_z_z_io_BVH_out_2 : 32'h0; // @[Top_1.scala 329:31 Top_1.scala 352:53 Top_1.scala 378:53]
  assign RAY_AABB_2_io_bvh_nz_w = memory_valid_2 ? BVH_RAM_z_w_io_BVH_out_2 : 32'h0; // @[Top_1.scala 329:31 Top_1.scala 353:52 Top_1.scala 379:51]
  assign RAY_AABB_2_io_bvh_temp_x = memory_valid_2 ? $signed(BVH_RAM_tmp_x_io_BVH_out_2) : $signed(32'sh0); // @[Top_1.scala 329:31 Top_1.scala 354:50 Top_1.scala 381:50]
  assign RAY_AABB_2_io_bvh_temp_y = memory_valid_2 ? $signed(BVH_RAM_tmp_y_io_BVH_out_2) : $signed(32'sh0); // @[Top_1.scala 329:31 Top_1.scala 355:50 Top_1.scala 382:50]
  assign RAY_AABB_2_io_rayid = memory_valid_2 ? ray_id_temp_2 : 32'h0; // @[Top_1.scala 329:31 Top_1.scala 356:59 Top_1.scala 383:59]
  assign RAY_AABB_2_io_valid_en = memory_valid_2; // @[Top_1.scala 329:31 Top_1.scala 357:55 Top_1.scala 384:55]
  assign Arbitration_1_clock = clock;
  assign Arbitration_1_reset = reset;
  assign Arbitration_1_io_node_id_0 = _T_96 & Stack_manage_io_pop_valid ? $signed(Stack_manage_io_node_id_out) :
    $signed(32'sh0); // @[Top_1.scala 451:81 Top_1.scala 452:47]
  assign Arbitration_1_io_ray_id_0 = {{32'd0}, _GEN_168}; // @[Top_1.scala 451:81 Top_1.scala 453:50]
  assign Arbitration_1_io_hit_0 = _T_96 & Stack_manage_io_pop_valid ? Stack_manage_io_hitT_out : 32'h0; // @[Top_1.scala 451:81 Top_1.scala 454:54]
  assign Arbitration_1_io_valid_0 = _T_96 & Stack_manage_io_pop_valid; // @[Top_1.scala 451:53]
  assign Arbitration_1_io_node_id_1 = RAY_AABB_io_back & RAY_AABB_io_valid_out ? $signed(RAY_AABB_io_nodeIdx_1) :
    $signed(32'sh0); // @[Top_1.scala 110:50 Top_1.scala 111:37 Top_1.scala 115:37]
  assign Arbitration_1_io_ray_id_1 = RAY_AABB_io_back & RAY_AABB_io_valid_out ? RAY_AABB_io_rayid_out : 32'h0; // @[Top_1.scala 110:50 Top_1.scala 112:40 Top_1.scala 116:40]
  assign Arbitration_1_io_valid_1 = RAY_AABB_io_back & RAY_AABB_io_valid_out & RAY_AABB_io_back; // @[Top_1.scala 110:50 Top_1.scala 113:42 Top_1.scala 117:42]
  assign Arbitration_1_io_ray_id_2 = Ray_Dispatch_io_ray_out ? Ray_Dispatch_io_rayid_id : 32'h0; // @[Top_1.scala 87:43 Top_1.scala 89:56 Top_1.scala 93:56]
  assign Arbitration_1_io_valid_2 = Ray_Dispatch_io_ray_out; // @[Top_1.scala 87:33]
  assign Arbitration_1_2_clock = clock;
  assign Arbitration_1_2_reset = reset;
  assign Arbitration_1_2_io_node_id_0 = _T_111 & Stack_manage_2_io_pop_valid ? $signed(Stack_manage_2_io_node_id_out) :
    $signed(32'sh0); // @[Top_1.scala 471:85 Top_1.scala 472:49]
  assign Arbitration_1_2_io_ray_id_0 = {{32'd0}, _GEN_182}; // @[Top_1.scala 471:85 Top_1.scala 473:52]
  assign Arbitration_1_2_io_hit_0 = _T_111 & Stack_manage_2_io_pop_valid ? Stack_manage_2_io_hitT_out : 32'h0; // @[Top_1.scala 471:85 Top_1.scala 474:56]
  assign Arbitration_1_2_io_valid_0 = _T_111 & Stack_manage_2_io_pop_valid; // @[Top_1.scala 471:55]
  assign Arbitration_1_2_io_node_id_1 = RAY_AABB_2_io_back & RAY_AABB_2_io_valid_out ? $signed(RAY_AABB_2_io_nodeIdx_1)
     : $signed(32'sh0); // @[Top_1.scala 119:54 Top_1.scala 120:39 Top_1.scala 124:39]
  assign Arbitration_1_2_io_ray_id_1 = RAY_AABB_2_io_back & RAY_AABB_2_io_valid_out ? RAY_AABB_2_io_rayid_out : 32'h0; // @[Top_1.scala 119:54 Top_1.scala 121:42 Top_1.scala 125:42]
  assign Arbitration_1_2_io_valid_1 = RAY_AABB_2_io_back & RAY_AABB_2_io_valid_out & RAY_AABB_2_io_back; // @[Top_1.scala 119:54 Top_1.scala 122:44 Top_1.scala 126:44]
  assign Arbitration_1_2_io_ray_id_2 = Ray_Dispatch_io_ray_out_2 ? Ray_Dispatch_io_rayid_id_2 : 32'h0; // @[Top_1.scala 97:45 Top_1.scala 99:58 Top_1.scala 103:58]
  assign Arbitration_1_2_io_valid_2 = Ray_Dispatch_io_ray_out_2; // @[Top_1.scala 97:35]
  assign Arbitration_2_clock = clock;
  assign Arbitration_2_reset = reset;
  assign Arbitration_2_io_ray_id_2_0 = Triangle_io_break_3 & Triangle_io_RAY_AABB_1_out_IST3 ? Triangle_io_ray_id_ist3
     : 32'h0; // @[Top_1.scala 639:63 Top_1.scala 641:46 Top_1.scala 646:46]
  assign Arbitration_2_io_hit_2_0 = Triangle_io_break_3 & Triangle_io_RAY_AABB_1_out_IST3 ? Triangle_io_hiT_out_3 : 32'h0
    ; // @[Top_1.scala 639:63 Top_1.scala 642:50 Top_1.scala 647:50]
  assign Arbitration_2_io_valid_2_0 = Triangle_io_break_3 & Triangle_io_RAY_AABB_1_out_IST3; // @[Top_1.scala 639:29]
  assign Arbitration_2_io_ray_id_2_1 = Triangle_io_break_2 & Triangle_io_RAY_AABB_1_out_IST2 ? Triangle_io_ray_id_ist2
     : 32'h0; // @[Top_1.scala 615:63 Top_1.scala 617:46 Top_1.scala 622:46]
  assign Arbitration_2_io_hit_2_1 = Triangle_io_break_2 & Triangle_io_RAY_AABB_1_out_IST2 ? Triangle_io_hiT_out_2 : 32'h0
    ; // @[Top_1.scala 615:63 Top_1.scala 618:50 Top_1.scala 623:50]
  assign Arbitration_2_io_valid_2_1 = Triangle_io_break_2 & Triangle_io_RAY_AABB_1_out_IST2; // @[Top_1.scala 615:29]
  assign Arbitration_2_io_ray_id_2_2 = Triangle_io_break_1 & Triangle_io_RAY_AABB_1_out_IST1 ? Triangle_io_ray_id_ist1
     : 32'h0; // @[Top_1.scala 590:63 Top_1.scala 592:46 Top_1.scala 597:46]
  assign Arbitration_2_io_hit_2_2 = Triangle_io_break_1 & Triangle_io_RAY_AABB_1_out_IST1 ? Triangle_io_hiT_out_1 : 32'h0
    ; // @[Top_1.scala 590:63 Top_1.scala 593:50 Top_1.scala 598:50]
  assign Arbitration_2_io_valid_2_2 = Triangle_io_break_1 & Triangle_io_RAY_AABB_1_out_IST1; // @[Top_1.scala 590:29]
  assign Arbitration_2_io_ray_id_2_3 = RAY_AABB_io_pop & RAY_AABB_io_valid_out ? RAY_AABB_io_rayid_out : 32'h0; // @[Top_1.scala 251:49 Top_1.scala 253:48 Top_1.scala 258:48]
  assign Arbitration_2_io_hit_2_3 = RAY_AABB_io_pop & RAY_AABB_io_valid_out ? RAY_AABB_io_hitT_out : 32'h0; // @[Top_1.scala 251:49 Top_1.scala 254:52 Top_1.scala 259:52]
  assign Arbitration_2_io_valid_2_3 = RAY_AABB_io_pop & RAY_AABB_io_valid_out; // @[Top_1.scala 251:25]
  assign Arbitration_2_2_clock = clock;
  assign Arbitration_2_2_reset = reset;
  assign Arbitration_2_2_io_ray_id_2_0 = Triangle_io_break_3 & Triangle_io_RAY_AABB_2_out_IST3 ? Triangle_io_ray_id_ist3
     : 32'h0; // @[Top_1.scala 651:60 Top_1.scala 653:48 Top_1.scala 658:48]
  assign Arbitration_2_2_io_hit_2_0 = Triangle_io_break_3 & Triangle_io_RAY_AABB_2_out_IST3 ? Triangle_io_hiT_out_3 : 32'h0
    ; // @[Top_1.scala 651:60 Top_1.scala 654:52 Top_1.scala 659:52]
  assign Arbitration_2_2_io_valid_2_0 = Triangle_io_break_3 & Triangle_io_RAY_AABB_2_out_IST3; // @[Top_1.scala 651:26]
  assign Arbitration_2_2_io_ray_id_2_1 = Triangle_io_break_2 & Triangle_io_RAY_AABB_2_out_IST2 ? Triangle_io_ray_id_ist2
     : 32'h0; // @[Top_1.scala 626:63 Top_1.scala 628:48 Top_1.scala 633:48]
  assign Arbitration_2_2_io_hit_2_1 = Triangle_io_break_2 & Triangle_io_RAY_AABB_2_out_IST2 ? Triangle_io_hiT_out_2 : 32'h0
    ; // @[Top_1.scala 626:63 Top_1.scala 629:52 Top_1.scala 634:52]
  assign Arbitration_2_2_io_valid_2_1 = Triangle_io_break_2 & Triangle_io_RAY_AABB_2_out_IST2; // @[Top_1.scala 626:29]
  assign Arbitration_2_2_io_ray_id_2_2 = Triangle_io_break_1 & Triangle_io_RAY_AABB_2_out_IST1 ? Triangle_io_ray_id_ist1
     : 32'h0; // @[Top_1.scala 602:63 Top_1.scala 604:48 Top_1.scala 609:48]
  assign Arbitration_2_2_io_hit_2_2 = Triangle_io_break_1 & Triangle_io_RAY_AABB_2_out_IST1 ? Triangle_io_hiT_out_1 : 32'h0
    ; // @[Top_1.scala 602:63 Top_1.scala 605:52 Top_1.scala 610:52]
  assign Arbitration_2_2_io_valid_2_2 = Triangle_io_break_1 & Triangle_io_RAY_AABB_2_out_IST1; // @[Top_1.scala 602:29]
  assign Arbitration_2_2_io_ray_id_2_3 = RAY_AABB_2_io_pop & RAY_AABB_2_io_valid_out ? RAY_AABB_2_io_rayid_out : 32'h0; // @[Top_1.scala 387:53 Top_1.scala 388:50 Top_1.scala 392:50]
  assign Arbitration_2_2_io_hit_2_3 = RAY_AABB_2_io_pop & RAY_AABB_2_io_valid_out ? RAY_AABB_2_io_hitT_out : 32'h0; // @[Top_1.scala 387:53 Top_1.scala 389:54 Top_1.scala 393:54]
  assign Arbitration_2_2_io_valid_2_3 = RAY_AABB_2_io_pop & RAY_AABB_2_io_valid_out; // @[Top_1.scala 387:27]
  assign Arbitration_3_clock = clock;
  assign Arbitration_3_reset = reset;
  assign Arbitration_3_io_node_id_3_0 = Triangle_io_pop_3 & Triangle_io_RAY_AABB_1_out_IST3 ? $signed(_T_144) : $signed(32'sh0
    ); // @[Top_1.scala 565:62 Top_1.scala 566:43 Top_1.scala 571:43]
  assign Arbitration_3_io_ray_id_3_0 = Triangle_io_pop_3 & Triangle_io_RAY_AABB_1_out_IST3 ? Triangle_io_ray_id_ist3 : 32'h0
    ; // @[Top_1.scala 565:62 Top_1.scala 567:46 Top_1.scala 572:46]
  assign Arbitration_3_io_hit_3_0 = Triangle_io_pop_3 & Triangle_io_RAY_AABB_1_out_IST3 ? Triangle_io_hiT_out_3 : 32'h0; // @[Top_1.scala 565:62 Top_1.scala 568:50 Top_1.scala 573:50]
  assign Arbitration_3_io_valid_3_0 = Triangle_io_pop_3 & Triangle_io_RAY_AABB_1_out_IST3; // @[Top_1.scala 565:28]
  assign Arbitration_3_io_node_id_3_1 = Triangle_io_pop_2 & Triangle_io_RAY_AABB_1_out_IST2 ? $signed(_T_136) : $signed(32'sh0
    ); // @[Top_1.scala 541:61 Top_1.scala 542:43 Top_1.scala 547:43]
  assign Arbitration_3_io_ray_id_3_1 = Triangle_io_pop_2 & Triangle_io_RAY_AABB_1_out_IST2 ? Triangle_io_ray_id_ist2 : 32'h0
    ; // @[Top_1.scala 541:61 Top_1.scala 543:46 Top_1.scala 548:46]
  assign Arbitration_3_io_hit_3_1 = Triangle_io_pop_2 & Triangle_io_RAY_AABB_1_out_IST2 ? Triangle_io_hiT_out_2 : 32'h0; // @[Top_1.scala 541:61 Top_1.scala 544:50 Top_1.scala 549:50]
  assign Arbitration_3_io_valid_3_1 = Triangle_io_pop_2 & Triangle_io_RAY_AABB_1_out_IST2; // @[Top_1.scala 541:27]
  assign Arbitration_3_io_node_id_3_2 = Triangle_io_pop_1 & Triangle_io_RAY_AABB_1_out_IST1 ? $signed(_T_128) : $signed(32'sh0
    ); // @[Top_1.scala 516:59 Top_1.scala 517:43 Top_1.scala 522:43]
  assign Arbitration_3_io_ray_id_3_2 = Triangle_io_pop_1 & Triangle_io_RAY_AABB_1_out_IST1 ? Triangle_io_ray_id_ist1 : 32'h0
    ; // @[Top_1.scala 516:59 Top_1.scala 518:46 Top_1.scala 523:46]
  assign Arbitration_3_io_hit_3_2 = Triangle_io_pop_1 & Triangle_io_RAY_AABB_1_out_IST1 ? Triangle_io_hiT_out_1 : 32'h0; // @[Top_1.scala 516:59 Top_1.scala 519:50 Top_1.scala 524:50]
  assign Arbitration_3_io_valid_3_2 = Triangle_io_pop_1 & Triangle_io_RAY_AABB_1_out_IST1; // @[Top_1.scala 516:25]
  assign Arbitration_3_io_node_id_3_3 = ~_T_96 & Stack_manage_io_pop_valid ? $signed(_T_109) : $signed(32'sh0); // @[Top_1.scala 456:87 Top_1.scala 457:44 Top_1.scala 466:44]
  assign Arbitration_3_io_ray_id_3_3 = ~_T_96 & Stack_manage_io_pop_valid ? Stack_manage_io_ray_id_out : 32'h0; // @[Top_1.scala 456:87 Top_1.scala 458:47 Top_1.scala 467:47]
  assign Arbitration_3_io_hit_3_3 = ~_T_96 & Stack_manage_io_pop_valid ? Stack_manage_io_hitT_out : 32'h0; // @[Top_1.scala 456:87 Top_1.scala 459:52 Top_1.scala 468:52]
  assign Arbitration_3_io_valid_3_3 = ~_T_96 & Stack_manage_io_pop_valid; // @[Top_1.scala 456:59]
  assign Arbitration_3_io_node_id_3_4 = RAY_AABB_io_leaf & RAY_AABB_io_valid_out ? $signed(_T_88) : $signed(32'sh0); // @[Top_1.scala 426:50 Top_1.scala 427:45 Top_1.scala 432:45]
  assign Arbitration_3_io_ray_id_3_4 = RAY_AABB_io_leaf & RAY_AABB_io_valid_out ? RAY_AABB_io_rayid_out : 32'h0; // @[Top_1.scala 426:50 Top_1.scala 428:48 Top_1.scala 433:48]
  assign Arbitration_3_io_hit_3_4 = RAY_AABB_io_leaf & RAY_AABB_io_valid_out ? RAY_AABB_io_hitT_out : 32'h0; // @[Top_1.scala 426:50 Top_1.scala 429:52 Top_1.scala 434:52]
  assign Arbitration_3_io_valid_3_4 = RAY_AABB_io_leaf & RAY_AABB_io_valid_out; // @[Top_1.scala 426:26]
  assign Arbitration_3_2_clock = clock;
  assign Arbitration_3_2_reset = reset;
  assign Arbitration_3_2_io_node_id_3_0 = Triangle_io_pop_3 & Triangle_io_RAY_AABB_2_out_IST3 ? $signed(_T_144) :
    $signed(32'sh0); // @[Top_1.scala 576:61 Top_1.scala 577:45 Top_1.scala 582:45]
  assign Arbitration_3_2_io_ray_id_3_0 = Triangle_io_pop_3 & Triangle_io_RAY_AABB_2_out_IST3 ? Triangle_io_ray_id_ist3
     : 32'h0; // @[Top_1.scala 576:61 Top_1.scala 578:48 Top_1.scala 583:48]
  assign Arbitration_3_2_io_hit_3_0 = Triangle_io_pop_3 & Triangle_io_RAY_AABB_2_out_IST3 ? Triangle_io_hiT_out_3 : 32'h0
    ; // @[Top_1.scala 576:61 Top_1.scala 579:52 Top_1.scala 584:52]
  assign Arbitration_3_2_io_valid_3_0 = Triangle_io_pop_3 & Triangle_io_RAY_AABB_2_out_IST3; // @[Top_1.scala 576:27]
  assign Arbitration_3_2_io_node_id_3_1 = Triangle_io_pop_2 & Triangle_io_RAY_AABB_2_out_IST2 ? $signed(_T_136) :
    $signed(32'sh0); // @[Top_1.scala 552:61 Top_1.scala 553:45 Top_1.scala 558:45]
  assign Arbitration_3_2_io_ray_id_3_1 = Triangle_io_pop_2 & Triangle_io_RAY_AABB_2_out_IST2 ? Triangle_io_ray_id_ist2
     : 32'h0; // @[Top_1.scala 552:61 Top_1.scala 554:48 Top_1.scala 559:48]
  assign Arbitration_3_2_io_hit_3_1 = Triangle_io_pop_2 & Triangle_io_RAY_AABB_2_out_IST2 ? Triangle_io_hiT_out_2 : 32'h0
    ; // @[Top_1.scala 552:61 Top_1.scala 555:52 Top_1.scala 560:52]
  assign Arbitration_3_2_io_valid_3_1 = Triangle_io_pop_2 & Triangle_io_RAY_AABB_2_out_IST2; // @[Top_1.scala 552:27]
  assign Arbitration_3_2_io_node_id_3_2 = Triangle_io_pop_1 & Triangle_io_RAY_AABB_2_out_IST1 ? $signed(_T_128) :
    $signed(32'sh0); // @[Top_1.scala 528:61 Top_1.scala 529:45 Top_1.scala 534:45]
  assign Arbitration_3_2_io_ray_id_3_2 = Triangle_io_pop_1 & Triangle_io_RAY_AABB_2_out_IST1 ? Triangle_io_ray_id_ist1
     : 32'h0; // @[Top_1.scala 528:61 Top_1.scala 530:48 Top_1.scala 535:48]
  assign Arbitration_3_2_io_hit_3_2 = Triangle_io_pop_1 & Triangle_io_RAY_AABB_2_out_IST1 ? Triangle_io_hiT_out_1 : 32'h0
    ; // @[Top_1.scala 528:61 Top_1.scala 531:52 Top_1.scala 536:52]
  assign Arbitration_3_2_io_valid_3_2 = Triangle_io_pop_1 & Triangle_io_RAY_AABB_2_out_IST1; // @[Top_1.scala 528:27]
  assign Arbitration_3_2_io_node_id_3_3 = ~_T_111 & Stack_manage_2_io_pop_valid ? $signed(_T_124) : $signed(32'sh0); // @[Top_1.scala 476:91 Top_1.scala 477:46 Top_1.scala 486:46]
  assign Arbitration_3_2_io_ray_id_3_3 = ~_T_111 & Stack_manage_2_io_pop_valid ? Stack_manage_2_io_ray_id_out : 32'h0; // @[Top_1.scala 476:91 Top_1.scala 478:49 Top_1.scala 487:49]
  assign Arbitration_3_2_io_hit_3_3 = ~_T_111 & Stack_manage_2_io_pop_valid ? Stack_manage_2_io_hitT_out : 32'h0; // @[Top_1.scala 476:91 Top_1.scala 479:54 Top_1.scala 488:54]
  assign Arbitration_3_2_io_valid_3_3 = ~_T_111 & Stack_manage_2_io_pop_valid; // @[Top_1.scala 476:61]
  assign Arbitration_3_2_io_node_id_3_4 = RAY_AABB_2_io_leaf & RAY_AABB_2_io_valid_out ? $signed(_T_94) : $signed(32'sh0
    ); // @[Top_1.scala 437:54 Top_1.scala 438:47 Top_1.scala 443:47]
  assign Arbitration_3_2_io_ray_id_3_4 = RAY_AABB_2_io_leaf & RAY_AABB_2_io_valid_out ? RAY_AABB_2_io_rayid_out : 32'h0; // @[Top_1.scala 437:54 Top_1.scala 439:50 Top_1.scala 444:50]
  assign Arbitration_3_2_io_hit_3_4 = RAY_AABB_2_io_leaf & RAY_AABB_2_io_valid_out ? RAY_AABB_2_io_hitT_out : 32'h0; // @[Top_1.scala 437:54 Top_1.scala 440:54 Top_1.scala 445:54]
  assign Arbitration_3_2_io_valid_3_4 = RAY_AABB_2_io_leaf & RAY_AABB_2_io_valid_out; // @[Top_1.scala 437:28]
  assign Arbitration_4_clock = clock;
  assign Arbitration_4_reset = reset;
  assign Arbitration_4_io_node_id_4_0 = Arbitration_3_io_valid_out ? $signed(Arbitration_3_io_node_id_out) : $signed(32'sh0
    ); // @[Top_1.scala 492:37 Top_1.scala 493:43 Top_1.scala 498:43]
  assign Arbitration_4_io_ray_id_4_0 = Arbitration_3_io_valid_out ? Arbitration_3_io_ray_id_out : 32'h0; // @[Top_1.scala 492:37 Top_1.scala 494:46 Top_1.scala 499:46]
  assign Arbitration_4_io_hit_4_0 = Arbitration_3_io_valid_out ? Arbitration_3_io_hit_out : 32'h0; // @[Top_1.scala 492:37 Top_1.scala 495:50 Top_1.scala 500:50]
  assign Arbitration_4_io_valid_4_0 = Arbitration_3_io_valid_out; // @[Top_1.scala 492:37 Top_1.scala 496:47 Top_1.scala 501:48]
  assign Arbitration_4_io_node_id_4_1 = Arbitration_3_2_io_valid_out ? $signed(Arbitration_3_2_io_node_id_out) :
    $signed(32'sh0); // @[Top_1.scala 504:39 Top_1.scala 505:43 Top_1.scala 510:43]
  assign Arbitration_4_io_ray_id_4_1 = Arbitration_3_2_io_valid_out ? Arbitration_3_2_io_ray_id_out : 32'h0; // @[Top_1.scala 504:39 Top_1.scala 506:46 Top_1.scala 511:46]
  assign Arbitration_4_io_hit_4_1 = Arbitration_3_2_io_valid_out ? Arbitration_3_2_io_hit_out : 32'h0; // @[Top_1.scala 504:39 Top_1.scala 507:50 Top_1.scala 512:50]
  assign Arbitration_4_io_valid_4_1 = Arbitration_3_2_io_valid_out; // @[Top_1.scala 504:39 Top_1.scala 508:47 Top_1.scala 513:47]
  assign Stack_manage_clock = clock;
  assign Stack_manage_reset = reset;
  assign Stack_manage_io_push = RAY_AABB_io_push & RAY_AABB_io_valid_out; // @[Top_1.scala 401:26]
  assign Stack_manage_io_push_en = RAY_AABB_io_push & RAY_AABB_io_valid_out; // @[Top_1.scala 401:26]
  assign Stack_manage_io_pop = Arbitration_2_io_valid_out; // @[Top_1.scala 755:46]
  assign Stack_manage_io_pop_en = Arbitration_2_io_valid_out; // @[Top_1.scala 756:42]
  assign Stack_manage_io_ray_id_push = RAY_AABB_io_push & RAY_AABB_io_valid_out ? RAY_AABB_io_rayid_out : 32'h0; // @[Top_1.scala 401:50 Top_1.scala 405:52 Top_1.scala 410:53]
  assign Stack_manage_io_ray_id_pop = Arbitration_2_io_ray_id_out; // @[Top_1.scala 757:38]
  assign Stack_manage_io_node_id_push_in = RAY_AABB_io_push & RAY_AABB_io_valid_out ? $signed(RAY_AABB_io_nodeIdx_0) :
    $signed(32'sh0); // @[Top_1.scala 401:50 Top_1.scala 404:45 Top_1.scala 409:47]
  assign Stack_manage_io_hitT_in = Arbitration_2_io_hit_out; // @[Top_1.scala 758:44]
  assign Stack_manage_2_clock = clock;
  assign Stack_manage_2_reset = reset;
  assign Stack_manage_2_io_push = RAY_AABB_2_io_push & RAY_AABB_2_io_valid_out; // @[Top_1.scala 413:28]
  assign Stack_manage_2_io_push_en = RAY_AABB_2_io_push & RAY_AABB_2_io_valid_out; // @[Top_1.scala 413:28]
  assign Stack_manage_2_io_pop = Arbitration_2_2_io_valid_out; // @[Top_1.scala 760:48]
  assign Stack_manage_2_io_pop_en = Arbitration_2_2_io_valid_out; // @[Top_1.scala 761:44]
  assign Stack_manage_2_io_ray_id_push = RAY_AABB_2_io_push & RAY_AABB_2_io_valid_out ? RAY_AABB_2_io_rayid_out : 32'h0; // @[Top_1.scala 413:54 Top_1.scala 417:54 Top_1.scala 422:55]
  assign Stack_manage_2_io_ray_id_pop = Arbitration_2_2_io_ray_id_out; // @[Top_1.scala 762:40]
  assign Stack_manage_2_io_node_id_push_in = RAY_AABB_2_io_push & RAY_AABB_2_io_valid_out ? $signed(
    RAY_AABB_2_io_nodeIdx_0) : $signed(32'sh0); // @[Top_1.scala 413:54 Top_1.scala 416:47 Top_1.scala 421:49]
  assign Stack_manage_2_io_hitT_in = Arbitration_2_2_io_hit_out; // @[Top_1.scala 763:46]
  assign Triangle_clock = clock;
  assign Triangle_reset = reset;
  assign Triangle_io_To_IST0_enable = leaf_memory_valid; // @[Top_1.scala 698:34 Top_1.scala 699:42 Top_1.scala 726:42]
  assign Triangle_io_nodeid_leaf = leaf_memory_valid ? $signed(leaf_node_id_temp) : $signed(32'sh0); // @[Top_1.scala 698:34 Top_1.scala 700:47 Top_1.scala 727:47]
  assign Triangle_io_rayid_leaf = leaf_memory_valid ? ray_leaf_temp : 32'h0; // @[Top_1.scala 698:34 Top_1.scala 701:50 Top_1.scala 728:50]
  assign Triangle_io_hiT_in = leaf_memory_valid ? hitT_temp : 32'h0; // @[Top_1.scala 698:34 Top_1.scala 702:54 Top_1.scala 729:54]
  assign Triangle_io_v00_in_x = leaf_memory_valid ? TRI_RAM_x_io_v00_out : 32'h0; // @[Top_1.scala 698:34 Top_1.scala 703:52 Top_1.scala 730:52]
  assign Triangle_io_v00_in_y = leaf_memory_valid ? TRI_RAM_y_io_v00_out : 32'h0; // @[Top_1.scala 698:34 Top_1.scala 705:52 Top_1.scala 732:52]
  assign Triangle_io_v00_in_z = leaf_memory_valid ? TRI_RAM_z_io_v00_out : 32'h0; // @[Top_1.scala 698:34 Top_1.scala 706:52 Top_1.scala 733:52]
  assign Triangle_io_v00_in_w = leaf_memory_valid ? TRI_RAM_w_io_v00_out : 32'h0; // @[Top_1.scala 698:34 Top_1.scala 707:51 Top_1.scala 734:51]
  assign Triangle_io_v11_in_x = leaf_memory_valid ? TRI_RAM_x_io_v11_out : 32'h0; // @[Top_1.scala 698:34 Top_1.scala 708:52 Top_1.scala 735:52]
  assign Triangle_io_v11_in_y = leaf_memory_valid ? TRI_RAM_y_io_v11_out : 32'h0; // @[Top_1.scala 698:34 Top_1.scala 709:52 Top_1.scala 736:52]
  assign Triangle_io_v11_in_z = leaf_memory_valid ? TRI_RAM_z_io_v11_out : 32'h0; // @[Top_1.scala 698:34 Top_1.scala 710:52 Top_1.scala 737:52]
  assign Triangle_io_v11_in_w = leaf_memory_valid ? TRI_RAM_w_io_v11_out : 32'h0; // @[Top_1.scala 698:34 Top_1.scala 711:51 Top_1.scala 738:51]
  assign Triangle_io_v22_in_x = leaf_memory_valid ? TRI_RAM_x_io_v22_out : 32'h0; // @[Top_1.scala 698:34 Top_1.scala 712:52 Top_1.scala 739:52]
  assign Triangle_io_v22_in_y = leaf_memory_valid ? TRI_RAM_y_io_v22_out : 32'h0; // @[Top_1.scala 698:34 Top_1.scala 713:52 Top_1.scala 740:52]
  assign Triangle_io_v22_in_z = leaf_memory_valid ? TRI_RAM_z_io_v22_out : 32'h0; // @[Top_1.scala 698:34 Top_1.scala 714:52 Top_1.scala 741:52]
  assign Triangle_io_v22_in_w = leaf_memory_valid ? TRI_RAM_w_io_v22_out : 32'h0; // @[Top_1.scala 698:34 Top_1.scala 715:51 Top_1.scala 742:51]
  assign Triangle_io_ray_o_in_x = leaf_memory_valid ? Ray_origx_io_Ray_out : 32'h0; // @[Top_1.scala 698:34 Top_1.scala 716:50 Top_1.scala 743:50]
  assign Triangle_io_ray_o_in_y = leaf_memory_valid ? Ray_origy_io_Ray_out : 32'h0; // @[Top_1.scala 698:34 Top_1.scala 717:50 Top_1.scala 744:50]
  assign Triangle_io_ray_o_in_z = leaf_memory_valid ? Ray_origz_io_Ray_out : 32'h0; // @[Top_1.scala 698:34 Top_1.scala 718:50 Top_1.scala 745:50]
  assign Triangle_io_ray_d_in_x = leaf_memory_valid ? Ray_dirx_io_Ray_out : 32'h0; // @[Top_1.scala 698:34 Top_1.scala 719:50 Top_1.scala 746:50]
  assign Triangle_io_ray_d_in_y = leaf_memory_valid ? Ray_diry_io_Ray_out : 32'h0; // @[Top_1.scala 698:34 Top_1.scala 720:50 Top_1.scala 747:50]
  assign Triangle_io_ray_d_in_z = leaf_memory_valid ? Ray_dirz_io_Ray_out : 32'h0; // @[Top_1.scala 698:34 Top_1.scala 721:50 Top_1.scala 748:50]
  assign Triangle_io_break_in = leaf_memory_valid & TRI_RAM_x_io_valid == 32'h80000000; // @[Top_1.scala 698:34 Top_1.scala 704:51 Top_1.scala 731:51]
  assign Triangle_io_RAY_AABB_1 = leaf_memory_valid & ray_aabb; // @[Top_1.scala 698:34 Top_1.scala 722:45 Top_1.scala 749:45]
  assign Triangle_io_RAY_AABB_2 = leaf_memory_valid & ray_aabb_2; // @[Top_1.scala 698:34 Top_1.scala 723:45 Top_1.scala 750:45]
  always @(posedge clock) begin
    if (reset) begin // @[Top_1.scala 79:42]
      clock_counter <= 64'h0; // @[Top_1.scala 79:42]
    end else begin
      clock_counter <= _T_1; // @[Top_1.scala 80:36]
    end
    if (reset) begin // @[Top_1.scala 129:54]
      memory_valid <= 1'h0; // @[Top_1.scala 129:54]
    end else begin
      memory_valid <= _GEN_31;
    end
    if (reset) begin // @[Top_1.scala 130:61]
      hit_temp <= 32'h0; // @[Top_1.scala 130:61]
    end else if (Arbitration_1_io_valid_out & Arbitration_1_io_hit_out != 32'h0) begin // @[Top_1.scala 134:70]
      hit_temp <= Arbitration_1_io_hit_out; // @[Top_1.scala 142:51]
    end else begin
      hit_temp <= 32'h0;
    end
    if (reset) begin // @[Top_1.scala 131:57]
      ray_id_temp <= 32'h0; // @[Top_1.scala 131:57]
    end else if (Arbitration_1_io_valid_out & Arbitration_1_io_hit_out != 32'h0) begin // @[Top_1.scala 134:70]
      ray_id_temp <= Arbitration_1_io_ray_id_out; // @[Top_1.scala 157:59]
    end else if (Arbitration_1_io_valid_out & Arbitration_1_io_hit_out == 32'h0) begin // @[Top_1.scala 159:76]
      ray_id_temp <= Arbitration_1_io_ray_id_out; // @[Top_1.scala 183:59]
    end
    if (reset) begin // @[Top_1.scala 132:57]
      hit_from_arb <= 1'h0; // @[Top_1.scala 132:57]
    end else begin
      hit_from_arb <= _T_8;
    end
    if (reset) begin // @[Top_1.scala 133:64]
      TRV_1 <= 64'h0; // @[Top_1.scala 133:64]
    end else if (memory_valid) begin // @[Top_1.scala 190:29]
      TRV_1 <= _T_42; // @[Top_1.scala 222:70]
    end
    if (reset) begin // @[Top_1.scala 264:56]
      memory_valid_2 <= 1'h0; // @[Top_1.scala 264:56]
    end else begin
      memory_valid_2 <= _GEN_98;
    end
    if (reset) begin // @[Top_1.scala 265:63]
      hit_temp_2 <= 32'h0; // @[Top_1.scala 265:63]
    end else if (Arbitration_1_2_io_valid_out & Arbitration_1_2_io_hit_out != 32'h0) begin // @[Top_1.scala 269:74]
      hit_temp_2 <= Arbitration_1_2_io_hit_out; // @[Top_1.scala 279:65]
    end else begin
      hit_temp_2 <= 32'h0;
    end
    if (reset) begin // @[Top_1.scala 266:59]
      ray_id_temp_2 <= 32'h0; // @[Top_1.scala 266:59]
    end else if (Arbitration_1_2_io_valid_out & Arbitration_1_2_io_hit_out != 32'h0) begin // @[Top_1.scala 269:74]
      ray_id_temp_2 <= Arbitration_1_2_io_ray_id_out; // @[Top_1.scala 294:61]
    end else if (Arbitration_1_2_io_valid_out & Arbitration_1_2_io_hit_out == 32'h0) begin // @[Top_1.scala 296:80]
      ray_id_temp_2 <= Arbitration_1_2_io_ray_id_out; // @[Top_1.scala 322:61]
    end
    if (reset) begin // @[Top_1.scala 267:59]
      hit_from_arb_2 <= 1'h0; // @[Top_1.scala 267:59]
    end else begin
      hit_from_arb_2 <= _T_45;
    end
    if (reset) begin // @[Top_1.scala 268:70]
      TRV_2 <= 64'h0; // @[Top_1.scala 268:70]
    end else if (memory_valid_2) begin // @[Top_1.scala 329:31]
      TRV_2 <= _T_79; // @[Top_1.scala 358:76]
    end
    if (reset) begin // @[Top_1.scala 666:58]
      leaf_memory_valid <= 1'h0; // @[Top_1.scala 666:58]
    end else begin
      leaf_memory_valid <= _GEN_239;
    end
    if (reset) begin // @[Top_1.scala 667:68]
      hitT_temp <= 32'h0; // @[Top_1.scala 667:68]
    end else if (Arbitration_4_io_valid_out) begin // @[Top_1.scala 673:37]
      hitT_temp <= Arbitration_4_io_hit_out; // @[Top_1.scala 685:55]
    end else begin
      hitT_temp <= 32'h0; // @[Top_1.scala 692:61]
    end
    if (reset) begin // @[Top_1.scala 668:64]
      ray_leaf_temp <= 32'h0; // @[Top_1.scala 668:64]
    end else if (Arbitration_4_io_valid_out) begin // @[Top_1.scala 673:37]
      ray_leaf_temp <= Arbitration_4_io_ray_id_out; // @[Top_1.scala 686:55]
    end else begin
      ray_leaf_temp <= 32'h0; // @[Top_1.scala 693:57]
    end
    if (reset) begin // @[Top_1.scala 669:57]
      leaf_node_id_temp <= 32'sh0; // @[Top_1.scala 669:57]
    end else if (Arbitration_4_io_valid_out) begin // @[Top_1.scala 673:37]
      leaf_node_id_temp <= Arbitration_4_io_node_id_out; // @[Top_1.scala 687:55]
    end else begin
      leaf_node_id_temp <= 32'sh0; // @[Top_1.scala 694:50]
    end
    if (reset) begin // @[Top_1.scala 670:69]
      ray_aabb <= 1'h0; // @[Top_1.scala 670:69]
    end else begin
      ray_aabb <= _GEN_245;
    end
    if (reset) begin // @[Top_1.scala 671:71]
      ray_aabb_2 <= 1'h0; // @[Top_1.scala 671:71]
    end else begin
      ray_aabb_2 <= _GEN_246;
    end
    if (reset) begin // @[Top_1.scala 672:75]
      IST_1 <= 64'h0; // @[Top_1.scala 672:75]
    end else if (leaf_memory_valid) begin // @[Top_1.scala 698:34]
      IST_1 <= _T_159; // @[Top_1.scala 724:67]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  clock_counter = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  memory_valid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  hit_temp = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  ray_id_temp = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  hit_from_arb = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  TRV_1 = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  memory_valid_2 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  hit_temp_2 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  ray_id_temp_2 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  hit_from_arb_2 = _RAND_9[0:0];
  _RAND_10 = {2{`RANDOM}};
  TRV_2 = _RAND_10[63:0];
  _RAND_11 = {1{`RANDOM}};
  leaf_memory_valid = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  hitT_temp = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  ray_leaf_temp = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  leaf_node_id_temp = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  ray_aabb = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  ray_aabb_2 = _RAND_16[0:0];
  _RAND_17 = {2{`RANDOM}};
  IST_1 = _RAND_17[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
